magic
tech sky130A
magscale 1 2
timestamp 1682557845
<< viali >>
rect 1593 24361 1627 24395
rect 6561 24361 6595 24395
rect 18153 24361 18187 24395
rect 19625 24361 19659 24395
rect 19993 24361 20027 24395
rect 22017 24361 22051 24395
rect 22458 24361 22492 24395
rect 23949 24361 23983 24395
rect 3985 24293 4019 24327
rect 17969 24293 18003 24327
rect 20177 24293 20211 24327
rect 21189 24293 21223 24327
rect 24593 24293 24627 24327
rect 3249 24225 3283 24259
rect 8401 24225 8435 24259
rect 10977 24225 11011 24259
rect 12817 24225 12851 24259
rect 14749 24225 14783 24259
rect 17417 24225 17451 24259
rect 17601 24225 17635 24259
rect 18705 24225 18739 24259
rect 20729 24225 20763 24259
rect 21833 24225 21867 24259
rect 22201 24225 22235 24259
rect 25237 24225 25271 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6745 24157 6779 24191
rect 7205 24157 7239 24191
rect 9781 24157 9815 24191
rect 11897 24157 11931 24191
rect 12357 24157 12391 24191
rect 14289 24157 14323 24191
rect 16313 24157 16347 24191
rect 18521 24157 18555 24191
rect 21373 24157 21407 24191
rect 24961 24157 24995 24191
rect 5825 24089 5859 24123
rect 17325 24089 17359 24123
rect 19533 24089 19567 24123
rect 20637 24089 20671 24123
rect 21557 24089 21591 24123
rect 1777 24021 1811 24055
rect 9137 24021 9171 24055
rect 11713 24021 11747 24055
rect 16129 24021 16163 24055
rect 16957 24021 16991 24055
rect 18613 24021 18647 24055
rect 19349 24021 19383 24055
rect 20545 24021 20579 24055
rect 25053 24021 25087 24055
rect 2329 23817 2363 23851
rect 13829 23817 13863 23851
rect 14473 23817 14507 23851
rect 16865 23817 16899 23851
rect 20361 23817 20395 23851
rect 15945 23749 15979 23783
rect 17233 23749 17267 23783
rect 20729 23749 20763 23783
rect 22937 23749 22971 23783
rect 1685 23681 1719 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 6561 23681 6595 23715
rect 6837 23681 6871 23715
rect 7941 23681 7975 23715
rect 9137 23681 9171 23715
rect 9965 23681 9999 23715
rect 10885 23681 10919 23715
rect 12081 23681 12115 23715
rect 15301 23681 15335 23715
rect 17325 23681 17359 23715
rect 20821 23681 20855 23715
rect 22201 23681 22235 23715
rect 25053 23681 25087 23715
rect 3985 23613 4019 23647
rect 5825 23613 5859 23647
rect 12541 23613 12575 23647
rect 14565 23613 14599 23647
rect 14657 23613 14691 23647
rect 16313 23613 16347 23647
rect 17509 23613 17543 23647
rect 18061 23613 18095 23647
rect 18337 23613 18371 23647
rect 20913 23613 20947 23647
rect 22661 23613 22695 23647
rect 14105 23545 14139 23579
rect 22017 23545 22051 23579
rect 25237 23545 25271 23579
rect 7481 23477 7515 23511
rect 11621 23477 11655 23511
rect 11713 23477 11747 23511
rect 16497 23477 16531 23511
rect 19809 23477 19843 23511
rect 21373 23477 21407 23511
rect 21557 23477 21591 23511
rect 24409 23477 24443 23511
rect 1593 23273 1627 23307
rect 4905 23273 4939 23307
rect 18981 23273 19015 23307
rect 21189 23273 21223 23307
rect 24409 23273 24443 23307
rect 18705 23205 18739 23239
rect 3249 23137 3283 23171
rect 6469 23137 6503 23171
rect 8217 23137 8251 23171
rect 10609 23137 10643 23171
rect 17785 23137 17819 23171
rect 19441 23137 19475 23171
rect 21649 23137 21683 23171
rect 25053 23137 25087 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 4261 23069 4295 23103
rect 5457 23069 5491 23103
rect 7205 23069 7239 23103
rect 9229 23069 9263 23103
rect 9505 23069 9539 23103
rect 13093 23069 13127 23103
rect 15025 23069 15059 23103
rect 17601 23069 17635 23103
rect 24961 23069 24995 23103
rect 9045 23001 9079 23035
rect 10885 23001 10919 23035
rect 14381 23001 14415 23035
rect 14565 23001 14599 23035
rect 15301 23001 15335 23035
rect 18521 23001 18555 23035
rect 19717 23001 19751 23035
rect 21925 23001 21959 23035
rect 1777 22933 1811 22967
rect 3985 22933 4019 22967
rect 10149 22933 10183 22967
rect 12357 22933 12391 22967
rect 12725 22933 12759 22967
rect 13737 22933 13771 22967
rect 16773 22933 16807 22967
rect 17233 22933 17267 22967
rect 17693 22933 17727 22967
rect 23397 22933 23431 22967
rect 23857 22933 23891 22967
rect 24593 22933 24627 22967
rect 6561 22729 6595 22763
rect 7021 22729 7055 22763
rect 18061 22729 18095 22763
rect 18521 22729 18555 22763
rect 20453 22729 20487 22763
rect 24869 22729 24903 22763
rect 3985 22661 4019 22695
rect 5733 22661 5767 22695
rect 8769 22661 8803 22695
rect 17233 22661 17267 22695
rect 1685 22593 1719 22627
rect 2973 22593 3007 22627
rect 4813 22593 4847 22627
rect 6929 22593 6963 22627
rect 7573 22593 7607 22627
rect 9413 22593 9447 22627
rect 11989 22593 12023 22627
rect 13185 22593 13219 22627
rect 13645 22593 13679 22627
rect 15945 22593 15979 22627
rect 16129 22593 16163 22627
rect 17325 22593 17359 22627
rect 18429 22593 18463 22627
rect 19625 22593 19659 22627
rect 20821 22593 20855 22627
rect 21465 22593 21499 22627
rect 22017 22593 22051 22627
rect 22937 22593 22971 22627
rect 23121 22593 23155 22627
rect 9689 22525 9723 22559
rect 11713 22525 11747 22559
rect 13921 22525 13955 22559
rect 17417 22525 17451 22559
rect 18705 22525 18739 22559
rect 19717 22525 19751 22559
rect 19809 22525 19843 22559
rect 20913 22525 20947 22559
rect 21005 22525 21039 22559
rect 22661 22525 22695 22559
rect 23397 22525 23431 22559
rect 25145 22525 25179 22559
rect 16405 22457 16439 22491
rect 16865 22457 16899 22491
rect 25329 22457 25363 22491
rect 2329 22389 2363 22423
rect 11161 22389 11195 22423
rect 13001 22389 13035 22423
rect 15393 22389 15427 22423
rect 19257 22389 19291 22423
rect 1593 22185 1627 22219
rect 13461 22185 13495 22219
rect 16018 22185 16052 22219
rect 20618 22185 20652 22219
rect 1777 22049 1811 22083
rect 3249 22049 3283 22083
rect 8125 22049 8159 22083
rect 9137 22049 9171 22083
rect 13001 22049 13035 22083
rect 14841 22049 14875 22083
rect 15761 22049 15795 22083
rect 18521 22049 18555 22083
rect 19717 22049 19751 22083
rect 22109 22049 22143 22083
rect 23857 22049 23891 22083
rect 25145 22049 25179 22083
rect 2053 21981 2087 22015
rect 4261 21981 4295 22015
rect 5457 21981 5491 22015
rect 7389 21981 7423 22015
rect 9505 21981 9539 22015
rect 10609 21981 10643 22015
rect 12817 21981 12851 22015
rect 13645 21981 13679 22015
rect 14657 21981 14691 22015
rect 18337 21981 18371 22015
rect 20361 21981 20395 22015
rect 22385 21981 22419 22015
rect 25053 21981 25087 22015
rect 6285 21913 6319 21947
rect 10149 21913 10183 21947
rect 11529 21913 11563 21947
rect 13921 21913 13955 21947
rect 14749 21913 14783 21947
rect 19533 21913 19567 21947
rect 22753 21913 22787 21947
rect 23121 21913 23155 21947
rect 3893 21845 3927 21879
rect 4905 21845 4939 21879
rect 9045 21845 9079 21879
rect 12449 21845 12483 21879
rect 12909 21845 12943 21879
rect 14289 21845 14323 21879
rect 15301 21845 15335 21879
rect 17509 21845 17543 21879
rect 17969 21845 18003 21879
rect 18429 21845 18463 21879
rect 18981 21845 19015 21879
rect 19993 21845 20027 21879
rect 22569 21845 22603 21879
rect 24593 21845 24627 21879
rect 24961 21845 24995 21879
rect 2329 21641 2363 21675
rect 11897 21641 11931 21675
rect 12633 21641 12667 21675
rect 16865 21641 16899 21675
rect 22477 21641 22511 21675
rect 25421 21641 25455 21675
rect 13737 21573 13771 21607
rect 18613 21573 18647 21607
rect 23581 21573 23615 21607
rect 1685 21505 1719 21539
rect 2789 21505 2823 21539
rect 4813 21505 4847 21539
rect 7113 21505 7147 21539
rect 8953 21505 8987 21539
rect 11069 21505 11103 21539
rect 11253 21505 11287 21539
rect 13461 21505 13495 21539
rect 15669 21505 15703 21539
rect 17233 21505 17267 21539
rect 18337 21505 18371 21539
rect 21097 21505 21131 21539
rect 23305 21505 23339 21539
rect 3525 21437 3559 21471
rect 5089 21437 5123 21471
rect 6745 21437 6779 21471
rect 7573 21437 7607 21471
rect 12725 21437 12759 21471
rect 12909 21437 12943 21471
rect 17325 21437 17359 21471
rect 17417 21437 17451 21471
rect 17877 21437 17911 21471
rect 20085 21437 20119 21471
rect 21189 21437 21223 21471
rect 21281 21437 21315 21471
rect 22569 21437 22603 21471
rect 22661 21437 22695 21471
rect 6469 21301 6503 21335
rect 6653 21301 6687 21335
rect 9210 21301 9244 21335
rect 10701 21301 10735 21335
rect 11621 21301 11655 21335
rect 11713 21301 11747 21335
rect 12265 21301 12299 21335
rect 15209 21301 15243 21335
rect 16313 21301 16347 21335
rect 20361 21301 20395 21335
rect 20729 21301 20763 21335
rect 22109 21301 22143 21335
rect 25053 21301 25087 21335
rect 1777 21097 1811 21131
rect 6469 21097 6503 21131
rect 9413 21097 9447 21131
rect 15301 21097 15335 21131
rect 1593 21029 1627 21063
rect 16497 21029 16531 21063
rect 21189 21029 21223 21063
rect 21557 21029 21591 21063
rect 24593 21029 24627 21063
rect 2789 20961 2823 20995
rect 4445 20961 4479 20995
rect 7389 20961 7423 20995
rect 9781 20961 9815 20995
rect 10425 20961 10459 20995
rect 10609 20961 10643 20995
rect 11161 20961 11195 20995
rect 15853 20961 15887 20995
rect 17049 20961 17083 20995
rect 18153 20961 18187 20995
rect 18245 20961 18279 20995
rect 19441 20961 19475 20995
rect 22753 20961 22787 20995
rect 23857 20961 23891 20995
rect 25145 20961 25179 20995
rect 2237 20893 2271 20927
rect 4077 20893 4111 20927
rect 5825 20893 5859 20927
rect 7113 20893 7147 20927
rect 8769 20893 8803 20927
rect 9321 20893 9355 20927
rect 10333 20893 10367 20927
rect 13553 20893 13587 20927
rect 13737 20893 13771 20927
rect 14289 20893 14323 20927
rect 15669 20893 15703 20927
rect 15761 20893 15795 20927
rect 16957 20893 16991 20927
rect 23765 20893 23799 20927
rect 24961 20893 24995 20927
rect 11437 20825 11471 20859
rect 14565 20825 14599 20859
rect 18705 20825 18739 20859
rect 19717 20825 19751 20859
rect 25053 20825 25087 20859
rect 9965 20757 9999 20791
rect 12909 20757 12943 20791
rect 16865 20757 16899 20791
rect 17693 20757 17727 20791
rect 18061 20757 18095 20791
rect 19073 20757 19107 20791
rect 21741 20757 21775 20791
rect 22109 20757 22143 20791
rect 22477 20757 22511 20791
rect 22569 20757 22603 20791
rect 23305 20757 23339 20791
rect 23673 20757 23707 20791
rect 1501 20553 1535 20587
rect 4721 20553 4755 20587
rect 6009 20553 6043 20587
rect 8493 20553 8527 20587
rect 15393 20553 15427 20587
rect 21097 20553 21131 20587
rect 22385 20553 22419 20587
rect 23121 20553 23155 20587
rect 7389 20485 7423 20519
rect 11069 20485 11103 20519
rect 12449 20485 12483 20519
rect 13277 20485 13311 20519
rect 13921 20485 13955 20519
rect 15945 20485 15979 20519
rect 16497 20485 16531 20519
rect 16773 20485 16807 20519
rect 1777 20417 1811 20451
rect 3065 20417 3099 20451
rect 4905 20417 4939 20451
rect 5365 20417 5399 20451
rect 6745 20417 6779 20451
rect 7849 20417 7883 20451
rect 8953 20417 8987 20451
rect 13185 20417 13219 20451
rect 13652 20417 13686 20451
rect 17141 20417 17175 20451
rect 19809 20417 19843 20451
rect 19901 20417 19935 20451
rect 21005 20417 21039 20451
rect 23489 20417 23523 20451
rect 3341 20349 3375 20383
rect 9229 20349 9263 20383
rect 11253 20349 11287 20383
rect 12541 20349 12575 20383
rect 12633 20349 12667 20383
rect 16129 20349 16163 20383
rect 17417 20349 17451 20383
rect 19993 20349 20027 20383
rect 21281 20349 21315 20383
rect 22477 20349 22511 20383
rect 22661 20349 22695 20383
rect 23765 20349 23799 20383
rect 11621 20281 11655 20315
rect 2421 20213 2455 20247
rect 6469 20213 6503 20247
rect 10701 20213 10735 20247
rect 11713 20213 11747 20247
rect 12081 20213 12115 20247
rect 18889 20213 18923 20247
rect 19349 20213 19383 20247
rect 19441 20213 19475 20247
rect 20637 20213 20671 20247
rect 22017 20213 22051 20247
rect 25237 20213 25271 20247
rect 3985 20009 4019 20043
rect 16129 20009 16163 20043
rect 17785 20009 17819 20043
rect 13277 19941 13311 19975
rect 13737 19941 13771 19975
rect 13921 19941 13955 19975
rect 19441 19941 19475 19975
rect 2789 19873 2823 19907
rect 9689 19873 9723 19907
rect 10885 19873 10919 19907
rect 15485 19873 15519 19907
rect 16681 19873 16715 19907
rect 17417 19873 17451 19907
rect 18337 19873 18371 19907
rect 19993 19873 20027 19907
rect 20913 19873 20947 19907
rect 23673 19873 23707 19907
rect 25145 19873 25179 19907
rect 2237 19805 2271 19839
rect 4169 19805 4203 19839
rect 4629 19805 4663 19839
rect 5733 19805 5767 19839
rect 6837 19805 6871 19839
rect 7481 19805 7515 19839
rect 7941 19805 7975 19839
rect 11529 19805 11563 19839
rect 15301 19805 15335 19839
rect 16589 19805 16623 19839
rect 17325 19805 17359 19839
rect 18245 19805 18279 19839
rect 24133 19805 24167 19839
rect 1777 19737 1811 19771
rect 8585 19737 8619 19771
rect 11805 19737 11839 19771
rect 15393 19737 15427 19771
rect 19901 19737 19935 19771
rect 20821 19737 20855 19771
rect 21189 19737 21223 19771
rect 25053 19737 25087 19771
rect 5273 19669 5307 19703
rect 6377 19669 6411 19703
rect 9137 19669 9171 19703
rect 9505 19669 9539 19703
rect 9597 19669 9631 19703
rect 10333 19669 10367 19703
rect 10701 19669 10735 19703
rect 10793 19669 10827 19703
rect 14289 19669 14323 19703
rect 14933 19669 14967 19703
rect 16497 19669 16531 19703
rect 17601 19669 17635 19703
rect 18153 19669 18187 19703
rect 18797 19669 18831 19703
rect 18981 19669 19015 19703
rect 19349 19669 19383 19703
rect 19809 19669 19843 19703
rect 20269 19669 20303 19703
rect 20453 19669 20487 19703
rect 22661 19669 22695 19703
rect 23121 19669 23155 19703
rect 23489 19669 23523 19703
rect 23581 19669 23615 19703
rect 24593 19669 24627 19703
rect 24961 19669 24995 19703
rect 3617 19465 3651 19499
rect 6009 19465 6043 19499
rect 7389 19465 7423 19499
rect 10701 19465 10735 19499
rect 14749 19465 14783 19499
rect 15209 19465 15243 19499
rect 19625 19465 19659 19499
rect 20913 19465 20947 19499
rect 22017 19465 22051 19499
rect 22385 19465 22419 19499
rect 25053 19465 25087 19499
rect 8493 19397 8527 19431
rect 12081 19397 12115 19431
rect 12817 19397 12851 19431
rect 19717 19397 19751 19431
rect 1961 19329 1995 19363
rect 3801 19329 3835 19363
rect 4261 19329 4295 19363
rect 5365 19329 5399 19363
rect 6745 19329 6779 19363
rect 7849 19329 7883 19363
rect 8953 19329 8987 19363
rect 11345 19329 11379 19363
rect 11897 19329 11931 19363
rect 12541 19329 12575 19363
rect 15117 19329 15151 19363
rect 16129 19329 16163 19363
rect 17049 19329 17083 19363
rect 20821 19329 20855 19363
rect 22477 19329 22511 19363
rect 23305 19329 23339 19363
rect 2237 19261 2271 19295
rect 4905 19261 4939 19295
rect 9229 19261 9263 19295
rect 11161 19261 11195 19295
rect 15301 19261 15335 19295
rect 17325 19261 17359 19295
rect 19809 19261 19843 19295
rect 21005 19261 21039 19295
rect 22661 19261 22695 19295
rect 23581 19261 23615 19295
rect 6377 19193 6411 19227
rect 25421 19193 25455 19227
rect 14289 19125 14323 19159
rect 16221 19125 16255 19159
rect 16773 19125 16807 19159
rect 18797 19125 18831 19159
rect 19257 19125 19291 19159
rect 20453 19125 20487 19159
rect 21465 19125 21499 19159
rect 9229 18921 9263 18955
rect 12449 18921 12483 18955
rect 14289 18921 14323 18955
rect 13001 18853 13035 18887
rect 17325 18853 17359 18887
rect 18061 18853 18095 18887
rect 23949 18853 23983 18887
rect 9781 18785 9815 18819
rect 13461 18785 13495 18819
rect 13645 18785 13679 18819
rect 14933 18785 14967 18819
rect 15853 18785 15887 18819
rect 18613 18785 18647 18819
rect 20269 18785 20303 18819
rect 20545 18785 20579 18819
rect 23121 18785 23155 18819
rect 25053 18785 25087 18819
rect 25145 18785 25179 18819
rect 1685 18717 1719 18751
rect 2789 18717 2823 18751
rect 4629 18717 4663 18751
rect 5733 18717 5767 18751
rect 6837 18717 6871 18751
rect 7941 18717 7975 18751
rect 10425 18717 10459 18751
rect 12725 18717 12759 18751
rect 15577 18717 15611 18751
rect 19625 18717 19659 18751
rect 22937 18717 22971 18751
rect 9597 18649 9631 18683
rect 13369 18649 13403 18683
rect 14749 18649 14783 18683
rect 23765 18649 23799 18683
rect 2329 18581 2363 18615
rect 3433 18581 3467 18615
rect 3985 18581 4019 18615
rect 5273 18581 5307 18615
rect 6377 18581 6411 18615
rect 7481 18581 7515 18615
rect 8585 18581 8619 18615
rect 9689 18581 9723 18615
rect 11713 18581 11747 18615
rect 14657 18581 14691 18615
rect 17601 18581 17635 18615
rect 18429 18581 18463 18615
rect 18521 18581 18555 18615
rect 19717 18581 19751 18615
rect 22017 18581 22051 18615
rect 22477 18581 22511 18615
rect 22845 18581 22879 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 3801 18377 3835 18411
rect 6009 18377 6043 18411
rect 6377 18377 6411 18411
rect 10701 18377 10735 18411
rect 14289 18377 14323 18411
rect 15025 18377 15059 18411
rect 15301 18377 15335 18411
rect 16037 18377 16071 18411
rect 16681 18377 16715 18411
rect 23305 18377 23339 18411
rect 24869 18377 24903 18411
rect 4905 18309 4939 18343
rect 9229 18309 9263 18343
rect 13001 18309 13035 18343
rect 18245 18309 18279 18343
rect 19993 18309 20027 18343
rect 22017 18309 22051 18343
rect 25329 18309 25363 18343
rect 2053 18241 2087 18275
rect 3157 18241 3191 18275
rect 4261 18241 4295 18275
rect 5365 18241 5399 18275
rect 6745 18241 6779 18275
rect 7849 18241 7883 18275
rect 8953 18241 8987 18275
rect 12173 18241 12207 18275
rect 15945 18241 15979 18275
rect 17417 18241 17451 18275
rect 20821 18241 20855 18275
rect 20913 18241 20947 18275
rect 21465 18241 21499 18275
rect 24225 18241 24259 18275
rect 2697 18173 2731 18207
rect 11253 18173 11287 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 16129 18173 16163 18207
rect 17509 18173 17543 18207
rect 17693 18173 17727 18207
rect 21005 18173 21039 18207
rect 15577 18105 15611 18139
rect 25145 18105 25179 18139
rect 1685 18037 1719 18071
rect 7389 18037 7423 18071
rect 8493 18037 8527 18071
rect 11161 18037 11195 18071
rect 11805 18037 11839 18071
rect 17049 18037 17083 18071
rect 20453 18037 20487 18071
rect 2329 17833 2363 17867
rect 5273 17833 5307 17867
rect 6377 17833 6411 17867
rect 11253 17833 11287 17867
rect 13461 17833 13495 17867
rect 13921 17833 13955 17867
rect 17141 17833 17175 17867
rect 3985 17765 4019 17799
rect 16681 17765 16715 17799
rect 22477 17765 22511 17799
rect 22845 17765 22879 17799
rect 8585 17697 8619 17731
rect 9505 17697 9539 17731
rect 11713 17697 11747 17731
rect 11989 17697 12023 17731
rect 14933 17697 14967 17731
rect 15209 17697 15243 17731
rect 17693 17697 17727 17731
rect 18337 17697 18371 17731
rect 18889 17697 18923 17731
rect 22937 17697 22971 17731
rect 23949 17697 23983 17731
rect 1685 17629 1719 17663
rect 2789 17629 2823 17663
rect 4169 17629 4203 17663
rect 4629 17629 4663 17663
rect 5733 17629 5767 17663
rect 6837 17629 6871 17663
rect 7941 17629 7975 17663
rect 9137 17629 9171 17663
rect 19533 17629 19567 17663
rect 19993 17629 20027 17663
rect 20729 17629 20763 17663
rect 23765 17629 23799 17663
rect 24593 17629 24627 17663
rect 3433 17561 3467 17595
rect 9781 17561 9815 17595
rect 14289 17561 14323 17595
rect 17601 17561 17635 17595
rect 21005 17561 21039 17595
rect 23673 17561 23707 17595
rect 7481 17493 7515 17527
rect 8953 17493 8987 17527
rect 17509 17493 17543 17527
rect 23305 17493 23339 17527
rect 25237 17493 25271 17527
rect 2697 17289 2731 17323
rect 3801 17289 3835 17323
rect 6469 17289 6503 17323
rect 7665 17289 7699 17323
rect 8769 17289 8803 17323
rect 14749 17289 14783 17323
rect 20177 17289 20211 17323
rect 21281 17289 21315 17323
rect 1777 17221 1811 17255
rect 4905 17221 4939 17255
rect 9505 17221 9539 17255
rect 12817 17221 12851 17255
rect 15853 17221 15887 17255
rect 16497 17221 16531 17255
rect 17233 17221 17267 17255
rect 18705 17221 18739 17255
rect 2053 17153 2087 17187
rect 3157 17153 3191 17187
rect 4261 17153 4295 17187
rect 5365 17153 5399 17187
rect 7021 17153 7055 17187
rect 8125 17153 8159 17187
rect 9229 17153 9263 17187
rect 11897 17153 11931 17187
rect 14933 17153 14967 17187
rect 15761 17153 15795 17187
rect 18429 17153 18463 17187
rect 20637 17153 20671 17187
rect 22477 17153 22511 17187
rect 24685 17153 24719 17187
rect 12541 17085 12575 17119
rect 15945 17085 15979 17119
rect 17325 17085 17359 17119
rect 17417 17085 17451 17119
rect 18153 17085 18187 17119
rect 22753 17085 22787 17119
rect 24225 17085 24259 17119
rect 11253 17017 11287 17051
rect 12081 17017 12115 17051
rect 25329 17017 25363 17051
rect 6009 16949 6043 16983
rect 6745 16949 6779 16983
rect 10977 16949 11011 16983
rect 14289 16949 14323 16983
rect 15393 16949 15427 16983
rect 16865 16949 16899 16983
rect 17877 16949 17911 16983
rect 21557 16949 21591 16983
rect 22017 16949 22051 16983
rect 22109 16949 22143 16983
rect 4629 16745 4663 16779
rect 16037 16677 16071 16711
rect 9045 16609 9079 16643
rect 11253 16609 11287 16643
rect 11345 16609 11379 16643
rect 14289 16609 14323 16643
rect 14565 16609 14599 16643
rect 17141 16609 17175 16643
rect 17417 16609 17451 16643
rect 19441 16609 19475 16643
rect 22293 16609 22327 16643
rect 22569 16609 22603 16643
rect 1685 16541 1719 16575
rect 2789 16541 2823 16575
rect 3985 16541 4019 16575
rect 5273 16541 5307 16575
rect 5733 16541 5767 16575
rect 6377 16541 6411 16575
rect 6837 16541 6871 16575
rect 7941 16541 7975 16575
rect 9689 16541 9723 16575
rect 11989 16541 12023 16575
rect 16681 16541 16715 16575
rect 21833 16541 21867 16575
rect 24593 16541 24627 16575
rect 9137 16473 9171 16507
rect 12265 16473 12299 16507
rect 19717 16473 19751 16507
rect 2329 16405 2363 16439
rect 3433 16405 3467 16439
rect 5089 16405 5123 16439
rect 7481 16405 7515 16439
rect 8585 16405 8619 16439
rect 9413 16405 9447 16439
rect 10333 16405 10367 16439
rect 10793 16405 10827 16439
rect 11161 16405 11195 16439
rect 13737 16405 13771 16439
rect 16497 16405 16531 16439
rect 18889 16405 18923 16439
rect 21189 16405 21223 16439
rect 21649 16405 21683 16439
rect 24041 16405 24075 16439
rect 25237 16405 25271 16439
rect 1593 16201 1627 16235
rect 4905 16201 4939 16235
rect 6009 16201 6043 16235
rect 6561 16201 6595 16235
rect 7849 16201 7883 16235
rect 11161 16201 11195 16235
rect 13461 16201 13495 16235
rect 15393 16201 15427 16235
rect 18337 16201 18371 16235
rect 19625 16201 19659 16235
rect 20821 16201 20855 16235
rect 23857 16201 23891 16235
rect 15025 16133 15059 16167
rect 15853 16133 15887 16167
rect 22385 16133 22419 16167
rect 23029 16133 23063 16167
rect 2053 16065 2087 16099
rect 3157 16065 3191 16099
rect 4261 16065 4295 16099
rect 5365 16065 5399 16099
rect 6745 16065 6779 16099
rect 7205 16065 7239 16099
rect 8309 16065 8343 16099
rect 8953 16065 8987 16099
rect 9413 16065 9447 16099
rect 10517 16065 10551 16099
rect 11713 16065 11747 16099
rect 14289 16065 14323 16099
rect 15761 16065 15795 16099
rect 17049 16065 17083 16099
rect 20269 16065 20303 16099
rect 21465 16065 21499 16099
rect 22477 16065 22511 16099
rect 23765 16065 23799 16099
rect 24593 16065 24627 16099
rect 1777 15997 1811 16031
rect 11989 15997 12023 16031
rect 14381 15997 14415 16031
rect 14565 15997 14599 16031
rect 15945 15997 15979 16031
rect 19717 15997 19751 16031
rect 19809 15997 19843 16031
rect 20913 15997 20947 16031
rect 21097 15997 21131 16031
rect 22569 15997 22603 16031
rect 24041 15997 24075 16031
rect 2697 15929 2731 15963
rect 19257 15929 19291 15963
rect 20453 15929 20487 15963
rect 3801 15861 3835 15895
rect 10057 15861 10091 15895
rect 13921 15861 13955 15895
rect 16405 15861 16439 15895
rect 16773 15861 16807 15895
rect 22017 15861 22051 15895
rect 23397 15861 23431 15895
rect 25237 15861 25271 15895
rect 3985 15657 4019 15691
rect 6377 15657 6411 15691
rect 10590 15657 10624 15691
rect 13829 15657 13863 15691
rect 16037 15657 16071 15691
rect 16589 15657 16623 15691
rect 18705 15657 18739 15691
rect 23765 15657 23799 15691
rect 2145 15589 2179 15623
rect 1593 15521 1627 15555
rect 10333 15521 10367 15555
rect 13185 15521 13219 15555
rect 14289 15521 14323 15555
rect 17233 15521 17267 15555
rect 19349 15521 19383 15555
rect 20085 15521 20119 15555
rect 20177 15521 20211 15555
rect 21281 15521 21315 15555
rect 21373 15521 21407 15555
rect 2605 15453 2639 15487
rect 2881 15453 2915 15487
rect 4169 15453 4203 15487
rect 4629 15453 4663 15487
rect 5733 15453 5767 15487
rect 6837 15453 6871 15487
rect 7941 15453 7975 15487
rect 9229 15453 9263 15487
rect 13737 15453 13771 15487
rect 16957 15453 16991 15487
rect 20729 15453 20763 15487
rect 21189 15453 21223 15487
rect 22017 15453 22051 15487
rect 23121 15453 23155 15487
rect 24593 15453 24627 15487
rect 1961 15385 1995 15419
rect 7481 15385 7515 15419
rect 13001 15385 13035 15419
rect 14565 15385 14599 15419
rect 19441 15385 19475 15419
rect 19993 15385 20027 15419
rect 5273 15317 5307 15351
rect 8585 15317 8619 15351
rect 9873 15317 9907 15351
rect 12081 15317 12115 15351
rect 12541 15317 12575 15351
rect 12909 15317 12943 15351
rect 16313 15317 16347 15351
rect 19073 15317 19107 15351
rect 19625 15317 19659 15351
rect 20821 15317 20855 15351
rect 22661 15317 22695 15351
rect 24133 15317 24167 15351
rect 25237 15317 25271 15351
rect 4905 15113 4939 15147
rect 6009 15113 6043 15147
rect 7849 15113 7883 15147
rect 14473 15113 14507 15147
rect 15577 15113 15611 15147
rect 11161 15045 11195 15079
rect 12173 15045 12207 15079
rect 16129 15045 16163 15079
rect 19625 15045 19659 15079
rect 21465 15045 21499 15079
rect 23029 15045 23063 15079
rect 3157 14977 3191 15011
rect 4261 14977 4295 15011
rect 5365 14977 5399 15011
rect 6745 14977 6779 15011
rect 7205 14977 7239 15011
rect 8309 14977 8343 15011
rect 9413 14977 9447 15011
rect 10517 14977 10551 15011
rect 11805 14977 11839 15011
rect 14933 14977 14967 15011
rect 22109 14977 22143 15011
rect 22753 14977 22787 15011
rect 25145 14977 25179 15011
rect 1869 14909 1903 14943
rect 2145 14909 2179 14943
rect 12725 14909 12759 14943
rect 13001 14909 13035 14943
rect 16865 14909 16899 14943
rect 17141 14909 17175 14943
rect 19349 14909 19383 14943
rect 24501 14909 24535 14943
rect 16313 14841 16347 14875
rect 19073 14841 19107 14875
rect 21097 14841 21131 14875
rect 22293 14841 22327 14875
rect 3801 14773 3835 14807
rect 6561 14773 6595 14807
rect 8953 14773 8987 14807
rect 10057 14773 10091 14807
rect 18613 14773 18647 14807
rect 21557 14773 21591 14807
rect 25237 14773 25271 14807
rect 7481 14569 7515 14603
rect 8585 14569 8619 14603
rect 9045 14569 9079 14603
rect 9229 14569 9263 14603
rect 12633 14569 12667 14603
rect 16037 14569 16071 14603
rect 18245 14569 18279 14603
rect 18705 14569 18739 14603
rect 22293 14569 22327 14603
rect 12357 14501 12391 14535
rect 6377 14433 6411 14467
rect 10609 14433 10643 14467
rect 10885 14433 10919 14467
rect 14289 14433 14323 14467
rect 16497 14433 16531 14467
rect 20085 14433 20119 14467
rect 23489 14433 23523 14467
rect 23581 14433 23615 14467
rect 25145 14433 25179 14467
rect 2145 14365 2179 14399
rect 2605 14365 2639 14399
rect 2881 14365 2915 14399
rect 4169 14365 4203 14399
rect 4629 14365 4663 14399
rect 5273 14365 5307 14399
rect 5733 14365 5767 14399
rect 6837 14365 6871 14399
rect 7941 14365 7975 14399
rect 9505 14365 9539 14399
rect 13093 14365 13127 14399
rect 18889 14365 18923 14399
rect 19901 14365 19935 14399
rect 25053 14365 25087 14399
rect 13737 14297 13771 14331
rect 14565 14297 14599 14331
rect 16773 14297 16807 14331
rect 20821 14297 20855 14331
rect 24041 14297 24075 14331
rect 1961 14229 1995 14263
rect 3985 14229 4019 14263
rect 10149 14229 10183 14263
rect 19441 14229 19475 14263
rect 19809 14229 19843 14263
rect 20453 14229 20487 14263
rect 23029 14229 23063 14263
rect 23397 14229 23431 14263
rect 24593 14229 24627 14263
rect 24961 14229 24995 14263
rect 2789 14025 2823 14059
rect 2881 14025 2915 14059
rect 4721 14025 4755 14059
rect 6561 14025 6595 14059
rect 11161 14025 11195 14059
rect 13185 14025 13219 14059
rect 17509 14025 17543 14059
rect 17877 14025 17911 14059
rect 19533 14025 19567 14059
rect 20361 14025 20395 14059
rect 20729 14025 20763 14059
rect 24041 14025 24075 14059
rect 25145 14025 25179 14059
rect 3157 13957 3191 13991
rect 18245 13957 18279 13991
rect 21189 13957 21223 13991
rect 1593 13889 1627 13923
rect 1869 13889 1903 13923
rect 3433 13889 3467 13923
rect 4905 13889 4939 13923
rect 5365 13889 5399 13923
rect 7205 13889 7239 13923
rect 8309 13889 8343 13923
rect 9413 13889 9447 13923
rect 11897 13889 11931 13923
rect 12081 13889 12115 13923
rect 12541 13889 12575 13923
rect 13645 13889 13679 13923
rect 15853 13889 15887 13923
rect 16865 13889 16899 13923
rect 21097 13889 21131 13923
rect 22293 13889 22327 13923
rect 24501 13889 24535 13923
rect 3709 13821 3743 13855
rect 6009 13821 6043 13855
rect 7849 13821 7883 13855
rect 8953 13821 8987 13855
rect 9689 13821 9723 13855
rect 15393 13821 15427 13855
rect 16037 13821 16071 13855
rect 20545 13821 20579 13855
rect 21281 13821 21315 13855
rect 21925 13821 21959 13855
rect 25513 13821 25547 13855
rect 13908 13685 13942 13719
rect 22556 13685 22590 13719
rect 2329 13481 2363 13515
rect 3249 13481 3283 13515
rect 5457 13481 5491 13515
rect 8585 13481 8619 13515
rect 8953 13481 8987 13515
rect 9229 13481 9263 13515
rect 10793 13481 10827 13515
rect 15025 13481 15059 13515
rect 23673 13481 23707 13515
rect 24041 13481 24075 13515
rect 25237 13481 25271 13515
rect 2789 13413 2823 13447
rect 13461 13413 13495 13447
rect 17969 13413 18003 13447
rect 3985 13345 4019 13379
rect 4261 13345 4295 13379
rect 11713 13345 11747 13379
rect 15669 13345 15703 13379
rect 18521 13345 18555 13379
rect 19717 13345 19751 13379
rect 21925 13345 21959 13379
rect 22201 13345 22235 13379
rect 1685 13277 1719 13311
rect 3433 13277 3467 13311
rect 5273 13277 5307 13311
rect 5733 13277 5767 13311
rect 6837 13277 6871 13311
rect 7941 13277 7975 13311
rect 9505 13277 9539 13311
rect 14381 13277 14415 13311
rect 24593 13277 24627 13311
rect 2973 13209 3007 13243
rect 7481 13209 7515 13243
rect 11989 13209 12023 13243
rect 15945 13209 15979 13243
rect 18429 13209 18463 13243
rect 19993 13209 20027 13243
rect 24225 13209 24259 13243
rect 6377 13141 6411 13175
rect 15393 13141 15427 13175
rect 17417 13141 17451 13175
rect 18337 13141 18371 13175
rect 18981 13141 19015 13175
rect 19441 13141 19475 13175
rect 21465 13141 21499 13175
rect 2053 12937 2087 12971
rect 4721 12937 4755 12971
rect 4997 12937 5031 12971
rect 5089 12937 5123 12971
rect 5825 12937 5859 12971
rect 6561 12937 6595 12971
rect 10057 12937 10091 12971
rect 11161 12937 11195 12971
rect 15025 12937 15059 12971
rect 16313 12937 16347 12971
rect 19441 12937 19475 12971
rect 20729 12937 20763 12971
rect 21557 12937 21591 12971
rect 21925 12937 21959 12971
rect 24133 12937 24167 12971
rect 4445 12869 4479 12903
rect 12817 12869 12851 12903
rect 13553 12869 13587 12903
rect 1961 12801 1995 12835
rect 3525 12801 3559 12835
rect 4629 12801 4663 12835
rect 6745 12801 6779 12835
rect 7205 12801 7239 12835
rect 8677 12801 8711 12835
rect 9137 12801 9171 12835
rect 9413 12801 9447 12835
rect 10517 12801 10551 12835
rect 12173 12801 12207 12835
rect 15669 12801 15703 12835
rect 16865 12801 16899 12835
rect 20637 12801 20671 12835
rect 21465 12801 21499 12835
rect 22385 12801 22419 12835
rect 24593 12801 24627 12835
rect 2605 12733 2639 12767
rect 3249 12733 3283 12767
rect 7481 12733 7515 12767
rect 13277 12733 13311 12767
rect 17141 12733 17175 12767
rect 18613 12733 18647 12767
rect 19533 12733 19567 12767
rect 19625 12733 19659 12767
rect 20913 12733 20947 12767
rect 8493 12665 8527 12699
rect 19073 12665 19107 12699
rect 15301 12597 15335 12631
rect 18889 12597 18923 12631
rect 20269 12597 20303 12631
rect 22642 12597 22676 12631
rect 25237 12597 25271 12631
rect 2605 12393 2639 12427
rect 9137 12393 9171 12427
rect 12633 12393 12667 12427
rect 18521 12393 18555 12427
rect 21189 12393 21223 12427
rect 23765 12393 23799 12427
rect 14933 12325 14967 12359
rect 15301 12325 15335 12359
rect 3249 12257 3283 12291
rect 4997 12257 5031 12291
rect 6653 12257 6687 12291
rect 6929 12257 6963 12291
rect 19441 12257 19475 12291
rect 19717 12257 19751 12291
rect 21557 12257 21591 12291
rect 1869 12189 1903 12223
rect 2789 12189 2823 12223
rect 4261 12189 4295 12223
rect 4721 12189 4755 12223
rect 6193 12189 6227 12223
rect 7941 12189 7975 12223
rect 9321 12189 9355 12223
rect 9781 12189 9815 12223
rect 10885 12189 10919 12223
rect 11989 12189 12023 12223
rect 13093 12189 13127 12223
rect 14289 12189 14323 12223
rect 15669 12189 15703 12223
rect 17877 12189 17911 12223
rect 18797 12189 18831 12223
rect 22017 12189 22051 12223
rect 24133 12189 24167 12223
rect 24593 12189 24627 12223
rect 10425 12121 10459 12155
rect 19073 12121 19107 12155
rect 22293 12121 22327 12155
rect 4077 12053 4111 12087
rect 6009 12053 6043 12087
rect 8585 12053 8619 12087
rect 11529 12053 11563 12087
rect 13737 12053 13771 12087
rect 16957 12053 16991 12087
rect 21649 12053 21683 12087
rect 25237 12053 25271 12087
rect 3157 11849 3191 11883
rect 9873 11849 9907 11883
rect 10977 11849 11011 11883
rect 11253 11849 11287 11883
rect 13461 11849 13495 11883
rect 14565 11849 14599 11883
rect 15025 11849 15059 11883
rect 16313 11849 16347 11883
rect 21557 11849 21591 11883
rect 12357 11781 12391 11815
rect 23305 11781 23339 11815
rect 25145 11781 25179 11815
rect 1593 11713 1627 11747
rect 2053 11713 2087 11747
rect 2697 11713 2731 11747
rect 3801 11713 3835 11747
rect 5181 11713 5215 11747
rect 6561 11713 6595 11747
rect 7941 11713 7975 11747
rect 9229 11713 9263 11747
rect 10333 11713 10367 11747
rect 11701 11713 11735 11747
rect 12817 11713 12851 11747
rect 13921 11713 13955 11747
rect 15669 11713 15703 11747
rect 17049 11713 17083 11747
rect 19349 11713 19383 11747
rect 22293 11713 22327 11747
rect 23949 11713 23983 11747
rect 4077 11645 4111 11679
rect 5457 11645 5491 11679
rect 6837 11645 6871 11679
rect 16773 11645 16807 11679
rect 17325 11645 17359 11679
rect 19625 11645 19659 11679
rect 1869 11577 1903 11611
rect 2513 11509 2547 11543
rect 8585 11509 8619 11543
rect 8861 11509 8895 11543
rect 18797 11509 18831 11543
rect 21097 11509 21131 11543
rect 1869 11305 1903 11339
rect 2789 11305 2823 11339
rect 3801 11305 3835 11339
rect 7849 11305 7883 11339
rect 8401 11305 8435 11339
rect 10333 11305 10367 11339
rect 13185 11305 13219 11339
rect 21189 11305 21223 11339
rect 5733 11237 5767 11271
rect 10793 11237 10827 11271
rect 18797 11237 18831 11271
rect 4537 11169 4571 11203
rect 4813 11169 4847 11203
rect 6653 11169 6687 11203
rect 9137 11169 9171 11203
rect 10517 11169 10551 11203
rect 15669 11169 15703 11203
rect 17417 11169 17451 11203
rect 22201 11169 22235 11203
rect 23857 11169 23891 11203
rect 2237 11101 2271 11135
rect 3433 11101 3467 11135
rect 6377 11101 6411 11135
rect 7757 11101 7791 11135
rect 8585 11101 8619 11135
rect 9413 11101 9447 11135
rect 10977 11101 11011 11135
rect 11437 11101 11471 11135
rect 12541 11101 12575 11135
rect 13461 11101 13495 11135
rect 14565 11101 14599 11135
rect 17877 11101 17911 11135
rect 19441 11101 19475 11135
rect 20545 11101 20579 11135
rect 21741 11101 21775 11135
rect 21925 11101 21959 11135
rect 22661 11101 22695 11135
rect 24593 11101 24627 11135
rect 2421 11033 2455 11067
rect 12081 11033 12115 11067
rect 15209 11033 15243 11067
rect 15945 11033 15979 11067
rect 18981 11033 19015 11067
rect 20085 11033 20119 11067
rect 25237 11033 25271 11067
rect 3249 10965 3283 10999
rect 18521 10965 18555 10999
rect 3341 10761 3375 10795
rect 7113 10761 7147 10795
rect 7757 10761 7791 10795
rect 8401 10761 8435 10795
rect 13553 10761 13587 10795
rect 15761 10761 15795 10795
rect 18705 10761 18739 10795
rect 20913 10761 20947 10795
rect 21465 10761 21499 10795
rect 3801 10693 3835 10727
rect 3985 10693 4019 10727
rect 19809 10693 19843 10727
rect 25145 10693 25179 10727
rect 2145 10625 2179 10659
rect 6745 10625 6779 10659
rect 7297 10625 7331 10659
rect 7941 10625 7975 10659
rect 8585 10625 8619 10659
rect 9229 10625 9263 10659
rect 9873 10625 9907 10659
rect 10609 10625 10643 10659
rect 11805 10625 11839 10659
rect 12909 10625 12943 10659
rect 14013 10625 14047 10659
rect 15117 10625 15151 10659
rect 16865 10625 16899 10659
rect 18061 10625 18095 10659
rect 19165 10625 19199 10659
rect 20269 10625 20303 10659
rect 22109 10625 22143 10659
rect 23949 10625 23983 10659
rect 2421 10557 2455 10591
rect 4445 10557 4479 10591
rect 4721 10557 4755 10591
rect 5825 10557 5859 10591
rect 10333 10557 10367 10591
rect 23305 10557 23339 10591
rect 5641 10489 5675 10523
rect 9689 10489 9723 10523
rect 21557 10489 21591 10523
rect 9045 10421 9079 10455
rect 12449 10421 12483 10455
rect 14657 10421 14691 10455
rect 16037 10421 16071 10455
rect 17509 10421 17543 10455
rect 21281 10421 21315 10455
rect 6745 10217 6779 10251
rect 9137 10217 9171 10251
rect 11713 10217 11747 10251
rect 16497 10217 16531 10251
rect 18981 10217 19015 10251
rect 19349 10217 19383 10251
rect 20361 10217 20395 10251
rect 24225 10217 24259 10251
rect 2329 10149 2363 10183
rect 5365 10149 5399 10183
rect 5917 10149 5951 10183
rect 8309 10149 8343 10183
rect 12633 10149 12667 10183
rect 18705 10149 18739 10183
rect 21005 10149 21039 10183
rect 24593 10149 24627 10183
rect 4077 10081 4111 10115
rect 21281 10081 21315 10115
rect 25053 10081 25087 10115
rect 25145 10081 25179 10115
rect 2145 10013 2179 10047
rect 4353 10013 4387 10047
rect 5641 10013 5675 10047
rect 6101 10013 6135 10047
rect 8493 10013 8527 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 10701 10013 10735 10047
rect 11989 10013 12023 10047
rect 13093 10013 13127 10047
rect 14105 10013 14139 10047
rect 14749 10013 14783 10047
rect 15853 10013 15887 10047
rect 16957 10013 16991 10047
rect 17601 10013 17635 10047
rect 18061 10013 18095 10047
rect 19717 10013 19751 10047
rect 20729 10013 20763 10047
rect 2789 9945 2823 9979
rect 6653 9945 6687 9979
rect 21557 9945 21591 9979
rect 23673 9945 23707 9979
rect 7665 9877 7699 9911
rect 11345 9877 11379 9911
rect 13737 9877 13771 9911
rect 15393 9877 15427 9911
rect 23029 9877 23063 9911
rect 23765 9877 23799 9911
rect 24409 9877 24443 9911
rect 24961 9877 24995 9911
rect 20453 9673 20487 9707
rect 4721 9605 4755 9639
rect 5181 9605 5215 9639
rect 15209 9605 15243 9639
rect 18797 9605 18831 9639
rect 23305 9605 23339 9639
rect 1869 9537 1903 9571
rect 2329 9537 2363 9571
rect 2973 9537 3007 9571
rect 3617 9537 3651 9571
rect 4261 9537 4295 9571
rect 5917 9537 5951 9571
rect 7205 9537 7239 9571
rect 7757 9537 7791 9571
rect 9321 9537 9355 9571
rect 10609 9537 10643 9571
rect 11897 9537 11931 9571
rect 12357 9537 12391 9571
rect 13461 9537 13495 9571
rect 14473 9537 14507 9571
rect 14565 9537 14599 9571
rect 15669 9537 15703 9571
rect 17049 9537 17083 9571
rect 18153 9537 18187 9571
rect 19809 9537 19843 9571
rect 21005 9537 21039 9571
rect 22201 9537 22235 9571
rect 23949 9537 23983 9571
rect 8033 9469 8067 9503
rect 9045 9469 9079 9503
rect 10333 9469 10367 9503
rect 24777 9469 24811 9503
rect 2145 9401 2179 9435
rect 2789 9401 2823 9435
rect 3433 9401 3467 9435
rect 5733 9401 5767 9435
rect 11713 9401 11747 9435
rect 14105 9401 14139 9435
rect 21189 9401 21223 9435
rect 4077 9333 4111 9367
rect 5365 9333 5399 9367
rect 7021 9333 7055 9367
rect 13001 9333 13035 9367
rect 16313 9333 16347 9367
rect 16681 9333 16715 9367
rect 17693 9333 17727 9367
rect 19073 9333 19107 9367
rect 21557 9333 21591 9367
rect 1593 9129 1627 9163
rect 1961 9129 1995 9163
rect 3249 9129 3283 9163
rect 5825 9129 5859 9163
rect 7297 9129 7331 9163
rect 7849 9129 7883 9163
rect 8953 9129 8987 9163
rect 12357 9129 12391 9163
rect 16865 9129 16899 9163
rect 17969 9129 18003 9163
rect 21189 9129 21223 9163
rect 25237 9129 25271 9163
rect 5181 9061 5215 9095
rect 9321 8993 9355 9027
rect 10057 8993 10091 9027
rect 12081 8993 12115 9027
rect 2145 8925 2179 8959
rect 2789 8925 2823 8959
rect 3433 8925 3467 8959
rect 4169 8925 4203 8959
rect 4905 8925 4939 8959
rect 6009 8925 6043 8959
rect 6745 8925 6779 8959
rect 7481 8925 7515 8959
rect 8585 8925 8619 8959
rect 13093 8925 13127 8959
rect 14381 8925 14415 8959
rect 15117 8925 15151 8959
rect 16221 8925 16255 8959
rect 17325 8925 17359 8959
rect 18429 8925 18463 8959
rect 19441 8925 19475 8959
rect 20545 8925 20579 8959
rect 22661 8925 22695 8959
rect 24593 8925 24627 8959
rect 8033 8857 8067 8891
rect 10333 8857 10367 8891
rect 18705 8857 18739 8891
rect 21741 8857 21775 8891
rect 22201 8857 22235 8891
rect 23857 8857 23891 8891
rect 2605 8789 2639 8823
rect 3985 8789 4019 8823
rect 4721 8789 4755 8823
rect 6561 8789 6595 8823
rect 8401 8789 8435 8823
rect 13737 8789 13771 8823
rect 15761 8789 15795 8823
rect 20085 8789 20119 8823
rect 21833 8789 21867 8823
rect 1961 8585 1995 8619
rect 2605 8585 2639 8619
rect 3249 8585 3283 8619
rect 4445 8585 4479 8619
rect 6837 8585 6871 8619
rect 8677 8585 8711 8619
rect 9689 8585 9723 8619
rect 15209 8585 15243 8619
rect 18613 8585 18647 8619
rect 20821 8585 20855 8619
rect 21281 8517 21315 8551
rect 25145 8517 25179 8551
rect 4169 8449 4203 8483
rect 4629 8449 4663 8483
rect 8861 8449 8895 8483
rect 9137 8449 9171 8483
rect 9413 8449 9447 8483
rect 9873 8449 9907 8483
rect 11989 8449 12023 8483
rect 13461 8449 13495 8483
rect 14565 8449 14599 8483
rect 15669 8449 15703 8483
rect 16865 8449 16899 8483
rect 17969 8449 18003 8483
rect 19073 8449 19107 8483
rect 20177 8449 20211 8483
rect 22109 8449 22143 8483
rect 23949 8449 23983 8483
rect 10333 8381 10367 8415
rect 10609 8381 10643 8415
rect 11713 8381 11747 8415
rect 16313 8381 16347 8415
rect 17509 8381 17543 8415
rect 23305 8381 23339 8415
rect 3985 8313 4019 8347
rect 14105 8313 14139 8347
rect 19717 8245 19751 8279
rect 2145 8041 2179 8075
rect 2881 8041 2915 8075
rect 3617 8041 3651 8075
rect 10517 8041 10551 8075
rect 12357 8041 12391 8075
rect 12909 8041 12943 8075
rect 14197 8041 14231 8075
rect 17325 8041 17359 8075
rect 18429 8041 18463 8075
rect 20085 8041 20119 8075
rect 2605 7973 2639 8007
rect 15117 7973 15151 8007
rect 11253 7905 11287 7939
rect 20821 7905 20855 7939
rect 2329 7837 2363 7871
rect 9873 7837 9907 7871
rect 10977 7837 11011 7871
rect 12541 7837 12575 7871
rect 13461 7837 13495 7871
rect 13737 7837 13771 7871
rect 14473 7837 14507 7871
rect 15577 7837 15611 7871
rect 16681 7837 16715 7871
rect 17785 7837 17819 7871
rect 19441 7837 19475 7871
rect 20637 7837 20671 7871
rect 21557 7837 21591 7871
rect 22845 7837 22879 7871
rect 24593 7837 24627 7871
rect 23857 7769 23891 7803
rect 13553 7701 13587 7735
rect 16221 7701 16255 7735
rect 22201 7701 22235 7735
rect 25237 7701 25271 7735
rect 10977 7497 11011 7531
rect 11805 7497 11839 7531
rect 15025 7497 15059 7531
rect 16129 7497 16163 7531
rect 16405 7497 16439 7531
rect 18797 7497 18831 7531
rect 19901 7429 19935 7463
rect 10517 7361 10551 7395
rect 10885 7361 10919 7395
rect 11161 7361 11195 7395
rect 12725 7361 12759 7395
rect 14013 7361 14047 7395
rect 15209 7361 15243 7395
rect 15853 7361 15887 7395
rect 18153 7361 18187 7395
rect 19257 7361 19291 7395
rect 20361 7361 20395 7395
rect 21281 7361 21315 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 12449 7293 12483 7327
rect 13737 7293 13771 7327
rect 16865 7293 16899 7327
rect 17141 7293 17175 7327
rect 23305 7293 23339 7327
rect 24777 7293 24811 7327
rect 10333 7157 10367 7191
rect 15669 7157 15703 7191
rect 21005 7157 21039 7191
rect 12679 6953 12713 6987
rect 18889 6953 18923 6987
rect 16773 6885 16807 6919
rect 19257 6885 19291 6919
rect 20361 6817 20395 6851
rect 11345 6749 11379 6783
rect 12449 6749 12483 6783
rect 14933 6749 14967 6783
rect 15577 6749 15611 6783
rect 16221 6749 16255 6783
rect 16589 6749 16623 6783
rect 17141 6749 17175 6783
rect 18245 6749 18279 6783
rect 19717 6749 19751 6783
rect 20821 6749 20855 6783
rect 22109 6749 22143 6783
rect 22661 6749 22695 6783
rect 24593 6749 24627 6783
rect 17785 6681 17819 6715
rect 23857 6681 23891 6715
rect 11161 6613 11195 6647
rect 11713 6613 11747 6647
rect 11805 6613 11839 6647
rect 14473 6613 14507 6647
rect 14749 6613 14783 6647
rect 15393 6613 15427 6647
rect 16037 6613 16071 6647
rect 21465 6613 21499 6647
rect 21925 6613 21959 6647
rect 25237 6613 25271 6647
rect 9321 6409 9355 6443
rect 11529 6409 11563 6443
rect 12909 6409 12943 6443
rect 15485 6409 15519 6443
rect 16037 6409 16071 6443
rect 16129 6409 16163 6443
rect 16957 6409 16991 6443
rect 22661 6409 22695 6443
rect 19165 6341 19199 6375
rect 19901 6341 19935 6375
rect 8677 6273 8711 6307
rect 13737 6273 13771 6307
rect 14197 6273 14231 6307
rect 15669 6273 15703 6307
rect 17417 6273 17451 6307
rect 18061 6273 18095 6307
rect 18521 6273 18555 6307
rect 19717 6273 19751 6307
rect 20821 6273 20855 6307
rect 22017 6273 22051 6307
rect 23949 6273 23983 6307
rect 12173 6205 12207 6239
rect 12265 6205 12299 6239
rect 14473 6205 14507 6239
rect 20177 6205 20211 6239
rect 20545 6205 20579 6239
rect 24777 6205 24811 6239
rect 23581 6137 23615 6171
rect 13553 6069 13587 6103
rect 16773 6069 16807 6103
rect 22937 6069 22971 6103
rect 16865 5865 16899 5899
rect 20269 5729 20303 5763
rect 21373 5729 21407 5763
rect 21649 5729 21683 5763
rect 14289 5661 14323 5695
rect 14565 5661 14599 5695
rect 15577 5661 15611 5695
rect 15853 5661 15887 5695
rect 17049 5661 17083 5695
rect 18245 5661 18279 5695
rect 19625 5661 19659 5695
rect 20913 5661 20947 5695
rect 22661 5661 22695 5695
rect 24593 5661 24627 5695
rect 17601 5593 17635 5627
rect 17785 5593 17819 5627
rect 18889 5593 18923 5627
rect 23857 5593 23891 5627
rect 12909 5525 12943 5559
rect 13553 5525 13587 5559
rect 19257 5525 19291 5559
rect 20729 5525 20763 5559
rect 25237 5525 25271 5559
rect 13553 5321 13587 5355
rect 14013 5321 14047 5355
rect 15577 5321 15611 5355
rect 16865 5321 16899 5355
rect 18245 5321 18279 5355
rect 23305 5253 23339 5287
rect 13737 5185 13771 5219
rect 15761 5185 15795 5219
rect 17049 5185 17083 5219
rect 17693 5185 17727 5219
rect 18613 5185 18647 5219
rect 19717 5185 19751 5219
rect 20361 5185 20395 5219
rect 20821 5185 20855 5219
rect 22293 5185 22327 5219
rect 23949 5185 23983 5219
rect 14933 5117 14967 5151
rect 16129 5117 16163 5151
rect 24685 5117 24719 5151
rect 16497 5049 16531 5083
rect 17509 5049 17543 5083
rect 17969 4981 18003 5015
rect 19257 4981 19291 5015
rect 21465 4981 21499 5015
rect 8585 4777 8619 4811
rect 16037 4777 16071 4811
rect 16681 4777 16715 4811
rect 17141 4777 17175 4811
rect 20361 4777 20395 4811
rect 25237 4777 25271 4811
rect 19349 4709 19383 4743
rect 14749 4641 14783 4675
rect 7941 4573 7975 4607
rect 15025 4573 15059 4607
rect 16221 4573 16255 4607
rect 16865 4573 16899 4607
rect 17325 4573 17359 4607
rect 18153 4573 18187 4607
rect 19717 4573 19751 4607
rect 21005 4573 21039 4607
rect 22661 4573 22695 4607
rect 24593 4573 24627 4607
rect 18705 4505 18739 4539
rect 18889 4505 18923 4539
rect 22017 4505 22051 4539
rect 23857 4505 23891 4539
rect 17969 4437 18003 4471
rect 16313 4233 16347 4267
rect 6837 4097 6871 4131
rect 17049 4097 17083 4131
rect 18337 4097 18371 4131
rect 18981 4097 19015 4131
rect 19625 4097 19659 4131
rect 20085 4097 20119 4131
rect 22109 4097 22143 4131
rect 23949 4097 23983 4131
rect 17417 4029 17451 4063
rect 17509 4029 17543 4063
rect 21281 4029 21315 4063
rect 23305 4029 23339 4063
rect 24777 4029 24811 4063
rect 16865 3961 16899 3995
rect 7481 3893 7515 3927
rect 18153 3893 18187 3927
rect 18797 3893 18831 3927
rect 19441 3893 19475 3927
rect 8217 3689 8251 3723
rect 16405 3689 16439 3723
rect 17417 3689 17451 3723
rect 18705 3689 18739 3723
rect 20361 3689 20395 3723
rect 25237 3689 25271 3723
rect 16773 3553 16807 3587
rect 6469 3485 6503 3519
rect 7573 3485 7607 3519
rect 17601 3485 17635 3519
rect 18245 3485 18279 3519
rect 18889 3485 18923 3519
rect 19717 3485 19751 3519
rect 21005 3485 21039 3519
rect 22661 3485 22695 3519
rect 24593 3485 24627 3519
rect 19441 3417 19475 3451
rect 22017 3417 22051 3451
rect 23857 3417 23891 3451
rect 7113 3349 7147 3383
rect 18061 3349 18095 3383
rect 9137 3145 9171 3179
rect 16865 3145 16899 3179
rect 16957 3145 16991 3179
rect 16497 3077 16531 3111
rect 19441 3077 19475 3111
rect 23305 3077 23339 3111
rect 7389 3009 7423 3043
rect 8493 3009 8527 3043
rect 17785 3009 17819 3043
rect 18429 3009 18463 3043
rect 20269 3009 20303 3043
rect 22109 3009 22143 3043
rect 24133 3009 24167 3043
rect 21281 2941 21315 2975
rect 24593 2941 24627 2975
rect 17601 2873 17635 2907
rect 8033 2805 8067 2839
rect 6745 2601 6779 2635
rect 8677 2601 8711 2635
rect 9781 2601 9815 2635
rect 17601 2601 17635 2635
rect 18889 2601 18923 2635
rect 22017 2601 22051 2635
rect 25237 2601 25271 2635
rect 16957 2533 16991 2567
rect 8033 2465 8067 2499
rect 18245 2465 18279 2499
rect 21281 2465 21315 2499
rect 5365 2397 5399 2431
rect 6929 2397 6963 2431
rect 7389 2397 7423 2431
rect 9137 2397 9171 2431
rect 17141 2397 17175 2431
rect 17785 2397 17819 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 24593 2397 24627 2431
rect 6009 2329 6043 2363
rect 23857 2329 23891 2363
rect 16497 2261 16531 2295
rect 19441 2261 19475 2295
<< metal1 >>
rect 1026 26324 1032 26376
rect 1084 26364 1090 26376
rect 22554 26364 22560 26376
rect 1084 26336 22560 26364
rect 1084 26324 1090 26336
rect 22554 26324 22560 26336
rect 22612 26324 22618 26376
rect 2130 26256 2136 26308
rect 2188 26296 2194 26308
rect 22186 26296 22192 26308
rect 2188 26268 22192 26296
rect 2188 26256 2194 26268
rect 22186 26256 22192 26268
rect 22244 26256 22250 26308
rect 5442 26188 5448 26240
rect 5500 26228 5506 26240
rect 21266 26228 21272 26240
rect 5500 26200 21272 26228
rect 5500 26188 5506 26200
rect 21266 26188 21272 26200
rect 21324 26188 21330 26240
rect 1578 26120 1584 26172
rect 1636 26160 1642 26172
rect 16666 26160 16672 26172
rect 1636 26132 16672 26160
rect 1636 26120 1642 26132
rect 16666 26120 16672 26132
rect 16724 26160 16730 26172
rect 17310 26160 17316 26172
rect 16724 26132 17316 26160
rect 16724 26120 16730 26132
rect 17310 26120 17316 26132
rect 17368 26120 17374 26172
rect 10962 25916 10968 25968
rect 11020 25956 11026 25968
rect 14182 25956 14188 25968
rect 11020 25928 14188 25956
rect 11020 25916 11026 25928
rect 14182 25916 14188 25928
rect 14240 25916 14246 25968
rect 1854 25848 1860 25900
rect 1912 25888 1918 25900
rect 13722 25888 13728 25900
rect 1912 25860 13728 25888
rect 1912 25848 1918 25860
rect 13722 25848 13728 25860
rect 13780 25848 13786 25900
rect 3418 25780 3424 25832
rect 3476 25820 3482 25832
rect 21726 25820 21732 25832
rect 3476 25792 21732 25820
rect 3476 25780 3482 25792
rect 21726 25780 21732 25792
rect 21784 25780 21790 25832
rect 566 25712 572 25764
rect 624 25752 630 25764
rect 20898 25752 20904 25764
rect 624 25724 20904 25752
rect 624 25712 630 25724
rect 20898 25712 20904 25724
rect 20956 25712 20962 25764
rect 2406 25644 2412 25696
rect 2464 25684 2470 25696
rect 15838 25684 15844 25696
rect 2464 25656 15844 25684
rect 2464 25644 2470 25656
rect 15838 25644 15844 25656
rect 15896 25644 15902 25696
rect 2590 25576 2596 25628
rect 2648 25616 2654 25628
rect 20530 25616 20536 25628
rect 2648 25588 20536 25616
rect 2648 25576 2654 25588
rect 20530 25576 20536 25588
rect 20588 25576 20594 25628
rect 7282 25508 7288 25560
rect 7340 25548 7346 25560
rect 22002 25548 22008 25560
rect 7340 25520 22008 25548
rect 7340 25508 7346 25520
rect 22002 25508 22008 25520
rect 22060 25508 22066 25560
rect 4522 25440 4528 25492
rect 4580 25480 4586 25492
rect 24210 25480 24216 25492
rect 4580 25452 24216 25480
rect 4580 25440 4586 25452
rect 24210 25440 24216 25452
rect 24268 25440 24274 25492
rect 5258 25372 5264 25424
rect 5316 25412 5322 25424
rect 24762 25412 24768 25424
rect 5316 25384 24768 25412
rect 5316 25372 5322 25384
rect 24762 25372 24768 25384
rect 24820 25372 24826 25424
rect 4798 25304 4804 25356
rect 4856 25344 4862 25356
rect 19518 25344 19524 25356
rect 4856 25316 19524 25344
rect 4856 25304 4862 25316
rect 19518 25304 19524 25316
rect 19576 25304 19582 25356
rect 4154 25236 4160 25288
rect 4212 25276 4218 25288
rect 17954 25276 17960 25288
rect 4212 25248 17960 25276
rect 4212 25236 4218 25248
rect 17954 25236 17960 25248
rect 18012 25236 18018 25288
rect 3234 25168 3240 25220
rect 3292 25208 3298 25220
rect 9490 25208 9496 25220
rect 3292 25180 9496 25208
rect 3292 25168 3298 25180
rect 9490 25168 9496 25180
rect 9548 25168 9554 25220
rect 12618 25168 12624 25220
rect 12676 25208 12682 25220
rect 24026 25208 24032 25220
rect 12676 25180 24032 25208
rect 12676 25168 12682 25180
rect 24026 25168 24032 25180
rect 24084 25168 24090 25220
rect 6730 25100 6736 25152
rect 6788 25140 6794 25152
rect 13906 25140 13912 25152
rect 6788 25112 13912 25140
rect 6788 25100 6794 25112
rect 13906 25100 13912 25112
rect 13964 25100 13970 25152
rect 14274 25072 14280 25084
rect 2746 25044 14280 25072
rect 1118 24964 1124 25016
rect 1176 25004 1182 25016
rect 2746 25004 2774 25044
rect 14274 25032 14280 25044
rect 14332 25032 14338 25084
rect 13078 25004 13084 25016
rect 1176 24976 2774 25004
rect 7576 24976 13084 25004
rect 1176 24964 1182 24976
rect 750 24896 756 24948
rect 808 24936 814 24948
rect 7576 24936 7604 24976
rect 13078 24964 13084 24976
rect 13136 24964 13142 25016
rect 17678 24964 17684 25016
rect 17736 25004 17742 25016
rect 17736 24976 19748 25004
rect 17736 24964 17742 24976
rect 808 24908 7604 24936
rect 808 24896 814 24908
rect 11606 24896 11612 24948
rect 11664 24936 11670 24948
rect 14734 24936 14740 24948
rect 11664 24908 14740 24936
rect 11664 24896 11670 24908
rect 14734 24896 14740 24908
rect 14792 24896 14798 24948
rect 16022 24896 16028 24948
rect 16080 24936 16086 24948
rect 19610 24936 19616 24948
rect 16080 24908 19616 24936
rect 16080 24896 16086 24908
rect 19610 24896 19616 24908
rect 19668 24896 19674 24948
rect 19720 24936 19748 24976
rect 23566 24936 23572 24948
rect 19720 24908 23572 24936
rect 23566 24896 23572 24908
rect 23624 24896 23630 24948
rect 8570 24828 8576 24880
rect 8628 24868 8634 24880
rect 19978 24868 19984 24880
rect 8628 24840 19984 24868
rect 8628 24828 8634 24840
rect 19978 24828 19984 24840
rect 20036 24828 20042 24880
rect 13630 24760 13636 24812
rect 13688 24800 13694 24812
rect 13688 24772 15792 24800
rect 13688 24760 13694 24772
rect 14458 24732 14464 24744
rect 9646 24704 14464 24732
rect 3694 24624 3700 24676
rect 3752 24664 3758 24676
rect 9646 24664 9674 24704
rect 14458 24692 14464 24704
rect 14516 24692 14522 24744
rect 3752 24636 9674 24664
rect 3752 24624 3758 24636
rect 12526 24624 12532 24676
rect 12584 24664 12590 24676
rect 13814 24664 13820 24676
rect 12584 24636 13820 24664
rect 12584 24624 12590 24636
rect 13814 24624 13820 24636
rect 13872 24624 13878 24676
rect 15764 24664 15792 24772
rect 15838 24760 15844 24812
rect 15896 24800 15902 24812
rect 19334 24800 19340 24812
rect 15896 24772 19340 24800
rect 15896 24760 15902 24772
rect 19334 24760 19340 24772
rect 19392 24760 19398 24812
rect 17586 24732 17592 24744
rect 17420 24704 17592 24732
rect 17420 24664 17448 24704
rect 17586 24692 17592 24704
rect 17644 24732 17650 24744
rect 17644 24704 21312 24732
rect 17644 24692 17650 24704
rect 15764 24636 17448 24664
rect 17494 24624 17500 24676
rect 17552 24664 17558 24676
rect 19058 24664 19064 24676
rect 17552 24636 19064 24664
rect 17552 24624 17558 24636
rect 19058 24624 19064 24636
rect 19116 24664 19122 24676
rect 21174 24664 21180 24676
rect 19116 24636 21180 24664
rect 19116 24624 19122 24636
rect 21174 24624 21180 24636
rect 21232 24624 21238 24676
rect 21284 24664 21312 24704
rect 23934 24664 23940 24676
rect 21284 24636 23940 24664
rect 23934 24624 23940 24636
rect 23992 24624 23998 24676
rect 2774 24556 2780 24608
rect 2832 24596 2838 24608
rect 16574 24596 16580 24608
rect 2832 24568 16580 24596
rect 2832 24556 2838 24568
rect 16574 24556 16580 24568
rect 16632 24556 16638 24608
rect 16666 24556 16672 24608
rect 16724 24596 16730 24608
rect 22186 24596 22192 24608
rect 16724 24568 22192 24596
rect 16724 24556 16730 24568
rect 22186 24556 22192 24568
rect 22244 24556 22250 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 1578 24352 1584 24404
rect 1636 24352 1642 24404
rect 6546 24352 6552 24404
rect 6604 24352 6610 24404
rect 8478 24352 8484 24404
rect 8536 24392 8542 24404
rect 15286 24392 15292 24404
rect 8536 24364 15292 24392
rect 8536 24352 8542 24364
rect 15286 24352 15292 24364
rect 15344 24352 15350 24404
rect 15672 24364 18092 24392
rect 3970 24284 3976 24336
rect 4028 24284 4034 24336
rect 6270 24284 6276 24336
rect 6328 24324 6334 24336
rect 6328 24296 6592 24324
rect 6328 24284 6334 24296
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 6454 24256 6460 24268
rect 3283 24228 6460 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 6454 24216 6460 24228
rect 6512 24216 6518 24268
rect 6564 24256 6592 24296
rect 6638 24284 6644 24336
rect 6696 24324 6702 24336
rect 15672 24324 15700 24364
rect 6696 24296 15700 24324
rect 6696 24284 6702 24296
rect 16482 24284 16488 24336
rect 16540 24324 16546 24336
rect 17957 24327 18015 24333
rect 17957 24324 17969 24327
rect 16540 24296 17969 24324
rect 16540 24284 16546 24296
rect 17957 24293 17969 24296
rect 18003 24293 18015 24327
rect 17957 24287 18015 24293
rect 8389 24259 8447 24265
rect 6564 24228 7328 24256
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2314 24188 2320 24200
rect 2271 24160 2320 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2314 24148 2320 24160
rect 2372 24148 2378 24200
rect 4154 24148 4160 24200
rect 4212 24188 4218 24200
rect 4430 24188 4436 24200
rect 4212 24160 4436 24188
rect 4212 24148 4218 24160
rect 4430 24148 4436 24160
rect 4488 24148 4494 24200
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 1762 24012 1768 24064
rect 1820 24012 1826 24064
rect 4816 24052 4844 24151
rect 5902 24148 5908 24200
rect 5960 24188 5966 24200
rect 6733 24191 6791 24197
rect 6733 24188 6745 24191
rect 5960 24160 6745 24188
rect 5960 24148 5966 24160
rect 6733 24157 6745 24160
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 7190 24148 7196 24200
rect 7248 24148 7254 24200
rect 7300 24188 7328 24228
rect 8389 24225 8401 24259
rect 8435 24256 8447 24259
rect 9674 24256 9680 24268
rect 8435 24228 9680 24256
rect 8435 24225 8447 24228
rect 8389 24219 8447 24225
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 11238 24256 11244 24268
rect 11011 24228 11244 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 11238 24216 11244 24228
rect 11296 24216 11302 24268
rect 12434 24216 12440 24268
rect 12492 24256 12498 24268
rect 12805 24259 12863 24265
rect 12805 24256 12817 24259
rect 12492 24228 12817 24256
rect 12492 24216 12498 24228
rect 12805 24225 12817 24228
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 14734 24216 14740 24268
rect 14792 24216 14798 24268
rect 17402 24216 17408 24268
rect 17460 24216 17466 24268
rect 17586 24216 17592 24268
rect 17644 24216 17650 24268
rect 9769 24191 9827 24197
rect 9769 24188 9781 24191
rect 7300 24160 9781 24188
rect 9769 24157 9781 24160
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 5813 24123 5871 24129
rect 5813 24089 5825 24123
rect 5859 24120 5871 24123
rect 8662 24120 8668 24132
rect 5859 24092 8668 24120
rect 5859 24089 5871 24092
rect 5813 24083 5871 24089
rect 8662 24080 8668 24092
rect 8720 24080 8726 24132
rect 11900 24120 11928 24151
rect 12342 24148 12348 24200
rect 12400 24148 12406 24200
rect 13446 24148 13452 24200
rect 13504 24188 13510 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 13504 24160 14289 24188
rect 13504 24148 13510 24160
rect 14277 24157 14289 24160
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24188 16359 24191
rect 16574 24188 16580 24200
rect 16347 24160 16580 24188
rect 16347 24157 16359 24160
rect 16301 24151 16359 24157
rect 16574 24148 16580 24160
rect 16632 24148 16638 24200
rect 16206 24120 16212 24132
rect 8772 24092 11836 24120
rect 11900 24092 16212 24120
rect 7006 24052 7012 24064
rect 4816 24024 7012 24052
rect 7006 24012 7012 24024
rect 7064 24012 7070 24064
rect 7742 24012 7748 24064
rect 7800 24052 7806 24064
rect 8772 24052 8800 24092
rect 7800 24024 8800 24052
rect 9125 24055 9183 24061
rect 7800 24012 7806 24024
rect 9125 24021 9137 24055
rect 9171 24052 9183 24055
rect 11238 24052 11244 24064
rect 9171 24024 11244 24052
rect 9171 24021 9183 24024
rect 9125 24015 9183 24021
rect 11238 24012 11244 24024
rect 11296 24012 11302 24064
rect 11698 24012 11704 24064
rect 11756 24012 11762 24064
rect 11808 24052 11836 24092
rect 16206 24080 16212 24092
rect 16264 24080 16270 24132
rect 16758 24080 16764 24132
rect 16816 24120 16822 24132
rect 17313 24123 17371 24129
rect 17313 24120 17325 24123
rect 16816 24092 17325 24120
rect 16816 24080 16822 24092
rect 17313 24089 17325 24092
rect 17359 24089 17371 24123
rect 17420 24120 17448 24216
rect 17972 24188 18000 24287
rect 18064 24256 18092 24364
rect 18138 24352 18144 24404
rect 18196 24352 18202 24404
rect 18322 24352 18328 24404
rect 18380 24392 18386 24404
rect 19426 24392 19432 24404
rect 18380 24364 19432 24392
rect 18380 24352 18386 24364
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 19610 24352 19616 24404
rect 19668 24352 19674 24404
rect 19978 24352 19984 24404
rect 20036 24352 20042 24404
rect 21726 24352 21732 24404
rect 21784 24392 21790 24404
rect 22005 24395 22063 24401
rect 22005 24392 22017 24395
rect 21784 24364 22017 24392
rect 21784 24352 21790 24364
rect 22005 24361 22017 24364
rect 22051 24392 22063 24395
rect 22446 24395 22504 24401
rect 22446 24392 22458 24395
rect 22051 24364 22458 24392
rect 22051 24361 22063 24364
rect 22005 24355 22063 24361
rect 22446 24361 22458 24364
rect 22492 24361 22504 24395
rect 22446 24355 22504 24361
rect 23934 24352 23940 24404
rect 23992 24392 23998 24404
rect 25498 24392 25504 24404
rect 23992 24364 25504 24392
rect 23992 24352 23998 24364
rect 25498 24352 25504 24364
rect 25556 24352 25562 24404
rect 18966 24284 18972 24336
rect 19024 24324 19030 24336
rect 20165 24327 20223 24333
rect 20165 24324 20177 24327
rect 19024 24296 20177 24324
rect 19024 24284 19030 24296
rect 20165 24293 20177 24296
rect 20211 24293 20223 24327
rect 20165 24287 20223 24293
rect 20254 24284 20260 24336
rect 20312 24324 20318 24336
rect 20312 24296 20852 24324
rect 20312 24284 20318 24296
rect 18693 24259 18751 24265
rect 18693 24256 18705 24259
rect 18064 24228 18705 24256
rect 18693 24225 18705 24228
rect 18739 24256 18751 24259
rect 19702 24256 19708 24268
rect 18739 24228 19708 24256
rect 18739 24225 18751 24228
rect 18693 24219 18751 24225
rect 19702 24216 19708 24228
rect 19760 24216 19766 24268
rect 19794 24216 19800 24268
rect 19852 24256 19858 24268
rect 20717 24259 20775 24265
rect 20717 24256 20729 24259
rect 19852 24228 20729 24256
rect 19852 24216 19858 24228
rect 20717 24225 20729 24228
rect 20763 24225 20775 24259
rect 20824 24256 20852 24296
rect 21174 24284 21180 24336
rect 21232 24284 21238 24336
rect 24581 24327 24639 24333
rect 24581 24293 24593 24327
rect 24627 24324 24639 24327
rect 25038 24324 25044 24336
rect 24627 24296 25044 24324
rect 24627 24293 24639 24296
rect 24581 24287 24639 24293
rect 25038 24284 25044 24296
rect 25096 24284 25102 24336
rect 21821 24259 21879 24265
rect 21821 24256 21833 24259
rect 20824 24228 21833 24256
rect 20717 24219 20775 24225
rect 21821 24225 21833 24228
rect 21867 24225 21879 24259
rect 21821 24219 21879 24225
rect 22189 24259 22247 24265
rect 22189 24225 22201 24259
rect 22235 24256 22247 24259
rect 22554 24256 22560 24268
rect 22235 24228 22560 24256
rect 22235 24225 22247 24228
rect 22189 24219 22247 24225
rect 22554 24216 22560 24228
rect 22612 24216 22618 24268
rect 25225 24259 25283 24265
rect 25225 24225 25237 24259
rect 25271 24256 25283 24259
rect 25314 24256 25320 24268
rect 25271 24228 25320 24256
rect 25271 24225 25283 24228
rect 25225 24219 25283 24225
rect 25314 24216 25320 24228
rect 25372 24216 25378 24268
rect 18509 24191 18567 24197
rect 18509 24188 18521 24191
rect 17972 24160 18521 24188
rect 18509 24157 18521 24160
rect 18555 24157 18567 24191
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 18509 24151 18567 24157
rect 18616 24160 21373 24188
rect 18616 24120 18644 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 23750 24148 23756 24200
rect 23808 24188 23814 24200
rect 24949 24191 25007 24197
rect 24949 24188 24961 24191
rect 23808 24160 24961 24188
rect 23808 24148 23814 24160
rect 24949 24157 24961 24160
rect 24995 24188 25007 24191
rect 25130 24188 25136 24200
rect 24995 24160 25136 24188
rect 24995 24157 25007 24160
rect 24949 24151 25007 24157
rect 25130 24148 25136 24160
rect 25188 24148 25194 24200
rect 17420 24092 18644 24120
rect 19521 24123 19579 24129
rect 17313 24083 17371 24089
rect 19521 24089 19533 24123
rect 19567 24089 19579 24123
rect 19521 24083 19579 24089
rect 15930 24052 15936 24064
rect 11808 24024 15936 24052
rect 15930 24012 15936 24024
rect 15988 24012 15994 24064
rect 16114 24012 16120 24064
rect 16172 24012 16178 24064
rect 16945 24055 17003 24061
rect 16945 24021 16957 24055
rect 16991 24052 17003 24055
rect 17218 24052 17224 24064
rect 16991 24024 17224 24052
rect 16991 24021 17003 24024
rect 16945 24015 17003 24021
rect 17218 24012 17224 24024
rect 17276 24012 17282 24064
rect 18598 24012 18604 24064
rect 18656 24012 18662 24064
rect 19334 24012 19340 24064
rect 19392 24052 19398 24064
rect 19536 24052 19564 24083
rect 19978 24080 19984 24132
rect 20036 24120 20042 24132
rect 20625 24123 20683 24129
rect 20625 24120 20637 24123
rect 20036 24092 20637 24120
rect 20036 24080 20042 24092
rect 20625 24089 20637 24092
rect 20671 24089 20683 24123
rect 20625 24083 20683 24089
rect 21266 24080 21272 24132
rect 21324 24120 21330 24132
rect 21545 24123 21603 24129
rect 21545 24120 21557 24123
rect 21324 24092 21557 24120
rect 21324 24080 21330 24092
rect 21545 24089 21557 24092
rect 21591 24089 21603 24123
rect 21545 24083 21603 24089
rect 22756 24092 22954 24120
rect 19392 24024 19564 24052
rect 19392 24012 19398 24024
rect 20530 24012 20536 24064
rect 20588 24012 20594 24064
rect 22370 24012 22376 24064
rect 22428 24052 22434 24064
rect 22756 24052 22784 24092
rect 23842 24052 23848 24064
rect 22428 24024 23848 24052
rect 22428 24012 22434 24024
rect 23842 24012 23848 24024
rect 23900 24012 23906 24064
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 25590 24052 25596 24064
rect 25087 24024 25596 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 25590 24012 25596 24024
rect 25648 24012 25654 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 2317 23851 2375 23857
rect 2317 23817 2329 23851
rect 2363 23848 2375 23851
rect 2363 23820 6884 23848
rect 2363 23817 2375 23820
rect 2317 23811 2375 23817
rect 6856 23780 6884 23820
rect 7374 23808 7380 23860
rect 7432 23848 7438 23860
rect 7432 23820 12296 23848
rect 7432 23808 7438 23820
rect 12158 23780 12164 23792
rect 6856 23752 12164 23780
rect 12158 23740 12164 23752
rect 12216 23740 12222 23792
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 2590 23712 2596 23724
rect 1719 23684 2596 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 2590 23672 2596 23684
rect 2648 23672 2654 23724
rect 2958 23672 2964 23724
rect 3016 23672 3022 23724
rect 4798 23672 4804 23724
rect 4856 23672 4862 23724
rect 6549 23715 6607 23721
rect 6549 23712 6561 23715
rect 5736 23684 6561 23712
rect 3973 23647 4031 23653
rect 3973 23613 3985 23647
rect 4019 23644 4031 23647
rect 5350 23644 5356 23656
rect 4019 23616 5356 23644
rect 4019 23613 4031 23616
rect 3973 23607 4031 23613
rect 5350 23604 5356 23616
rect 5408 23604 5414 23656
rect 1762 23468 1768 23520
rect 1820 23508 1826 23520
rect 5736 23508 5764 23684
rect 6549 23681 6561 23684
rect 6595 23712 6607 23715
rect 6638 23712 6644 23724
rect 6595 23684 6644 23712
rect 6595 23681 6607 23684
rect 6549 23675 6607 23681
rect 6638 23672 6644 23684
rect 6696 23672 6702 23724
rect 6822 23672 6828 23724
rect 6880 23672 6886 23724
rect 7834 23672 7840 23724
rect 7892 23712 7898 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7892 23684 7941 23712
rect 7892 23672 7898 23684
rect 7929 23681 7941 23684
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 9125 23715 9183 23721
rect 9125 23681 9137 23715
rect 9171 23712 9183 23715
rect 9582 23712 9588 23724
rect 9171 23684 9588 23712
rect 9171 23681 9183 23684
rect 9125 23675 9183 23681
rect 9582 23672 9588 23684
rect 9640 23672 9646 23724
rect 9950 23672 9956 23724
rect 10008 23672 10014 23724
rect 10870 23672 10876 23724
rect 10928 23672 10934 23724
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 10980 23684 12081 23712
rect 5813 23647 5871 23653
rect 5813 23613 5825 23647
rect 5859 23644 5871 23647
rect 7558 23644 7564 23656
rect 5859 23616 7564 23644
rect 5859 23613 5871 23616
rect 5813 23607 5871 23613
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 9214 23604 9220 23656
rect 9272 23644 9278 23656
rect 10980 23644 11008 23684
rect 12069 23681 12081 23684
rect 12115 23681 12127 23715
rect 12268 23712 12296 23820
rect 12434 23808 12440 23860
rect 12492 23848 12498 23860
rect 13630 23848 13636 23860
rect 12492 23820 13636 23848
rect 12492 23808 12498 23820
rect 13630 23808 13636 23820
rect 13688 23808 13694 23860
rect 13817 23851 13875 23857
rect 13817 23817 13829 23851
rect 13863 23848 13875 23851
rect 13906 23848 13912 23860
rect 13863 23820 13912 23848
rect 13863 23817 13875 23820
rect 13817 23811 13875 23817
rect 13906 23808 13912 23820
rect 13964 23848 13970 23860
rect 14461 23851 14519 23857
rect 14461 23848 14473 23851
rect 13964 23820 14473 23848
rect 13964 23808 13970 23820
rect 14461 23817 14473 23820
rect 14507 23817 14519 23851
rect 14461 23811 14519 23817
rect 15562 23808 15568 23860
rect 15620 23848 15626 23860
rect 16853 23851 16911 23857
rect 15620 23820 16620 23848
rect 15620 23808 15626 23820
rect 13354 23740 13360 23792
rect 13412 23780 13418 23792
rect 15933 23783 15991 23789
rect 15933 23780 15945 23783
rect 13412 23752 15945 23780
rect 13412 23740 13418 23752
rect 15933 23749 15945 23752
rect 15979 23749 15991 23783
rect 16592 23780 16620 23820
rect 16853 23817 16865 23851
rect 16899 23848 16911 23851
rect 18506 23848 18512 23860
rect 16899 23820 18512 23848
rect 16899 23817 16911 23820
rect 16853 23811 16911 23817
rect 18506 23808 18512 23820
rect 18564 23808 18570 23860
rect 18598 23808 18604 23860
rect 18656 23848 18662 23860
rect 20349 23851 20407 23857
rect 20349 23848 20361 23851
rect 18656 23820 20361 23848
rect 18656 23808 18662 23820
rect 20349 23817 20361 23820
rect 20395 23817 20407 23851
rect 22370 23848 22376 23860
rect 20349 23811 20407 23817
rect 20456 23820 22376 23848
rect 17221 23783 17279 23789
rect 17221 23780 17233 23783
rect 16592 23752 17233 23780
rect 15933 23743 15991 23749
rect 17221 23749 17233 23752
rect 17267 23780 17279 23783
rect 18322 23780 18328 23792
rect 17267 23752 18328 23780
rect 17267 23749 17279 23752
rect 17221 23743 17279 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 20162 23780 20168 23792
rect 19550 23752 20168 23780
rect 20162 23740 20168 23752
rect 20220 23780 20226 23792
rect 20456 23780 20484 23820
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 20220 23752 20484 23780
rect 20220 23740 20226 23752
rect 20714 23740 20720 23792
rect 20772 23740 20778 23792
rect 22462 23740 22468 23792
rect 22520 23780 22526 23792
rect 22925 23783 22983 23789
rect 22925 23780 22937 23783
rect 22520 23752 22937 23780
rect 22520 23740 22526 23752
rect 22925 23749 22937 23752
rect 22971 23749 22983 23783
rect 22925 23743 22983 23749
rect 23382 23740 23388 23792
rect 23440 23740 23446 23792
rect 12268 23684 12664 23712
rect 12069 23675 12127 23681
rect 9272 23616 11008 23644
rect 9272 23604 9278 23616
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12032 23616 12541 23644
rect 12032 23604 12038 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12636 23644 12664 23684
rect 15286 23672 15292 23724
rect 15344 23672 15350 23724
rect 17310 23672 17316 23724
rect 17368 23672 17374 23724
rect 20809 23715 20867 23721
rect 20809 23681 20821 23715
rect 20855 23712 20867 23715
rect 21358 23712 21364 23724
rect 20855 23684 21364 23712
rect 20855 23681 20867 23684
rect 20809 23675 20867 23681
rect 21358 23672 21364 23684
rect 21416 23672 21422 23724
rect 22186 23672 22192 23724
rect 22244 23672 22250 23724
rect 25041 23715 25099 23721
rect 25041 23681 25053 23715
rect 25087 23712 25099 23715
rect 25406 23712 25412 23724
rect 25087 23684 25412 23712
rect 25087 23681 25099 23684
rect 25041 23675 25099 23681
rect 25406 23672 25412 23684
rect 25464 23672 25470 23724
rect 14553 23647 14611 23653
rect 12636 23616 13860 23644
rect 12529 23607 12587 23613
rect 7190 23576 7196 23588
rect 5828 23548 7196 23576
rect 5828 23520 5856 23548
rect 7190 23536 7196 23548
rect 7248 23536 7254 23588
rect 9674 23536 9680 23588
rect 9732 23576 9738 23588
rect 9732 23548 12434 23576
rect 9732 23536 9738 23548
rect 1820 23480 5764 23508
rect 1820 23468 1826 23480
rect 5810 23468 5816 23520
rect 5868 23468 5874 23520
rect 6638 23468 6644 23520
rect 6696 23508 6702 23520
rect 7469 23511 7527 23517
rect 7469 23508 7481 23511
rect 6696 23480 7481 23508
rect 6696 23468 6702 23480
rect 7469 23477 7481 23480
rect 7515 23477 7527 23511
rect 7469 23471 7527 23477
rect 11606 23468 11612 23520
rect 11664 23468 11670 23520
rect 11698 23468 11704 23520
rect 11756 23468 11762 23520
rect 12406 23508 12434 23548
rect 13722 23508 13728 23520
rect 12406 23480 13728 23508
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 13832 23508 13860 23616
rect 14553 23613 14565 23647
rect 14599 23613 14611 23647
rect 14553 23607 14611 23613
rect 14090 23536 14096 23588
rect 14148 23536 14154 23588
rect 14568 23576 14596 23607
rect 14642 23604 14648 23656
rect 14700 23604 14706 23656
rect 16301 23647 16359 23653
rect 16301 23613 16313 23647
rect 16347 23644 16359 23647
rect 16942 23644 16948 23656
rect 16347 23616 16948 23644
rect 16347 23613 16359 23616
rect 16301 23607 16359 23613
rect 16942 23604 16948 23616
rect 17000 23604 17006 23656
rect 17497 23647 17555 23653
rect 17497 23613 17509 23647
rect 17543 23613 17555 23647
rect 17497 23607 17555 23613
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23613 18107 23647
rect 18049 23607 18107 23613
rect 18325 23647 18383 23653
rect 18325 23613 18337 23647
rect 18371 23644 18383 23647
rect 18782 23644 18788 23656
rect 18371 23616 18788 23644
rect 18371 23613 18383 23616
rect 18325 23607 18383 23613
rect 14568 23548 16896 23576
rect 14826 23508 14832 23520
rect 13832 23480 14832 23508
rect 14826 23468 14832 23480
rect 14884 23468 14890 23520
rect 16482 23468 16488 23520
rect 16540 23468 16546 23520
rect 16868 23508 16896 23548
rect 17034 23536 17040 23588
rect 17092 23576 17098 23588
rect 17512 23576 17540 23607
rect 17092 23548 17540 23576
rect 17092 23536 17098 23548
rect 17770 23508 17776 23520
rect 16868 23480 17776 23508
rect 17770 23468 17776 23480
rect 17828 23468 17834 23520
rect 18064 23508 18092 23607
rect 18782 23604 18788 23616
rect 18840 23604 18846 23656
rect 19702 23604 19708 23656
rect 19760 23644 19766 23656
rect 20714 23644 20720 23656
rect 19760 23616 20720 23644
rect 19760 23604 19766 23616
rect 20714 23604 20720 23616
rect 20772 23604 20778 23656
rect 20898 23604 20904 23656
rect 20956 23604 20962 23656
rect 20990 23604 20996 23656
rect 21048 23644 21054 23656
rect 22462 23644 22468 23656
rect 21048 23616 22468 23644
rect 21048 23604 21054 23616
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 22646 23604 22652 23656
rect 22704 23604 22710 23656
rect 21082 23536 21088 23588
rect 21140 23576 21146 23588
rect 22005 23579 22063 23585
rect 22005 23576 22017 23579
rect 21140 23548 22017 23576
rect 21140 23536 21146 23548
rect 22005 23545 22017 23548
rect 22051 23545 22063 23579
rect 22005 23539 22063 23545
rect 25222 23536 25228 23588
rect 25280 23536 25286 23588
rect 18322 23508 18328 23520
rect 18064 23480 18328 23508
rect 18322 23468 18328 23480
rect 18380 23468 18386 23520
rect 19794 23468 19800 23520
rect 19852 23468 19858 23520
rect 20070 23468 20076 23520
rect 20128 23508 20134 23520
rect 21361 23511 21419 23517
rect 21361 23508 21373 23511
rect 20128 23480 21373 23508
rect 20128 23468 20134 23480
rect 21361 23477 21373 23480
rect 21407 23477 21419 23511
rect 21361 23471 21419 23477
rect 21542 23468 21548 23520
rect 21600 23468 21606 23520
rect 24394 23468 24400 23520
rect 24452 23468 24458 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 1581 23307 1639 23313
rect 1581 23273 1593 23307
rect 1627 23304 1639 23307
rect 3694 23304 3700 23316
rect 1627 23276 3700 23304
rect 1627 23273 1639 23276
rect 1581 23267 1639 23273
rect 3694 23264 3700 23276
rect 3752 23264 3758 23316
rect 4893 23307 4951 23313
rect 4893 23273 4905 23307
rect 4939 23304 4951 23307
rect 9674 23304 9680 23316
rect 4939 23276 9680 23304
rect 4939 23273 4951 23276
rect 4893 23267 4951 23273
rect 9674 23264 9680 23276
rect 9732 23264 9738 23316
rect 11882 23264 11888 23316
rect 11940 23304 11946 23316
rect 12526 23304 12532 23316
rect 11940 23276 12532 23304
rect 11940 23264 11946 23276
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 12618 23264 12624 23316
rect 12676 23304 12682 23316
rect 13446 23304 13452 23316
rect 12676 23276 13452 23304
rect 12676 23264 12682 23276
rect 13446 23264 13452 23276
rect 13504 23264 13510 23316
rect 13538 23264 13544 23316
rect 13596 23304 13602 23316
rect 15838 23304 15844 23316
rect 13596 23276 15844 23304
rect 13596 23264 13602 23276
rect 15838 23264 15844 23276
rect 15896 23264 15902 23316
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 17862 23304 17868 23316
rect 16632 23276 17868 23304
rect 16632 23264 16638 23276
rect 17862 23264 17868 23276
rect 17920 23304 17926 23316
rect 18969 23307 19027 23313
rect 18969 23304 18981 23307
rect 17920 23276 18981 23304
rect 17920 23264 17926 23276
rect 18969 23273 18981 23276
rect 19015 23273 19027 23307
rect 20254 23304 20260 23316
rect 18969 23267 19027 23273
rect 19076 23276 20260 23304
rect 3142 23196 3148 23248
rect 3200 23236 3206 23248
rect 3200 23208 10732 23236
rect 3200 23196 3206 23208
rect 3237 23171 3295 23177
rect 3237 23137 3249 23171
rect 3283 23168 3295 23171
rect 4614 23168 4620 23180
rect 3283 23140 4620 23168
rect 3283 23137 3295 23140
rect 3237 23131 3295 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 6457 23171 6515 23177
rect 6457 23137 6469 23171
rect 6503 23168 6515 23171
rect 7650 23168 7656 23180
rect 6503 23140 7656 23168
rect 6503 23137 6515 23140
rect 6457 23131 6515 23137
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23168 8263 23171
rect 9306 23168 9312 23180
rect 8251 23140 9312 23168
rect 8251 23137 8263 23140
rect 8205 23131 8263 23137
rect 9306 23128 9312 23140
rect 9364 23128 9370 23180
rect 9398 23128 9404 23180
rect 9456 23168 9462 23180
rect 10597 23171 10655 23177
rect 10597 23168 10609 23171
rect 9456 23140 10609 23168
rect 9456 23128 9462 23140
rect 10597 23137 10609 23140
rect 10643 23137 10655 23171
rect 10704 23168 10732 23208
rect 12986 23196 12992 23248
rect 13044 23236 13050 23248
rect 13044 23208 15148 23236
rect 13044 23196 13050 23208
rect 14642 23168 14648 23180
rect 10704 23140 14648 23168
rect 10597 23131 10655 23137
rect 14642 23128 14648 23140
rect 14700 23128 14706 23180
rect 15120 23168 15148 23208
rect 16298 23196 16304 23248
rect 16356 23236 16362 23248
rect 16356 23208 17908 23236
rect 16356 23196 16362 23208
rect 17402 23168 17408 23180
rect 15120 23140 17408 23168
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 17494 23128 17500 23180
rect 17552 23168 17558 23180
rect 17773 23171 17831 23177
rect 17773 23168 17785 23171
rect 17552 23140 17785 23168
rect 17552 23128 17558 23140
rect 17773 23137 17785 23140
rect 17819 23137 17831 23171
rect 17880 23168 17908 23208
rect 18690 23196 18696 23248
rect 18748 23196 18754 23248
rect 18874 23196 18880 23248
rect 18932 23236 18938 23248
rect 19076 23236 19104 23276
rect 20254 23264 20260 23276
rect 20312 23264 20318 23316
rect 20714 23264 20720 23316
rect 20772 23304 20778 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 20772 23276 21189 23304
rect 20772 23264 20778 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 24302 23264 24308 23316
rect 24360 23304 24366 23316
rect 24397 23307 24455 23313
rect 24397 23304 24409 23307
rect 24360 23276 24409 23304
rect 24360 23264 24366 23276
rect 24397 23273 24409 23276
rect 24443 23273 24455 23307
rect 24397 23267 24455 23273
rect 18932 23208 19104 23236
rect 18932 23196 18938 23208
rect 19429 23171 19487 23177
rect 17880 23140 19104 23168
rect 17773 23131 17831 23137
rect 2222 23060 2228 23112
rect 2280 23060 2286 23112
rect 4246 23060 4252 23112
rect 4304 23060 4310 23112
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23100 5503 23103
rect 6546 23100 6552 23112
rect 5491 23072 6552 23100
rect 5491 23069 5503 23072
rect 5445 23063 5503 23069
rect 6546 23060 6552 23072
rect 6604 23060 6610 23112
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 1765 22967 1823 22973
rect 1765 22933 1777 22967
rect 1811 22964 1823 22967
rect 3694 22964 3700 22976
rect 1811 22936 3700 22964
rect 1811 22933 1823 22936
rect 1765 22927 1823 22933
rect 3694 22924 3700 22936
rect 3752 22924 3758 22976
rect 3973 22967 4031 22973
rect 3973 22933 3985 22967
rect 4019 22964 4031 22967
rect 4614 22964 4620 22976
rect 4019 22936 4620 22964
rect 4019 22933 4031 22936
rect 3973 22927 4031 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 6178 22924 6184 22976
rect 6236 22964 6242 22976
rect 7208 22964 7236 23063
rect 7282 23060 7288 23112
rect 7340 23100 7346 23112
rect 9214 23100 9220 23112
rect 7340 23072 9220 23100
rect 7340 23060 7346 23072
rect 9214 23060 9220 23072
rect 9272 23060 9278 23112
rect 9490 23060 9496 23112
rect 9548 23060 9554 23112
rect 13081 23103 13139 23109
rect 13081 23069 13093 23103
rect 13127 23100 13139 23103
rect 13354 23100 13360 23112
rect 13127 23072 13360 23100
rect 13127 23069 13139 23072
rect 13081 23063 13139 23069
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 13630 23060 13636 23112
rect 13688 23100 13694 23112
rect 15013 23103 15071 23109
rect 15013 23100 15025 23103
rect 13688 23072 15025 23100
rect 13688 23060 13694 23072
rect 15013 23069 15025 23072
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 16666 23060 16672 23112
rect 16724 23100 16730 23112
rect 17034 23100 17040 23112
rect 16724 23072 17040 23100
rect 16724 23060 16730 23072
rect 17034 23060 17040 23072
rect 17092 23060 17098 23112
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23100 17647 23103
rect 18966 23100 18972 23112
rect 17635 23072 18972 23100
rect 17635 23069 17647 23072
rect 17589 23063 17647 23069
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 9033 23035 9091 23041
rect 9033 23001 9045 23035
rect 9079 23032 9091 23035
rect 9508 23032 9536 23060
rect 9079 23004 9536 23032
rect 9079 23001 9091 23004
rect 9033 22995 9091 23001
rect 10594 22992 10600 23044
rect 10652 23032 10658 23044
rect 10873 23035 10931 23041
rect 10873 23032 10885 23035
rect 10652 23004 10885 23032
rect 10652 22992 10658 23004
rect 10873 23001 10885 23004
rect 10919 23001 10931 23035
rect 12250 23032 12256 23044
rect 12098 23004 12256 23032
rect 10873 22995 10931 23001
rect 6236 22936 7236 22964
rect 10137 22967 10195 22973
rect 6236 22924 6242 22936
rect 10137 22933 10149 22967
rect 10183 22964 10195 22967
rect 10778 22964 10784 22976
rect 10183 22936 10784 22964
rect 10183 22933 10195 22936
rect 10137 22927 10195 22933
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 11606 22924 11612 22976
rect 11664 22964 11670 22976
rect 12176 22964 12204 23004
rect 12250 22992 12256 23004
rect 12308 22992 12314 23044
rect 13170 22992 13176 23044
rect 13228 23032 13234 23044
rect 13228 23004 14320 23032
rect 13228 22992 13234 23004
rect 11664 22936 12204 22964
rect 11664 22924 11670 22936
rect 12342 22924 12348 22976
rect 12400 22924 12406 22976
rect 12618 22924 12624 22976
rect 12676 22964 12682 22976
rect 12713 22967 12771 22973
rect 12713 22964 12725 22967
rect 12676 22936 12725 22964
rect 12676 22924 12682 22936
rect 12713 22933 12725 22936
rect 12759 22933 12771 22967
rect 12713 22927 12771 22933
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 13725 22967 13783 22973
rect 13725 22964 13737 22967
rect 12860 22936 13737 22964
rect 12860 22924 12866 22936
rect 13725 22933 13737 22936
rect 13771 22933 13783 22967
rect 14292 22964 14320 23004
rect 14366 22992 14372 23044
rect 14424 22992 14430 23044
rect 14550 22992 14556 23044
rect 14608 22992 14614 23044
rect 14734 22992 14740 23044
rect 14792 23032 14798 23044
rect 15289 23035 15347 23041
rect 15289 23032 15301 23035
rect 14792 23004 15301 23032
rect 14792 22992 14798 23004
rect 15289 23001 15301 23004
rect 15335 23001 15347 23035
rect 16942 23032 16948 23044
rect 16514 23004 16948 23032
rect 15289 22995 15347 23001
rect 16942 22992 16948 23004
rect 17000 22992 17006 23044
rect 18509 23035 18567 23041
rect 18509 23001 18521 23035
rect 18555 23032 18567 23035
rect 18874 23032 18880 23044
rect 18555 23004 18880 23032
rect 18555 23001 18567 23004
rect 18509 22995 18567 23001
rect 18874 22992 18880 23004
rect 18932 22992 18938 23044
rect 16761 22967 16819 22973
rect 16761 22964 16773 22967
rect 14292 22936 16773 22964
rect 13725 22927 13783 22933
rect 16761 22933 16773 22936
rect 16807 22964 16819 22967
rect 17126 22964 17132 22976
rect 16807 22936 17132 22964
rect 16807 22933 16819 22936
rect 16761 22927 16819 22933
rect 17126 22924 17132 22936
rect 17184 22924 17190 22976
rect 17218 22924 17224 22976
rect 17276 22924 17282 22976
rect 17678 22924 17684 22976
rect 17736 22924 17742 22976
rect 19076 22964 19104 23140
rect 19429 23137 19441 23171
rect 19475 23168 19487 23171
rect 21637 23171 21695 23177
rect 21637 23168 21649 23171
rect 19475 23140 21649 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 21637 23137 21649 23140
rect 21683 23168 21695 23171
rect 22646 23168 22652 23180
rect 21683 23140 22652 23168
rect 21683 23137 21695 23140
rect 21637 23131 21695 23137
rect 22646 23128 22652 23140
rect 22704 23128 22710 23180
rect 24412 23168 24440 23267
rect 25041 23171 25099 23177
rect 25041 23168 25053 23171
rect 24412 23140 25053 23168
rect 25041 23137 25053 23140
rect 25087 23137 25099 23171
rect 25041 23131 25099 23137
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 23382 23100 23388 23112
rect 23046 23072 23388 23100
rect 23382 23060 23388 23072
rect 23440 23060 23446 23112
rect 24946 23060 24952 23112
rect 25004 23100 25010 23112
rect 25222 23100 25228 23112
rect 25004 23072 25228 23100
rect 25004 23060 25010 23072
rect 25222 23060 25228 23072
rect 25280 23060 25286 23112
rect 19702 22992 19708 23044
rect 19760 22992 19766 23044
rect 20162 22992 20168 23044
rect 20220 22992 20226 23044
rect 21910 22992 21916 23044
rect 21968 22992 21974 23044
rect 26878 23032 26884 23044
rect 23216 23004 26884 23032
rect 20530 22964 20536 22976
rect 19076 22936 20536 22964
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 22278 22924 22284 22976
rect 22336 22964 22342 22976
rect 23216 22964 23244 23004
rect 26878 22992 26884 23004
rect 26936 22992 26942 23044
rect 22336 22936 23244 22964
rect 22336 22924 22342 22936
rect 23382 22924 23388 22976
rect 23440 22924 23446 22976
rect 23842 22924 23848 22976
rect 23900 22924 23906 22976
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 2498 22720 2504 22772
rect 2556 22760 2562 22772
rect 3418 22760 3424 22772
rect 2556 22732 3424 22760
rect 2556 22720 2562 22732
rect 3418 22720 3424 22732
rect 3476 22720 3482 22772
rect 5994 22720 6000 22772
rect 6052 22760 6058 22772
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 6052 22732 6561 22760
rect 6052 22720 6058 22732
rect 6549 22729 6561 22732
rect 6595 22760 6607 22763
rect 6730 22760 6736 22772
rect 6595 22732 6736 22760
rect 6595 22729 6607 22732
rect 6549 22723 6607 22729
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 7006 22720 7012 22772
rect 7064 22720 7070 22772
rect 11790 22720 11796 22772
rect 11848 22760 11854 22772
rect 14734 22760 14740 22772
rect 11848 22732 14740 22760
rect 11848 22720 11854 22732
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 15286 22760 15292 22772
rect 15212 22732 15292 22760
rect 3142 22692 3148 22704
rect 1688 22664 3148 22692
rect 1688 22633 1716 22664
rect 3142 22652 3148 22664
rect 3200 22652 3206 22704
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 4154 22692 4160 22704
rect 4019 22664 4160 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 4154 22652 4160 22664
rect 4212 22652 4218 22704
rect 5718 22652 5724 22704
rect 5776 22652 5782 22704
rect 8754 22652 8760 22704
rect 8812 22652 8818 22704
rect 11606 22692 11612 22704
rect 10902 22664 11612 22692
rect 11606 22652 11612 22664
rect 11664 22652 11670 22704
rect 12526 22652 12532 22704
rect 12584 22692 12590 22704
rect 13538 22692 13544 22704
rect 12584 22664 13544 22692
rect 12584 22652 12590 22664
rect 13538 22652 13544 22664
rect 13596 22652 13602 22704
rect 15212 22692 15240 22732
rect 15286 22720 15292 22732
rect 15344 22760 15350 22772
rect 16942 22760 16948 22772
rect 15344 22732 16948 22760
rect 15344 22720 15350 22732
rect 16942 22720 16948 22732
rect 17000 22720 17006 22772
rect 17126 22720 17132 22772
rect 17184 22760 17190 22772
rect 18049 22763 18107 22769
rect 17184 22732 18000 22760
rect 17184 22720 17190 22732
rect 15134 22664 15240 22692
rect 15470 22652 15476 22704
rect 15528 22692 15534 22704
rect 17221 22695 17279 22701
rect 17221 22692 17233 22695
rect 15528 22664 17233 22692
rect 15528 22652 15534 22664
rect 17221 22661 17233 22664
rect 17267 22692 17279 22695
rect 17862 22692 17868 22704
rect 17267 22664 17868 22692
rect 17267 22661 17279 22664
rect 17221 22655 17279 22661
rect 17862 22652 17868 22664
rect 17920 22652 17926 22704
rect 17972 22692 18000 22732
rect 18049 22729 18061 22763
rect 18095 22760 18107 22763
rect 18414 22760 18420 22772
rect 18095 22732 18420 22760
rect 18095 22729 18107 22732
rect 18049 22723 18107 22729
rect 18414 22720 18420 22732
rect 18472 22720 18478 22772
rect 18509 22763 18567 22769
rect 18509 22729 18521 22763
rect 18555 22760 18567 22763
rect 20441 22763 20499 22769
rect 20441 22760 20453 22763
rect 18555 22732 20453 22760
rect 18555 22729 18567 22732
rect 18509 22723 18567 22729
rect 20441 22729 20453 22732
rect 20487 22729 20499 22763
rect 20441 22723 20499 22729
rect 20530 22720 20536 22772
rect 20588 22760 20594 22772
rect 22554 22760 22560 22772
rect 20588 22732 22560 22760
rect 20588 22720 20594 22732
rect 22554 22720 22560 22732
rect 22612 22720 22618 22772
rect 23106 22720 23112 22772
rect 23164 22760 23170 22772
rect 24857 22763 24915 22769
rect 24857 22760 24869 22763
rect 23164 22732 24869 22760
rect 23164 22720 23170 22732
rect 24857 22729 24869 22732
rect 24903 22760 24915 22763
rect 24946 22760 24952 22772
rect 24903 22732 24952 22760
rect 24903 22729 24915 22732
rect 24857 22723 24915 22729
rect 24946 22720 24952 22732
rect 25004 22720 25010 22772
rect 17972 22664 21680 22692
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22593 1731 22627
rect 1673 22587 1731 22593
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 3602 22624 3608 22636
rect 3007 22596 3608 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 3602 22584 3608 22596
rect 3660 22584 3666 22636
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7098 22624 7104 22636
rect 6963 22596 7104 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7098 22584 7104 22596
rect 7156 22584 7162 22636
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 6362 22516 6368 22568
rect 6420 22556 6426 22568
rect 7576 22556 7604 22587
rect 8938 22584 8944 22636
rect 8996 22624 9002 22636
rect 9398 22624 9404 22636
rect 8996 22596 9404 22624
rect 8996 22584 9002 22596
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 11146 22584 11152 22636
rect 11204 22624 11210 22636
rect 11977 22627 12035 22633
rect 11977 22624 11989 22627
rect 11204 22596 11989 22624
rect 11204 22584 11210 22596
rect 11977 22593 11989 22596
rect 12023 22593 12035 22627
rect 11977 22587 12035 22593
rect 12158 22584 12164 22636
rect 12216 22624 12222 22636
rect 12216 22596 12572 22624
rect 12216 22584 12222 22596
rect 6420 22528 7604 22556
rect 9677 22559 9735 22565
rect 6420 22516 6426 22528
rect 9677 22525 9689 22559
rect 9723 22556 9735 22559
rect 9766 22556 9772 22568
rect 9723 22528 9772 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 9766 22516 9772 22528
rect 9824 22516 9830 22568
rect 11698 22516 11704 22568
rect 11756 22516 11762 22568
rect 12066 22516 12072 22568
rect 12124 22556 12130 22568
rect 12434 22556 12440 22568
rect 12124 22528 12440 22556
rect 12124 22516 12130 22528
rect 12434 22516 12440 22528
rect 12492 22516 12498 22568
rect 12544 22556 12572 22596
rect 12710 22584 12716 22636
rect 12768 22624 12774 22636
rect 13173 22627 13231 22633
rect 13173 22624 13185 22627
rect 12768 22596 13185 22624
rect 12768 22584 12774 22596
rect 13173 22593 13185 22596
rect 13219 22624 13231 22627
rect 13446 22624 13452 22636
rect 13219 22596 13452 22624
rect 13219 22593 13231 22596
rect 13173 22587 13231 22593
rect 13446 22584 13452 22596
rect 13504 22584 13510 22636
rect 13630 22584 13636 22636
rect 13688 22584 13694 22636
rect 15930 22584 15936 22636
rect 15988 22584 15994 22636
rect 16022 22584 16028 22636
rect 16080 22624 16086 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 16080 22596 16129 22624
rect 16080 22584 16086 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 17313 22627 17371 22633
rect 17313 22624 17325 22627
rect 16117 22587 16175 22593
rect 17144 22596 17325 22624
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 12544 22528 13921 22556
rect 13909 22525 13921 22528
rect 13955 22525 13967 22559
rect 13909 22519 13967 22525
rect 13998 22516 14004 22568
rect 14056 22556 14062 22568
rect 14056 22528 16896 22556
rect 14056 22516 14062 22528
rect 5534 22448 5540 22500
rect 5592 22488 5598 22500
rect 9398 22488 9404 22500
rect 5592 22460 9404 22488
rect 5592 22448 5598 22460
rect 9398 22448 9404 22460
rect 9456 22448 9462 22500
rect 10704 22460 12434 22488
rect 1670 22380 1676 22432
rect 1728 22420 1734 22432
rect 2317 22423 2375 22429
rect 2317 22420 2329 22423
rect 1728 22392 2329 22420
rect 1728 22380 1734 22392
rect 2317 22389 2329 22392
rect 2363 22389 2375 22423
rect 2317 22383 2375 22389
rect 3418 22380 3424 22432
rect 3476 22420 3482 22432
rect 10704 22420 10732 22460
rect 3476 22392 10732 22420
rect 11149 22423 11207 22429
rect 3476 22380 3482 22392
rect 11149 22389 11161 22423
rect 11195 22420 11207 22423
rect 11330 22420 11336 22432
rect 11195 22392 11336 22420
rect 11195 22389 11207 22392
rect 11149 22383 11207 22389
rect 11330 22380 11336 22392
rect 11388 22380 11394 22432
rect 12406 22420 12434 22460
rect 12912 22460 13124 22488
rect 12912 22420 12940 22460
rect 12406 22392 12940 22420
rect 12986 22380 12992 22432
rect 13044 22380 13050 22432
rect 13096 22420 13124 22460
rect 15746 22448 15752 22500
rect 15804 22488 15810 22500
rect 16868 22497 16896 22528
rect 16942 22516 16948 22568
rect 17000 22556 17006 22568
rect 17144 22556 17172 22596
rect 17313 22593 17325 22596
rect 17359 22593 17371 22627
rect 17313 22587 17371 22593
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22624 18475 22627
rect 18598 22624 18604 22636
rect 18463 22596 18604 22624
rect 18463 22593 18475 22596
rect 18417 22587 18475 22593
rect 18598 22584 18604 22596
rect 18656 22584 18662 22636
rect 19610 22584 19616 22636
rect 19668 22584 19674 22636
rect 17000 22528 17172 22556
rect 17405 22559 17463 22565
rect 17000 22516 17006 22528
rect 17405 22525 17417 22559
rect 17451 22525 17463 22559
rect 17405 22519 17463 22525
rect 16393 22491 16451 22497
rect 16393 22488 16405 22491
rect 15804 22460 16405 22488
rect 15804 22448 15810 22460
rect 16393 22457 16405 22460
rect 16439 22457 16451 22491
rect 16393 22451 16451 22457
rect 16853 22491 16911 22497
rect 16853 22457 16865 22491
rect 16899 22457 16911 22491
rect 17420 22488 17448 22519
rect 17586 22516 17592 22568
rect 17644 22556 17650 22568
rect 18693 22559 18751 22565
rect 17644 22528 18644 22556
rect 17644 22516 17650 22528
rect 16853 22451 16911 22457
rect 16960 22460 17448 22488
rect 13906 22420 13912 22432
rect 13096 22392 13912 22420
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 14642 22380 14648 22432
rect 14700 22420 14706 22432
rect 15381 22423 15439 22429
rect 15381 22420 15393 22423
rect 14700 22392 15393 22420
rect 14700 22380 14706 22392
rect 15381 22389 15393 22392
rect 15427 22389 15439 22423
rect 15381 22383 15439 22389
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 16960 22420 16988 22460
rect 17770 22448 17776 22500
rect 17828 22488 17834 22500
rect 17828 22460 18184 22488
rect 17828 22448 17834 22460
rect 15896 22392 16988 22420
rect 18156 22420 18184 22460
rect 18230 22448 18236 22500
rect 18288 22488 18294 22500
rect 18414 22488 18420 22500
rect 18288 22460 18420 22488
rect 18288 22448 18294 22460
rect 18414 22448 18420 22460
rect 18472 22448 18478 22500
rect 18616 22488 18644 22528
rect 18693 22525 18705 22559
rect 18739 22556 18751 22559
rect 18966 22556 18972 22568
rect 18739 22528 18972 22556
rect 18739 22525 18751 22528
rect 18693 22519 18751 22525
rect 18966 22516 18972 22528
rect 19024 22516 19030 22568
rect 19812 22565 19840 22664
rect 20806 22584 20812 22636
rect 20864 22584 20870 22636
rect 20916 22596 21312 22624
rect 20916 22565 20944 22596
rect 19705 22559 19763 22565
rect 19705 22556 19717 22559
rect 19076 22528 19717 22556
rect 19076 22488 19104 22528
rect 19705 22525 19717 22528
rect 19751 22525 19763 22559
rect 19705 22519 19763 22525
rect 19797 22559 19855 22565
rect 19797 22525 19809 22559
rect 19843 22525 19855 22559
rect 20901 22559 20959 22565
rect 20901 22556 20913 22559
rect 19797 22519 19855 22525
rect 19904 22528 20913 22556
rect 18616 22460 19104 22488
rect 19150 22448 19156 22500
rect 19208 22488 19214 22500
rect 19720 22488 19748 22519
rect 19904 22488 19932 22528
rect 20901 22525 20913 22528
rect 20947 22525 20959 22559
rect 20901 22519 20959 22525
rect 20993 22559 21051 22565
rect 20993 22525 21005 22559
rect 21039 22525 21051 22559
rect 21284 22556 21312 22596
rect 21450 22584 21456 22636
rect 21508 22584 21514 22636
rect 21542 22556 21548 22568
rect 21284 22528 21548 22556
rect 20993 22519 21051 22525
rect 19208 22460 19380 22488
rect 19720 22460 19932 22488
rect 19208 22448 19214 22460
rect 19245 22423 19303 22429
rect 19245 22420 19257 22423
rect 18156 22392 19257 22420
rect 15896 22380 15902 22392
rect 19245 22389 19257 22392
rect 19291 22389 19303 22423
rect 19352 22420 19380 22460
rect 20714 22448 20720 22500
rect 20772 22488 20778 22500
rect 21008 22488 21036 22519
rect 21542 22516 21548 22528
rect 21600 22516 21606 22568
rect 21652 22488 21680 22664
rect 22646 22652 22652 22704
rect 22704 22692 22710 22704
rect 23290 22692 23296 22704
rect 22704 22664 23296 22692
rect 22704 22652 22710 22664
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22624 22063 22627
rect 22278 22624 22284 22636
rect 22051 22596 22284 22624
rect 22051 22593 22063 22596
rect 22005 22587 22063 22593
rect 22278 22584 22284 22596
rect 22336 22584 22342 22636
rect 23124 22633 23152 22664
rect 23290 22652 23296 22664
rect 23348 22652 23354 22704
rect 23934 22652 23940 22704
rect 23992 22652 23998 22704
rect 22925 22627 22983 22633
rect 22925 22624 22937 22627
rect 22480 22596 22937 22624
rect 21726 22516 21732 22568
rect 21784 22556 21790 22568
rect 22480 22556 22508 22596
rect 22925 22593 22937 22596
rect 22971 22593 22983 22627
rect 22925 22587 22983 22593
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 21784 22528 22508 22556
rect 21784 22516 21790 22528
rect 22554 22516 22560 22568
rect 22612 22556 22618 22568
rect 22649 22559 22707 22565
rect 22649 22556 22661 22559
rect 22612 22528 22661 22556
rect 22612 22516 22618 22528
rect 22649 22525 22661 22528
rect 22695 22525 22707 22559
rect 22940 22556 22968 22587
rect 23385 22559 23443 22565
rect 23385 22556 23397 22559
rect 22940 22528 23397 22556
rect 22649 22519 22707 22525
rect 23385 22525 23397 22528
rect 23431 22525 23443 22559
rect 23385 22519 23443 22525
rect 24854 22516 24860 22568
rect 24912 22556 24918 22568
rect 25133 22559 25191 22565
rect 25133 22556 25145 22559
rect 24912 22528 25145 22556
rect 24912 22516 24918 22528
rect 25133 22525 25145 22528
rect 25179 22525 25191 22559
rect 25133 22519 25191 22525
rect 25317 22491 25375 22497
rect 25317 22488 25329 22491
rect 20772 22460 21036 22488
rect 21100 22460 21588 22488
rect 21652 22460 23244 22488
rect 20772 22448 20778 22460
rect 21100 22420 21128 22460
rect 19352 22392 21128 22420
rect 21560 22420 21588 22460
rect 23106 22420 23112 22432
rect 21560 22392 23112 22420
rect 19245 22383 19303 22389
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 23216 22420 23244 22460
rect 24412 22460 25329 22488
rect 24412 22420 24440 22460
rect 25317 22457 25329 22460
rect 25363 22457 25375 22491
rect 25317 22451 25375 22457
rect 23216 22392 24440 22420
rect 26050 22380 26056 22432
rect 26108 22420 26114 22432
rect 26694 22420 26700 22432
rect 26108 22392 26700 22420
rect 26108 22380 26114 22392
rect 26694 22380 26700 22392
rect 26752 22380 26758 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 1581 22219 1639 22225
rect 1581 22185 1593 22219
rect 1627 22216 1639 22219
rect 1854 22216 1860 22228
rect 1627 22188 1860 22216
rect 1627 22185 1639 22188
rect 1581 22179 1639 22185
rect 1854 22176 1860 22188
rect 1912 22176 1918 22228
rect 5626 22176 5632 22228
rect 5684 22216 5690 22228
rect 13354 22216 13360 22228
rect 5684 22188 13360 22216
rect 5684 22176 5690 22188
rect 13354 22176 13360 22188
rect 13412 22176 13418 22228
rect 13446 22176 13452 22228
rect 13504 22176 13510 22228
rect 14182 22176 14188 22228
rect 14240 22216 14246 22228
rect 15194 22216 15200 22228
rect 14240 22188 15200 22216
rect 14240 22176 14246 22188
rect 15194 22176 15200 22188
rect 15252 22176 15258 22228
rect 15746 22176 15752 22228
rect 15804 22216 15810 22228
rect 16006 22219 16064 22225
rect 16006 22216 16018 22219
rect 15804 22188 16018 22216
rect 15804 22176 15810 22188
rect 16006 22185 16018 22188
rect 16052 22185 16064 22219
rect 16006 22179 16064 22185
rect 16206 22176 16212 22228
rect 16264 22216 16270 22228
rect 16264 22188 18276 22216
rect 16264 22176 16270 22188
rect 9398 22108 9404 22160
rect 9456 22148 9462 22160
rect 12342 22148 12348 22160
rect 9456 22120 12348 22148
rect 9456 22108 9462 22120
rect 12342 22108 12348 22120
rect 12400 22108 12406 22160
rect 17402 22108 17408 22160
rect 17460 22148 17466 22160
rect 17770 22148 17776 22160
rect 17460 22120 17776 22148
rect 17460 22108 17466 22120
rect 17770 22108 17776 22120
rect 17828 22108 17834 22160
rect 18248 22148 18276 22188
rect 19978 22176 19984 22228
rect 20036 22216 20042 22228
rect 20606 22219 20664 22225
rect 20606 22216 20618 22219
rect 20036 22188 20618 22216
rect 20036 22176 20042 22188
rect 20606 22185 20618 22188
rect 20652 22185 20664 22219
rect 20606 22179 20664 22185
rect 20990 22176 20996 22228
rect 21048 22216 21054 22228
rect 24486 22216 24492 22228
rect 21048 22188 24492 22216
rect 21048 22176 21054 22188
rect 24486 22176 24492 22188
rect 24544 22176 24550 22228
rect 18248 22120 18368 22148
rect 1765 22083 1823 22089
rect 1765 22049 1777 22083
rect 1811 22080 1823 22083
rect 2498 22080 2504 22092
rect 1811 22052 2504 22080
rect 1811 22049 1823 22052
rect 1765 22043 1823 22049
rect 2498 22040 2504 22052
rect 2556 22040 2562 22092
rect 3237 22083 3295 22089
rect 3237 22049 3249 22083
rect 3283 22080 3295 22083
rect 3326 22080 3332 22092
rect 3283 22052 3332 22080
rect 3283 22049 3295 22052
rect 3237 22043 3295 22049
rect 3326 22040 3332 22052
rect 3384 22040 3390 22092
rect 3786 22040 3792 22092
rect 3844 22080 3850 22092
rect 7834 22080 7840 22092
rect 3844 22052 7840 22080
rect 3844 22040 3850 22052
rect 7834 22040 7840 22052
rect 7892 22040 7898 22092
rect 8113 22083 8171 22089
rect 8113 22049 8125 22083
rect 8159 22080 8171 22083
rect 8202 22080 8208 22106
rect 8159 22054 8208 22080
rect 8260 22094 8266 22106
rect 8260 22066 8339 22094
rect 8260 22054 8266 22066
rect 8159 22052 8248 22054
rect 8159 22049 8171 22052
rect 8113 22043 8171 22049
rect 8846 22040 8852 22092
rect 8904 22080 8910 22092
rect 9125 22083 9183 22089
rect 9125 22080 9137 22083
rect 8904 22052 9137 22080
rect 8904 22040 8910 22052
rect 9125 22049 9137 22052
rect 9171 22080 9183 22083
rect 9214 22080 9220 22092
rect 9171 22052 9220 22080
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 9214 22040 9220 22052
rect 9272 22040 9278 22092
rect 12618 22080 12624 22092
rect 9646 22052 12624 22080
rect 1854 21972 1860 22024
rect 1912 22012 1918 22024
rect 2041 22015 2099 22021
rect 2041 22012 2053 22015
rect 1912 21984 2053 22012
rect 1912 21972 1918 21984
rect 2041 21981 2053 21984
rect 2087 21981 2099 22015
rect 2041 21975 2099 21981
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 21981 4307 22015
rect 4249 21975 4307 21981
rect 3970 21904 3976 21956
rect 4028 21944 4034 21956
rect 4264 21944 4292 21975
rect 5442 21972 5448 22024
rect 5500 21972 5506 22024
rect 7282 22012 7288 22024
rect 5552 21984 7288 22012
rect 5552 21944 5580 21984
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 7374 21972 7380 22024
rect 7432 21972 7438 22024
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 22012 9551 22015
rect 9646 22012 9674 22052
rect 12618 22040 12624 22052
rect 12676 22040 12682 22092
rect 12986 22040 12992 22092
rect 13044 22040 13050 22092
rect 14826 22040 14832 22092
rect 14884 22040 14890 22092
rect 15749 22083 15807 22089
rect 15749 22049 15761 22083
rect 15795 22080 15807 22083
rect 17034 22080 17040 22092
rect 15795 22052 17040 22080
rect 15795 22049 15807 22052
rect 15749 22043 15807 22049
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 18046 22080 18052 22092
rect 17144 22052 18052 22080
rect 17144 22024 17172 22052
rect 18046 22040 18052 22052
rect 18104 22040 18110 22092
rect 18340 22080 18368 22120
rect 19058 22108 19064 22160
rect 19116 22148 19122 22160
rect 20346 22148 20352 22160
rect 19116 22120 20352 22148
rect 19116 22108 19122 22120
rect 20346 22108 20352 22120
rect 20404 22108 20410 22160
rect 25498 22148 25504 22160
rect 21744 22120 23520 22148
rect 18509 22083 18567 22089
rect 18509 22080 18521 22083
rect 18340 22052 18521 22080
rect 18509 22049 18521 22052
rect 18555 22049 18567 22083
rect 19426 22080 19432 22092
rect 18509 22043 18567 22049
rect 18708 22052 19432 22080
rect 9539 21984 9674 22012
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10597 22015 10655 22021
rect 10597 22012 10609 22015
rect 10100 21984 10609 22012
rect 10100 21972 10106 21984
rect 10597 21981 10609 21984
rect 10643 21981 10655 22015
rect 10597 21975 10655 21981
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 12805 22015 12863 22021
rect 12805 22012 12817 22015
rect 12492 21984 12817 22012
rect 12492 21972 12498 21984
rect 12805 21981 12817 21984
rect 12851 22012 12863 22015
rect 13633 22015 13691 22021
rect 13633 22012 13645 22015
rect 12851 21984 13645 22012
rect 12851 21981 12863 21984
rect 12805 21975 12863 21981
rect 13633 21981 13645 21984
rect 13679 21981 13691 22015
rect 14458 22012 14464 22024
rect 13633 21975 13691 21981
rect 13832 21984 14464 22012
rect 4028 21916 5580 21944
rect 4028 21904 4034 21916
rect 6086 21904 6092 21956
rect 6144 21944 6150 21956
rect 6273 21947 6331 21953
rect 6273 21944 6285 21947
rect 6144 21916 6285 21944
rect 6144 21904 6150 21916
rect 6273 21913 6285 21916
rect 6319 21913 6331 21947
rect 6273 21907 6331 21913
rect 6730 21904 6736 21956
rect 6788 21944 6794 21956
rect 10137 21947 10195 21953
rect 10137 21944 10149 21947
rect 6788 21916 10149 21944
rect 6788 21904 6794 21916
rect 10137 21913 10149 21916
rect 10183 21913 10195 21947
rect 10137 21907 10195 21913
rect 11054 21904 11060 21956
rect 11112 21944 11118 21956
rect 11517 21947 11575 21953
rect 11517 21944 11529 21947
rect 11112 21916 11529 21944
rect 11112 21904 11118 21916
rect 11517 21913 11529 21916
rect 11563 21913 11575 21947
rect 11517 21907 11575 21913
rect 12618 21904 12624 21956
rect 12676 21944 12682 21956
rect 13832 21944 13860 21984
rect 14458 21972 14464 21984
rect 14516 21972 14522 22024
rect 14645 22015 14703 22021
rect 14645 21981 14657 22015
rect 14691 22012 14703 22015
rect 15654 22012 15660 22024
rect 14691 21984 15660 22012
rect 14691 21981 14703 21984
rect 14645 21975 14703 21981
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 17126 21972 17132 22024
rect 17184 21972 17190 22024
rect 17862 21972 17868 22024
rect 17920 22012 17926 22024
rect 17920 21984 18092 22012
rect 17920 21972 17926 21984
rect 12676 21916 13860 21944
rect 13909 21947 13967 21953
rect 12676 21904 12682 21916
rect 13909 21913 13921 21947
rect 13955 21944 13967 21947
rect 14366 21944 14372 21956
rect 13955 21916 14372 21944
rect 13955 21913 13967 21916
rect 13909 21907 13967 21913
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 14737 21947 14795 21953
rect 14737 21913 14749 21947
rect 14783 21944 14795 21947
rect 18064 21944 18092 21984
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 18325 22015 18383 22021
rect 18325 22012 18337 22015
rect 18288 21984 18337 22012
rect 18288 21972 18294 21984
rect 18325 21981 18337 21984
rect 18371 21981 18383 22015
rect 18325 21975 18383 21981
rect 18414 21972 18420 22024
rect 18472 22012 18478 22024
rect 18708 22012 18736 22052
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 19518 22040 19524 22092
rect 19576 22080 19582 22092
rect 19705 22083 19763 22089
rect 19705 22080 19717 22083
rect 19576 22052 19717 22080
rect 19576 22040 19582 22052
rect 19705 22049 19717 22052
rect 19751 22049 19763 22083
rect 19705 22043 19763 22049
rect 18472 21984 18736 22012
rect 18472 21972 18478 21984
rect 19058 21972 19064 22024
rect 19116 22012 19122 22024
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 19116 21984 20361 22012
rect 19116 21972 19122 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 14783 21916 16436 21944
rect 14783 21913 14795 21916
rect 14737 21907 14795 21913
rect 3881 21879 3939 21885
rect 3881 21845 3893 21879
rect 3927 21876 3939 21879
rect 4614 21876 4620 21888
rect 3927 21848 4620 21876
rect 3927 21845 3939 21848
rect 3881 21839 3939 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 4893 21879 4951 21885
rect 4893 21845 4905 21879
rect 4939 21876 4951 21879
rect 4982 21876 4988 21888
rect 4939 21848 4988 21876
rect 4939 21845 4951 21848
rect 4893 21839 4951 21845
rect 4982 21836 4988 21848
rect 5040 21836 5046 21888
rect 5350 21836 5356 21888
rect 5408 21876 5414 21888
rect 8846 21876 8852 21888
rect 5408 21848 8852 21876
rect 5408 21836 5414 21848
rect 8846 21836 8852 21848
rect 8904 21836 8910 21888
rect 9030 21836 9036 21888
rect 9088 21836 9094 21888
rect 9214 21836 9220 21888
rect 9272 21876 9278 21888
rect 9674 21876 9680 21888
rect 9272 21848 9680 21876
rect 9272 21836 9278 21848
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 9858 21836 9864 21888
rect 9916 21876 9922 21888
rect 11146 21876 11152 21888
rect 9916 21848 11152 21876
rect 9916 21836 9922 21848
rect 11146 21836 11152 21848
rect 11204 21836 11210 21888
rect 12434 21836 12440 21888
rect 12492 21836 12498 21888
rect 12897 21879 12955 21885
rect 12897 21845 12909 21879
rect 12943 21876 12955 21879
rect 13998 21876 14004 21888
rect 12943 21848 14004 21876
rect 12943 21845 12955 21848
rect 12897 21839 12955 21845
rect 13998 21836 14004 21848
rect 14056 21836 14062 21888
rect 14274 21836 14280 21888
rect 14332 21836 14338 21888
rect 15286 21836 15292 21888
rect 15344 21836 15350 21888
rect 16408 21876 16436 21916
rect 17420 21916 18000 21944
rect 18064 21916 18552 21944
rect 17420 21876 17448 21916
rect 16408 21848 17448 21876
rect 17494 21836 17500 21888
rect 17552 21836 17558 21888
rect 17972 21885 18000 21916
rect 17957 21879 18015 21885
rect 17957 21845 17969 21879
rect 18003 21845 18015 21879
rect 17957 21839 18015 21845
rect 18138 21836 18144 21888
rect 18196 21876 18202 21888
rect 18417 21879 18475 21885
rect 18417 21876 18429 21879
rect 18196 21848 18429 21876
rect 18196 21836 18202 21848
rect 18417 21845 18429 21848
rect 18463 21845 18475 21879
rect 18524 21876 18552 21916
rect 18874 21904 18880 21956
rect 18932 21944 18938 21956
rect 19521 21947 19579 21953
rect 19521 21944 19533 21947
rect 18932 21916 19533 21944
rect 18932 21904 18938 21916
rect 19521 21913 19533 21916
rect 19567 21913 19579 21947
rect 19521 21907 19579 21913
rect 18969 21879 19027 21885
rect 18969 21876 18981 21879
rect 18524 21848 18981 21876
rect 18417 21839 18475 21845
rect 18969 21845 18981 21848
rect 19015 21845 19027 21879
rect 18969 21839 19027 21845
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19981 21879 20039 21885
rect 19981 21876 19993 21879
rect 19484 21848 19993 21876
rect 19484 21836 19490 21848
rect 19981 21845 19993 21848
rect 20027 21876 20039 21879
rect 20070 21876 20076 21888
rect 20027 21848 20076 21876
rect 20027 21845 20039 21848
rect 19981 21839 20039 21845
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 20714 21836 20720 21888
rect 20772 21876 20778 21888
rect 21744 21876 21772 22120
rect 23492 22092 23520 22120
rect 25148 22120 25504 22148
rect 22097 22083 22155 22089
rect 22097 22049 22109 22083
rect 22143 22080 22155 22083
rect 22143 22052 22876 22080
rect 22143 22049 22155 22052
rect 22097 22043 22155 22049
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22244 21984 22385 22012
rect 22244 21972 22250 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22848 22012 22876 22052
rect 23474 22040 23480 22092
rect 23532 22080 23538 22092
rect 25148 22089 25176 22120
rect 25498 22108 25504 22120
rect 25556 22108 25562 22160
rect 23845 22083 23903 22089
rect 23845 22080 23857 22083
rect 23532 22052 23857 22080
rect 23532 22040 23538 22052
rect 23845 22049 23857 22052
rect 23891 22049 23903 22083
rect 23845 22043 23903 22049
rect 25133 22083 25191 22089
rect 25133 22049 25145 22083
rect 25179 22049 25191 22083
rect 25133 22043 25191 22049
rect 23014 22012 23020 22024
rect 22848 21984 23020 22012
rect 22373 21975 22431 21981
rect 23014 21972 23020 21984
rect 23072 21972 23078 22024
rect 25041 22015 25099 22021
rect 25041 21981 25053 22015
rect 25087 22012 25099 22015
rect 25682 22012 25688 22024
rect 25087 21984 25688 22012
rect 25087 21981 25099 21984
rect 25041 21975 25099 21981
rect 25682 21972 25688 21984
rect 25740 21972 25746 22024
rect 22002 21904 22008 21956
rect 22060 21944 22066 21956
rect 22741 21947 22799 21953
rect 22741 21944 22753 21947
rect 22060 21916 22753 21944
rect 22060 21904 22066 21916
rect 22741 21913 22753 21916
rect 22787 21913 22799 21947
rect 22741 21907 22799 21913
rect 23106 21904 23112 21956
rect 23164 21904 23170 21956
rect 20772 21848 21772 21876
rect 20772 21836 20778 21848
rect 22278 21836 22284 21888
rect 22336 21876 22342 21888
rect 22557 21879 22615 21885
rect 22557 21876 22569 21879
rect 22336 21848 22569 21876
rect 22336 21836 22342 21848
rect 22557 21845 22569 21848
rect 22603 21845 22615 21879
rect 22557 21839 22615 21845
rect 24578 21836 24584 21888
rect 24636 21836 24642 21888
rect 24854 21836 24860 21888
rect 24912 21876 24918 21888
rect 24949 21879 25007 21885
rect 24949 21876 24961 21879
rect 24912 21848 24961 21876
rect 24912 21836 24918 21848
rect 24949 21845 24961 21848
rect 24995 21845 25007 21879
rect 24949 21839 25007 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 2317 21675 2375 21681
rect 2317 21641 2329 21675
rect 2363 21672 2375 21675
rect 4246 21672 4252 21684
rect 2363 21644 4252 21672
rect 2363 21641 2375 21644
rect 2317 21635 2375 21641
rect 4246 21632 4252 21644
rect 4304 21632 4310 21684
rect 4798 21632 4804 21684
rect 4856 21672 4862 21684
rect 5350 21672 5356 21684
rect 4856 21644 5356 21672
rect 4856 21632 4862 21644
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 5718 21632 5724 21684
rect 5776 21672 5782 21684
rect 5902 21672 5908 21684
rect 5776 21644 5908 21672
rect 5776 21632 5782 21644
rect 5902 21632 5908 21644
rect 5960 21632 5966 21684
rect 6086 21632 6092 21684
rect 6144 21672 6150 21684
rect 9214 21672 9220 21684
rect 6144 21644 9220 21672
rect 6144 21632 6150 21644
rect 9214 21632 9220 21644
rect 9272 21632 9278 21684
rect 11885 21675 11943 21681
rect 11885 21672 11897 21675
rect 9324 21644 11897 21672
rect 842 21564 848 21616
rect 900 21604 906 21616
rect 9324 21604 9352 21644
rect 11885 21641 11897 21644
rect 11931 21672 11943 21675
rect 12621 21675 12679 21681
rect 12621 21672 12633 21675
rect 11931 21644 12633 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12621 21641 12633 21644
rect 12667 21641 12679 21675
rect 12621 21635 12679 21641
rect 13906 21632 13912 21684
rect 13964 21672 13970 21684
rect 16482 21672 16488 21684
rect 13964 21644 16488 21672
rect 13964 21632 13970 21644
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 16853 21675 16911 21681
rect 16853 21641 16865 21675
rect 16899 21672 16911 21675
rect 17678 21672 17684 21684
rect 16899 21644 17684 21672
rect 16899 21641 16911 21644
rect 16853 21635 16911 21641
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 20438 21672 20444 21684
rect 17972 21644 18368 21672
rect 900 21576 9352 21604
rect 900 21564 906 21576
rect 11330 21564 11336 21616
rect 11388 21604 11394 21616
rect 11388 21576 12204 21604
rect 11388 21564 11394 21576
rect 1670 21496 1676 21548
rect 1728 21496 1734 21548
rect 2130 21496 2136 21548
rect 2188 21536 2194 21548
rect 2777 21539 2835 21545
rect 2777 21536 2789 21539
rect 2188 21508 2789 21536
rect 2188 21496 2194 21508
rect 2777 21505 2789 21508
rect 2823 21505 2835 21539
rect 2777 21499 2835 21505
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21505 4859 21539
rect 4801 21499 4859 21505
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 4816 21400 4844 21499
rect 5166 21496 5172 21548
rect 5224 21536 5230 21548
rect 7101 21539 7159 21545
rect 7101 21536 7113 21539
rect 5224 21508 7113 21536
rect 5224 21496 5230 21508
rect 7101 21505 7113 21508
rect 7147 21505 7159 21539
rect 7101 21499 7159 21505
rect 8938 21496 8944 21548
rect 8996 21496 9002 21548
rect 11054 21536 11060 21548
rect 10350 21508 11060 21536
rect 11054 21496 11060 21508
rect 11112 21536 11118 21548
rect 11241 21539 11299 21545
rect 11241 21536 11253 21539
rect 11112 21508 11253 21536
rect 11112 21496 11118 21508
rect 11241 21505 11253 21508
rect 11287 21536 11299 21539
rect 11974 21536 11980 21548
rect 11287 21508 11980 21536
rect 11287 21505 11299 21508
rect 11241 21499 11299 21505
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 5074 21428 5080 21480
rect 5132 21428 5138 21480
rect 5902 21428 5908 21480
rect 5960 21468 5966 21480
rect 6270 21468 6276 21480
rect 5960 21440 6276 21468
rect 5960 21428 5966 21440
rect 6270 21428 6276 21440
rect 6328 21468 6334 21480
rect 6733 21471 6791 21477
rect 6733 21468 6745 21471
rect 6328 21440 6745 21468
rect 6328 21428 6334 21440
rect 6733 21437 6745 21440
rect 6779 21437 6791 21471
rect 6733 21431 6791 21437
rect 6914 21428 6920 21480
rect 6972 21468 6978 21480
rect 7282 21468 7288 21480
rect 6972 21440 7288 21468
rect 6972 21428 6978 21440
rect 7282 21428 7288 21440
rect 7340 21428 7346 21480
rect 7466 21428 7472 21480
rect 7524 21468 7530 21480
rect 7561 21471 7619 21477
rect 7561 21468 7573 21471
rect 7524 21440 7573 21468
rect 7524 21428 7530 21440
rect 7561 21437 7573 21440
rect 7607 21437 7619 21471
rect 10962 21468 10968 21480
rect 7561 21431 7619 21437
rect 7668 21440 10968 21468
rect 7668 21400 7696 21440
rect 10962 21428 10968 21440
rect 11020 21428 11026 21480
rect 11606 21428 11612 21480
rect 11664 21468 11670 21480
rect 12066 21468 12072 21480
rect 11664 21440 12072 21468
rect 11664 21428 11670 21440
rect 12066 21428 12072 21440
rect 12124 21428 12130 21480
rect 12176 21468 12204 21576
rect 12250 21564 12256 21616
rect 12308 21604 12314 21616
rect 12986 21604 12992 21616
rect 12308 21576 12992 21604
rect 12308 21564 12314 21576
rect 12986 21564 12992 21576
rect 13044 21564 13050 21616
rect 13630 21604 13636 21616
rect 13464 21576 13636 21604
rect 13464 21545 13492 21576
rect 13630 21564 13636 21576
rect 13688 21564 13694 21616
rect 13722 21564 13728 21616
rect 13780 21564 13786 21616
rect 13998 21564 14004 21616
rect 14056 21604 14062 21616
rect 14056 21576 14214 21604
rect 14056 21564 14062 21576
rect 15102 21564 15108 21616
rect 15160 21604 15166 21616
rect 16390 21604 16396 21616
rect 15160 21576 16396 21604
rect 15160 21564 15166 21576
rect 16390 21564 16396 21576
rect 16448 21564 16454 21616
rect 17310 21564 17316 21616
rect 17368 21604 17374 21616
rect 17972 21604 18000 21644
rect 17368 21576 18000 21604
rect 18340 21604 18368 21644
rect 18524 21644 20444 21672
rect 18524 21604 18552 21644
rect 20438 21632 20444 21644
rect 20496 21632 20502 21684
rect 22002 21672 22008 21684
rect 21100 21644 22008 21672
rect 18340 21576 18552 21604
rect 17368 21564 17374 21576
rect 18598 21564 18604 21616
rect 18656 21564 18662 21616
rect 20162 21604 20168 21616
rect 19826 21576 20168 21604
rect 20162 21564 20168 21576
rect 20220 21564 20226 21616
rect 21100 21604 21128 21644
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22370 21632 22376 21684
rect 22428 21672 22434 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 22428 21644 22477 21672
rect 22428 21632 22434 21644
rect 22465 21641 22477 21644
rect 22511 21672 22523 21675
rect 23750 21672 23756 21684
rect 22511 21644 23756 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 23750 21632 23756 21644
rect 23808 21632 23814 21684
rect 23934 21632 23940 21684
rect 23992 21672 23998 21684
rect 24210 21672 24216 21684
rect 23992 21644 24216 21672
rect 23992 21632 23998 21644
rect 24210 21632 24216 21644
rect 24268 21672 24274 21684
rect 25409 21675 25467 21681
rect 25409 21672 25421 21675
rect 24268 21644 25421 21672
rect 24268 21632 24274 21644
rect 25409 21641 25421 21644
rect 25455 21641 25467 21675
rect 25409 21635 25467 21641
rect 21634 21604 21640 21616
rect 20272 21576 21128 21604
rect 21192 21576 21640 21604
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 15657 21539 15715 21545
rect 15657 21505 15669 21539
rect 15703 21536 15715 21539
rect 15703 21508 16436 21536
rect 15703 21505 15715 21508
rect 15657 21499 15715 21505
rect 12618 21468 12624 21480
rect 12176 21440 12624 21468
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 12710 21428 12716 21480
rect 12768 21428 12774 21480
rect 12897 21471 12955 21477
rect 12897 21437 12909 21471
rect 12943 21468 12955 21471
rect 12943 21440 13492 21468
rect 12943 21437 12955 21440
rect 12897 21431 12955 21437
rect 13464 21412 13492 21440
rect 14366 21428 14372 21480
rect 14424 21468 14430 21480
rect 16022 21468 16028 21480
rect 14424 21440 16028 21468
rect 14424 21428 14430 21440
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 4816 21372 7696 21400
rect 10612 21372 13400 21400
rect 1302 21292 1308 21344
rect 1360 21332 1366 21344
rect 6086 21332 6092 21344
rect 1360 21304 6092 21332
rect 1360 21292 1366 21304
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 6454 21292 6460 21344
rect 6512 21292 6518 21344
rect 6638 21292 6644 21344
rect 6696 21292 6702 21344
rect 7558 21292 7564 21344
rect 7616 21332 7622 21344
rect 9198 21335 9256 21341
rect 9198 21332 9210 21335
rect 7616 21304 9210 21332
rect 7616 21292 7622 21304
rect 9198 21301 9210 21304
rect 9244 21301 9256 21335
rect 9198 21295 9256 21301
rect 9582 21292 9588 21344
rect 9640 21332 9646 21344
rect 10612 21332 10640 21372
rect 9640 21304 10640 21332
rect 9640 21292 9646 21304
rect 10686 21292 10692 21344
rect 10744 21292 10750 21344
rect 11606 21292 11612 21344
rect 11664 21292 11670 21344
rect 11698 21292 11704 21344
rect 11756 21292 11762 21344
rect 12066 21292 12072 21344
rect 12124 21332 12130 21344
rect 12253 21335 12311 21341
rect 12253 21332 12265 21335
rect 12124 21304 12265 21332
rect 12124 21292 12130 21304
rect 12253 21301 12265 21304
rect 12299 21301 12311 21335
rect 13372 21332 13400 21372
rect 13446 21360 13452 21412
rect 13504 21360 13510 21412
rect 16206 21400 16212 21412
rect 15212 21372 16212 21400
rect 15212 21341 15240 21372
rect 16206 21360 16212 21372
rect 16264 21360 16270 21412
rect 15197 21335 15255 21341
rect 15197 21332 15209 21335
rect 13372 21304 15209 21332
rect 12253 21295 12311 21301
rect 15197 21301 15209 21304
rect 15243 21301 15255 21335
rect 15197 21295 15255 21301
rect 15286 21292 15292 21344
rect 15344 21332 15350 21344
rect 16301 21335 16359 21341
rect 16301 21332 16313 21335
rect 15344 21304 16313 21332
rect 15344 21292 15350 21304
rect 16301 21301 16313 21304
rect 16347 21301 16359 21335
rect 16408 21332 16436 21508
rect 17218 21496 17224 21548
rect 17276 21536 17282 21548
rect 18230 21536 18236 21548
rect 17276 21508 18236 21536
rect 17276 21496 17282 21508
rect 18230 21496 18236 21508
rect 18288 21496 18294 21548
rect 18322 21496 18328 21548
rect 18380 21496 18386 21548
rect 20272 21536 20300 21576
rect 19812 21508 20300 21536
rect 21085 21539 21143 21545
rect 16482 21428 16488 21480
rect 16540 21468 16546 21480
rect 16942 21468 16948 21480
rect 16540 21440 16948 21468
rect 16540 21428 16546 21440
rect 16942 21428 16948 21440
rect 17000 21468 17006 21480
rect 17313 21471 17371 21477
rect 17313 21468 17325 21471
rect 17000 21440 17325 21468
rect 17000 21428 17006 21440
rect 17313 21437 17325 21440
rect 17359 21437 17371 21471
rect 17313 21431 17371 21437
rect 17402 21428 17408 21480
rect 17460 21468 17466 21480
rect 17865 21471 17923 21477
rect 17865 21468 17877 21471
rect 17460 21440 17877 21468
rect 17460 21428 17466 21440
rect 17865 21437 17877 21440
rect 17911 21468 17923 21471
rect 17911 21440 19748 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 19720 21412 19748 21440
rect 17034 21360 17040 21412
rect 17092 21400 17098 21412
rect 18322 21400 18328 21412
rect 17092 21372 18328 21400
rect 17092 21360 17098 21372
rect 18322 21360 18328 21372
rect 18380 21360 18386 21412
rect 19702 21360 19708 21412
rect 19760 21360 19766 21412
rect 17862 21332 17868 21344
rect 16408 21304 17868 21332
rect 16301 21295 16359 21301
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 18966 21292 18972 21344
rect 19024 21332 19030 21344
rect 19812 21332 19840 21508
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 21192 21536 21220 21576
rect 21634 21564 21640 21576
rect 21692 21564 21698 21616
rect 23566 21564 23572 21616
rect 23624 21564 23630 21616
rect 23952 21604 23980 21632
rect 23952 21576 24058 21604
rect 21450 21536 21456 21548
rect 21131 21508 21220 21536
rect 21284 21508 21456 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 20070 21428 20076 21480
rect 20128 21428 20134 21480
rect 21174 21428 21180 21480
rect 21232 21428 21238 21480
rect 21284 21477 21312 21508
rect 21450 21496 21456 21508
rect 21508 21496 21514 21548
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22152 21508 22692 21536
rect 22152 21496 22158 21508
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21437 21327 21471
rect 21269 21431 21327 21437
rect 21358 21428 21364 21480
rect 21416 21468 21422 21480
rect 22278 21468 22284 21480
rect 21416 21440 22284 21468
rect 21416 21428 21422 21440
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 22554 21428 22560 21480
rect 22612 21428 22618 21480
rect 22664 21477 22692 21508
rect 23290 21496 23296 21548
rect 23348 21496 23354 21548
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 23014 21428 23020 21480
rect 23072 21468 23078 21480
rect 23566 21468 23572 21480
rect 23072 21440 23572 21468
rect 23072 21428 23078 21440
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 19886 21360 19892 21412
rect 19944 21400 19950 21412
rect 21726 21400 21732 21412
rect 19944 21372 21732 21400
rect 19944 21360 19950 21372
rect 21726 21360 21732 21372
rect 21784 21360 21790 21412
rect 21818 21360 21824 21412
rect 21876 21400 21882 21412
rect 23106 21400 23112 21412
rect 21876 21372 23112 21400
rect 21876 21360 21882 21372
rect 23106 21360 23112 21372
rect 23164 21360 23170 21412
rect 25590 21360 25596 21412
rect 25648 21400 25654 21412
rect 26050 21400 26056 21412
rect 25648 21372 26056 21400
rect 25648 21360 25654 21372
rect 26050 21360 26056 21372
rect 26108 21360 26114 21412
rect 19024 21304 19840 21332
rect 19024 21292 19030 21304
rect 20162 21292 20168 21344
rect 20220 21332 20226 21344
rect 20349 21335 20407 21341
rect 20349 21332 20361 21335
rect 20220 21304 20361 21332
rect 20220 21292 20226 21304
rect 20349 21301 20361 21304
rect 20395 21301 20407 21335
rect 20349 21295 20407 21301
rect 20717 21335 20775 21341
rect 20717 21301 20729 21335
rect 20763 21332 20775 21335
rect 21542 21332 21548 21344
rect 20763 21304 21548 21332
rect 20763 21301 20775 21304
rect 20717 21295 20775 21301
rect 21542 21292 21548 21304
rect 21600 21292 21606 21344
rect 22097 21335 22155 21341
rect 22097 21301 22109 21335
rect 22143 21332 22155 21335
rect 23382 21332 23388 21344
rect 22143 21304 23388 21332
rect 22143 21301 22155 21304
rect 22097 21295 22155 21301
rect 23382 21292 23388 21304
rect 23440 21292 23446 21344
rect 25041 21335 25099 21341
rect 25041 21301 25053 21335
rect 25087 21332 25099 21335
rect 25314 21332 25320 21344
rect 25087 21304 25320 21332
rect 25087 21301 25099 21304
rect 25041 21295 25099 21301
rect 25314 21292 25320 21304
rect 25372 21332 25378 21344
rect 25498 21332 25504 21344
rect 25372 21304 25504 21332
rect 25372 21292 25378 21304
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 1765 21131 1823 21137
rect 1765 21097 1777 21131
rect 1811 21128 1823 21131
rect 3970 21128 3976 21140
rect 1811 21100 3976 21128
rect 1811 21097 1823 21100
rect 1765 21091 1823 21097
rect 3970 21088 3976 21100
rect 4028 21088 4034 21140
rect 6457 21131 6515 21137
rect 6457 21097 6469 21131
rect 6503 21128 6515 21131
rect 6822 21128 6828 21140
rect 6503 21100 6828 21128
rect 6503 21097 6515 21100
rect 6457 21091 6515 21097
rect 6822 21088 6828 21100
rect 6880 21088 6886 21140
rect 7374 21088 7380 21140
rect 7432 21128 7438 21140
rect 9401 21131 9459 21137
rect 9401 21128 9413 21131
rect 7432 21100 9413 21128
rect 7432 21088 7438 21100
rect 9401 21097 9413 21100
rect 9447 21097 9459 21131
rect 15289 21131 15347 21137
rect 15289 21128 15301 21131
rect 9401 21091 9459 21097
rect 10520 21100 15301 21128
rect 1581 21063 1639 21069
rect 1581 21029 1593 21063
rect 1627 21060 1639 21063
rect 3326 21060 3332 21072
rect 1627 21032 3332 21060
rect 1627 21029 1639 21032
rect 1581 21023 1639 21029
rect 3326 21020 3332 21032
rect 3384 21060 3390 21072
rect 5718 21060 5724 21072
rect 3384 21032 5724 21060
rect 3384 21020 3390 21032
rect 5718 21020 5724 21032
rect 5776 21020 5782 21072
rect 10042 21060 10048 21072
rect 6932 21032 10048 21060
rect 2774 20952 2780 21004
rect 2832 20952 2838 21004
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 4614 20952 4620 21004
rect 4672 20992 4678 21004
rect 6822 20992 6828 21004
rect 4672 20964 6828 20992
rect 4672 20952 4678 20964
rect 6822 20952 6828 20964
rect 6880 20952 6886 21004
rect 2222 20884 2228 20936
rect 2280 20884 2286 20936
rect 4062 20884 4068 20936
rect 4120 20884 4126 20936
rect 5813 20927 5871 20933
rect 5813 20893 5825 20927
rect 5859 20893 5871 20927
rect 5813 20887 5871 20893
rect 2498 20816 2504 20868
rect 2556 20856 2562 20868
rect 4706 20856 4712 20868
rect 2556 20828 4712 20856
rect 2556 20816 2562 20828
rect 4706 20816 4712 20828
rect 4764 20816 4770 20868
rect 5828 20856 5856 20887
rect 6454 20884 6460 20936
rect 6512 20924 6518 20936
rect 6932 20924 6960 21032
rect 10042 21020 10048 21032
rect 10100 21020 10106 21072
rect 10520 21060 10548 21100
rect 15289 21097 15301 21100
rect 15335 21097 15347 21131
rect 15289 21091 15347 21097
rect 15654 21088 15660 21140
rect 15712 21128 15718 21140
rect 18598 21128 18604 21140
rect 15712 21100 18604 21128
rect 15712 21088 15718 21100
rect 18598 21088 18604 21100
rect 18656 21088 18662 21140
rect 18690 21088 18696 21140
rect 18748 21128 18754 21140
rect 21358 21128 21364 21140
rect 18748 21100 21364 21128
rect 18748 21088 18754 21100
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 21468 21100 22232 21128
rect 10428 21032 10548 21060
rect 7282 20952 7288 21004
rect 7340 20992 7346 21004
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 7340 20964 7389 20992
rect 7340 20952 7346 20964
rect 7377 20961 7389 20964
rect 7423 20961 7435 20995
rect 9582 20992 9588 21004
rect 7377 20955 7435 20961
rect 8680 20964 9588 20992
rect 6512 20896 6960 20924
rect 7101 20927 7159 20933
rect 6512 20884 6518 20896
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7742 20924 7748 20936
rect 7147 20896 7748 20924
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7742 20884 7748 20896
rect 7800 20884 7806 20936
rect 8680 20856 8708 20964
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 10428 21001 10456 21032
rect 12710 21020 12716 21072
rect 12768 21060 12774 21072
rect 16485 21063 16543 21069
rect 16485 21060 16497 21063
rect 12768 21032 16497 21060
rect 12768 21020 12774 21032
rect 16485 21029 16497 21032
rect 16531 21029 16543 21063
rect 17218 21060 17224 21072
rect 16485 21023 16543 21029
rect 16592 21032 17224 21060
rect 9769 20995 9827 21001
rect 9769 20992 9781 20995
rect 9732 20964 9781 20992
rect 9732 20952 9738 20964
rect 9769 20961 9781 20964
rect 9815 20992 9827 20995
rect 10413 20995 10471 21001
rect 9815 20964 10364 20992
rect 9815 20961 9827 20964
rect 9769 20955 9827 20961
rect 8754 20884 8760 20936
rect 8812 20924 8818 20936
rect 10336 20933 10364 20964
rect 10413 20961 10425 20995
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 10594 20952 10600 21004
rect 10652 20952 10658 21004
rect 11149 20995 11207 21001
rect 11149 20961 11161 20995
rect 11195 20992 11207 20995
rect 11514 20992 11520 21004
rect 11195 20964 11520 20992
rect 11195 20961 11207 20964
rect 11149 20955 11207 20961
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 12618 20952 12624 21004
rect 12676 20992 12682 21004
rect 15841 20995 15899 21001
rect 15841 20992 15853 20995
rect 12676 20964 15853 20992
rect 12676 20952 12682 20964
rect 15841 20961 15853 20964
rect 15887 20961 15899 20995
rect 15841 20955 15899 20961
rect 9309 20927 9367 20933
rect 9309 20924 9321 20927
rect 8812 20896 9321 20924
rect 8812 20884 8818 20896
rect 9309 20893 9321 20896
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 13538 20884 13544 20936
rect 13596 20884 13602 20936
rect 13722 20884 13728 20936
rect 13780 20884 13786 20936
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 13832 20896 14289 20924
rect 11425 20859 11483 20865
rect 11425 20856 11437 20859
rect 5828 20828 8708 20856
rect 9416 20828 11437 20856
rect 2038 20748 2044 20800
rect 2096 20788 2102 20800
rect 2774 20788 2780 20800
rect 2096 20760 2780 20788
rect 2096 20748 2102 20760
rect 2774 20748 2780 20760
rect 2832 20748 2838 20800
rect 3510 20748 3516 20800
rect 3568 20788 3574 20800
rect 5534 20788 5540 20800
rect 3568 20760 5540 20788
rect 3568 20748 3574 20760
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 5994 20748 6000 20800
rect 6052 20788 6058 20800
rect 9416 20788 9444 20828
rect 11425 20825 11437 20828
rect 11471 20825 11483 20859
rect 12710 20856 12716 20868
rect 12650 20828 12716 20856
rect 11425 20819 11483 20825
rect 12710 20816 12716 20828
rect 12768 20856 12774 20868
rect 13170 20856 13176 20868
rect 12768 20828 13176 20856
rect 12768 20816 12774 20828
rect 13170 20816 13176 20828
rect 13228 20816 13234 20868
rect 13262 20816 13268 20868
rect 13320 20856 13326 20868
rect 13832 20856 13860 20896
rect 14277 20893 14289 20896
rect 14323 20924 14335 20927
rect 14366 20924 14372 20936
rect 14323 20896 14372 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 14516 20896 15332 20924
rect 14516 20884 14522 20896
rect 13320 20828 13860 20856
rect 13320 20816 13326 20828
rect 13998 20816 14004 20868
rect 14056 20856 14062 20868
rect 14553 20859 14611 20865
rect 14553 20856 14565 20859
rect 14056 20828 14565 20856
rect 14056 20816 14062 20828
rect 14553 20825 14565 20828
rect 14599 20825 14611 20859
rect 15304 20856 15332 20896
rect 15378 20884 15384 20936
rect 15436 20924 15442 20936
rect 15657 20927 15715 20933
rect 15657 20924 15669 20927
rect 15436 20896 15669 20924
rect 15436 20884 15442 20896
rect 15657 20893 15669 20896
rect 15703 20893 15715 20927
rect 15657 20887 15715 20893
rect 15749 20927 15807 20933
rect 15749 20893 15761 20927
rect 15795 20924 15807 20927
rect 16022 20924 16028 20936
rect 15795 20896 16028 20924
rect 15795 20893 15807 20896
rect 15749 20887 15807 20893
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 16592 20924 16620 21032
rect 17218 21020 17224 21032
rect 17276 21020 17282 21072
rect 19242 21060 19248 21072
rect 18248 21032 19248 21060
rect 17037 20995 17095 21001
rect 17037 20992 17049 20995
rect 16540 20896 16620 20924
rect 16684 20964 17049 20992
rect 16540 20884 16546 20896
rect 16684 20856 16712 20964
rect 17037 20961 17049 20964
rect 17083 20961 17095 20995
rect 17037 20955 17095 20961
rect 17770 20952 17776 21004
rect 17828 20992 17834 21004
rect 18248 21001 18276 21032
rect 19242 21020 19248 21032
rect 19300 21020 19306 21072
rect 21177 21063 21235 21069
rect 21177 21029 21189 21063
rect 21223 21060 21235 21063
rect 21266 21060 21272 21072
rect 21223 21032 21272 21060
rect 21223 21029 21235 21032
rect 21177 21023 21235 21029
rect 21266 21020 21272 21032
rect 21324 21020 21330 21072
rect 18141 20995 18199 21001
rect 18141 20992 18153 20995
rect 17828 20964 18153 20992
rect 17828 20952 17834 20964
rect 18141 20961 18153 20964
rect 18187 20961 18199 20995
rect 18141 20955 18199 20961
rect 18233 20995 18291 21001
rect 18233 20961 18245 20995
rect 18279 20961 18291 20995
rect 18233 20955 18291 20961
rect 18322 20952 18328 21004
rect 18380 20992 18386 21004
rect 19058 20992 19064 21004
rect 18380 20964 19064 20992
rect 18380 20952 18386 20964
rect 19058 20952 19064 20964
rect 19116 20992 19122 21004
rect 19429 20995 19487 21001
rect 19429 20992 19441 20995
rect 19116 20964 19441 20992
rect 19116 20952 19122 20964
rect 19429 20961 19441 20964
rect 19475 20992 19487 20995
rect 20254 20992 20260 21004
rect 19475 20964 20260 20992
rect 19475 20961 19487 20964
rect 19429 20955 19487 20961
rect 20254 20952 20260 20964
rect 20312 20952 20318 21004
rect 20438 20952 20444 21004
rect 20496 20992 20502 21004
rect 21468 20992 21496 21100
rect 21545 21063 21603 21069
rect 21545 21029 21557 21063
rect 21591 21060 21603 21063
rect 21634 21060 21640 21072
rect 21591 21032 21640 21060
rect 21591 21029 21603 21032
rect 21545 21023 21603 21029
rect 21634 21020 21640 21032
rect 21692 21020 21698 21072
rect 22204 21060 22232 21100
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 25222 21128 25228 21140
rect 22336 21100 25228 21128
rect 22336 21088 22342 21100
rect 25222 21088 25228 21100
rect 25280 21088 25286 21140
rect 24581 21063 24639 21069
rect 22204 21032 23980 21060
rect 20496 20964 21496 20992
rect 21652 20992 21680 21020
rect 22462 20992 22468 21004
rect 21652 20964 22468 20992
rect 20496 20952 20502 20964
rect 22462 20952 22468 20964
rect 22520 20952 22526 21004
rect 22741 20995 22799 21001
rect 22741 20961 22753 20995
rect 22787 20992 22799 20995
rect 22922 20992 22928 21004
rect 22787 20964 22928 20992
rect 22787 20961 22799 20964
rect 22741 20955 22799 20961
rect 22922 20952 22928 20964
rect 22980 20952 22986 21004
rect 23566 20952 23572 21004
rect 23624 20992 23630 21004
rect 23845 20995 23903 21001
rect 23845 20992 23857 20995
rect 23624 20964 23857 20992
rect 23624 20952 23630 20964
rect 23845 20961 23857 20964
rect 23891 20961 23903 20995
rect 23845 20955 23903 20961
rect 16942 20884 16948 20936
rect 17000 20884 17006 20936
rect 21358 20884 21364 20936
rect 21416 20924 21422 20936
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 21416 20896 23765 20924
rect 21416 20884 21422 20896
rect 23753 20893 23765 20896
rect 23799 20893 23811 20927
rect 23753 20887 23811 20893
rect 15304 20828 16712 20856
rect 14553 20819 14611 20825
rect 16758 20816 16764 20868
rect 16816 20856 16822 20868
rect 16816 20828 18092 20856
rect 16816 20816 16822 20828
rect 6052 20760 9444 20788
rect 6052 20748 6058 20760
rect 9950 20748 9956 20800
rect 10008 20748 10014 20800
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 12897 20791 12955 20797
rect 12897 20788 12909 20791
rect 11204 20760 12909 20788
rect 11204 20748 11210 20760
rect 12897 20757 12909 20760
rect 12943 20788 12955 20791
rect 15838 20788 15844 20800
rect 12943 20760 15844 20788
rect 12943 20757 12955 20760
rect 12897 20751 12955 20757
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 16850 20748 16856 20800
rect 16908 20748 16914 20800
rect 17678 20748 17684 20800
rect 17736 20748 17742 20800
rect 18064 20797 18092 20828
rect 18230 20816 18236 20868
rect 18288 20856 18294 20868
rect 18693 20859 18751 20865
rect 18693 20856 18705 20859
rect 18288 20828 18705 20856
rect 18288 20816 18294 20828
rect 18693 20825 18705 20828
rect 18739 20825 18751 20859
rect 18693 20819 18751 20825
rect 18984 20828 19334 20856
rect 18049 20791 18107 20797
rect 18049 20757 18061 20791
rect 18095 20788 18107 20791
rect 18984 20788 19012 20828
rect 18095 20760 19012 20788
rect 18095 20757 18107 20760
rect 18049 20751 18107 20757
rect 19058 20748 19064 20800
rect 19116 20748 19122 20800
rect 19306 20788 19334 20828
rect 19702 20816 19708 20868
rect 19760 20816 19766 20868
rect 20714 20816 20720 20868
rect 20772 20816 20778 20868
rect 23952 20856 23980 21032
rect 24581 21029 24593 21063
rect 24627 21060 24639 21063
rect 24670 21060 24676 21072
rect 24627 21032 24676 21060
rect 24627 21029 24639 21032
rect 24581 21023 24639 21029
rect 24670 21020 24676 21032
rect 24728 21020 24734 21072
rect 24946 21020 24952 21072
rect 25004 21020 25010 21072
rect 24964 20992 24992 21020
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 24964 20964 25145 20992
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 24578 20884 24584 20936
rect 24636 20924 24642 20936
rect 24949 20927 25007 20933
rect 24949 20924 24961 20927
rect 24636 20896 24961 20924
rect 24636 20884 24642 20896
rect 24949 20893 24961 20896
rect 24995 20893 25007 20927
rect 24949 20887 25007 20893
rect 25041 20859 25099 20865
rect 25041 20856 25053 20859
rect 22204 20828 23888 20856
rect 23952 20828 25053 20856
rect 21634 20788 21640 20800
rect 19306 20760 21640 20788
rect 21634 20748 21640 20760
rect 21692 20748 21698 20800
rect 21726 20748 21732 20800
rect 21784 20748 21790 20800
rect 22097 20791 22155 20797
rect 22097 20757 22109 20791
rect 22143 20788 22155 20791
rect 22204 20788 22232 20828
rect 22143 20760 22232 20788
rect 22143 20757 22155 20760
rect 22097 20751 22155 20757
rect 22278 20748 22284 20800
rect 22336 20788 22342 20800
rect 22465 20791 22523 20797
rect 22465 20788 22477 20791
rect 22336 20760 22477 20788
rect 22336 20748 22342 20760
rect 22465 20757 22477 20760
rect 22511 20757 22523 20791
rect 22465 20751 22523 20757
rect 22554 20748 22560 20800
rect 22612 20748 22618 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 22704 20760 23305 20788
rect 22704 20748 22710 20760
rect 23293 20757 23305 20760
rect 23339 20757 23351 20791
rect 23293 20751 23351 20757
rect 23658 20748 23664 20800
rect 23716 20748 23722 20800
rect 23860 20788 23888 20828
rect 25041 20825 25053 20828
rect 25087 20825 25099 20859
rect 25041 20819 25099 20825
rect 25406 20788 25412 20800
rect 23860 20760 25412 20788
rect 25406 20748 25412 20760
rect 25464 20748 25470 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 1489 20587 1547 20593
rect 1489 20553 1501 20587
rect 1535 20584 1547 20587
rect 4430 20584 4436 20596
rect 1535 20556 4436 20584
rect 1535 20553 1547 20556
rect 1489 20547 1547 20553
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 4706 20544 4712 20596
rect 4764 20544 4770 20596
rect 5994 20544 6000 20596
rect 6052 20544 6058 20596
rect 8478 20544 8484 20596
rect 8536 20544 8542 20596
rect 9600 20556 13952 20584
rect 7282 20516 7288 20528
rect 1780 20488 7288 20516
rect 1780 20457 1808 20488
rect 7282 20476 7288 20488
rect 7340 20476 7346 20528
rect 7377 20519 7435 20525
rect 7377 20485 7389 20519
rect 7423 20516 7435 20519
rect 9600 20516 9628 20556
rect 11054 20516 11060 20528
rect 7423 20488 9628 20516
rect 10442 20488 11060 20516
rect 7423 20485 7435 20488
rect 7377 20479 7435 20485
rect 11054 20476 11060 20488
rect 11112 20476 11118 20528
rect 11238 20476 11244 20528
rect 11296 20516 11302 20528
rect 12437 20519 12495 20525
rect 12437 20516 12449 20519
rect 11296 20488 12449 20516
rect 11296 20476 11302 20488
rect 12437 20485 12449 20488
rect 12483 20485 12495 20519
rect 12437 20479 12495 20485
rect 13262 20476 13268 20528
rect 13320 20476 13326 20528
rect 13538 20516 13544 20528
rect 13372 20488 13544 20516
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20417 1823 20451
rect 1765 20411 1823 20417
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20448 3111 20451
rect 4893 20451 4951 20457
rect 3099 20420 4292 20448
rect 3099 20417 3111 20420
rect 3053 20411 3111 20417
rect 2958 20340 2964 20392
rect 3016 20380 3022 20392
rect 3329 20383 3387 20389
rect 3329 20380 3341 20383
rect 3016 20352 3341 20380
rect 3016 20340 3022 20352
rect 3329 20349 3341 20352
rect 3375 20349 3387 20383
rect 4264 20380 4292 20420
rect 4893 20417 4905 20451
rect 4939 20448 4951 20451
rect 5074 20448 5080 20460
rect 4939 20420 5080 20448
rect 4939 20417 4951 20420
rect 4893 20411 4951 20417
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20448 5411 20451
rect 5994 20448 6000 20460
rect 5399 20420 6000 20448
rect 5399 20417 5411 20420
rect 5353 20411 5411 20417
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 6733 20451 6791 20457
rect 6733 20448 6745 20451
rect 6604 20420 6745 20448
rect 6604 20408 6610 20420
rect 6733 20417 6745 20420
rect 6779 20417 6791 20451
rect 6733 20411 6791 20417
rect 7834 20408 7840 20460
rect 7892 20408 7898 20460
rect 8938 20408 8944 20460
rect 8996 20408 9002 20460
rect 10962 20408 10968 20460
rect 11020 20448 11026 20460
rect 11020 20420 12940 20448
rect 11020 20408 11026 20420
rect 5626 20380 5632 20392
rect 4264 20352 5632 20380
rect 3329 20343 3387 20349
rect 5626 20340 5632 20352
rect 5684 20340 5690 20392
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 9217 20383 9275 20389
rect 9217 20380 9229 20383
rect 8352 20352 9229 20380
rect 8352 20340 8358 20352
rect 9217 20349 9229 20352
rect 9263 20349 9275 20383
rect 9217 20343 9275 20349
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 11241 20383 11299 20389
rect 11241 20380 11253 20383
rect 9732 20352 11253 20380
rect 9732 20340 9738 20352
rect 11241 20349 11253 20352
rect 11287 20380 11299 20383
rect 12529 20383 12587 20389
rect 11287 20352 12434 20380
rect 11287 20349 11299 20352
rect 11241 20343 11299 20349
rect 2314 20272 2320 20324
rect 2372 20312 2378 20324
rect 3694 20312 3700 20324
rect 2372 20284 3700 20312
rect 2372 20272 2378 20284
rect 3694 20272 3700 20284
rect 3752 20272 3758 20324
rect 3970 20272 3976 20324
rect 4028 20312 4034 20324
rect 8846 20312 8852 20324
rect 4028 20284 8852 20312
rect 4028 20272 4034 20284
rect 8846 20272 8852 20284
rect 8904 20272 8910 20324
rect 11609 20315 11667 20321
rect 10244 20284 11284 20312
rect 2409 20247 2467 20253
rect 2409 20213 2421 20247
rect 2455 20244 2467 20247
rect 4246 20244 4252 20256
rect 2455 20216 4252 20244
rect 2455 20213 2467 20216
rect 2409 20207 2467 20213
rect 4246 20204 4252 20216
rect 4304 20204 4310 20256
rect 5074 20204 5080 20256
rect 5132 20244 5138 20256
rect 6457 20247 6515 20253
rect 6457 20244 6469 20247
rect 5132 20216 6469 20244
rect 5132 20204 5138 20216
rect 6457 20213 6469 20216
rect 6503 20244 6515 20247
rect 6546 20244 6552 20256
rect 6503 20216 6552 20244
rect 6503 20213 6515 20216
rect 6457 20207 6515 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 7834 20204 7840 20256
rect 7892 20244 7898 20256
rect 10244 20244 10272 20284
rect 11256 20256 11284 20284
rect 11609 20281 11621 20315
rect 11655 20312 11667 20315
rect 11974 20312 11980 20324
rect 11655 20284 11980 20312
rect 11655 20281 11667 20284
rect 11609 20275 11667 20281
rect 11974 20272 11980 20284
rect 12032 20272 12038 20324
rect 7892 20216 10272 20244
rect 7892 20204 7898 20216
rect 10502 20204 10508 20256
rect 10560 20244 10566 20256
rect 10689 20247 10747 20253
rect 10689 20244 10701 20247
rect 10560 20216 10701 20244
rect 10560 20204 10566 20216
rect 10689 20213 10701 20216
rect 10735 20213 10747 20247
rect 10689 20207 10747 20213
rect 11238 20204 11244 20256
rect 11296 20204 11302 20256
rect 11698 20204 11704 20256
rect 11756 20204 11762 20256
rect 12066 20204 12072 20256
rect 12124 20204 12130 20256
rect 12406 20244 12434 20352
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 12544 20312 12572 20343
rect 12618 20340 12624 20392
rect 12676 20340 12682 20392
rect 12912 20380 12940 20420
rect 13170 20408 13176 20460
rect 13228 20448 13234 20460
rect 13372 20448 13400 20488
rect 13538 20476 13544 20488
rect 13596 20476 13602 20528
rect 13924 20525 13952 20556
rect 15378 20544 15384 20596
rect 15436 20544 15442 20596
rect 15948 20556 20576 20584
rect 13909 20519 13967 20525
rect 13909 20485 13921 20519
rect 13955 20485 13967 20519
rect 13909 20479 13967 20485
rect 13998 20476 14004 20528
rect 14056 20516 14062 20528
rect 15948 20525 15976 20556
rect 15933 20519 15991 20525
rect 14056 20488 14398 20516
rect 14056 20476 14062 20488
rect 15933 20485 15945 20519
rect 15979 20485 15991 20519
rect 15933 20479 15991 20485
rect 16482 20476 16488 20528
rect 16540 20476 16546 20528
rect 16761 20519 16819 20525
rect 16761 20485 16773 20519
rect 16807 20516 16819 20519
rect 16942 20516 16948 20528
rect 16807 20488 16948 20516
rect 16807 20485 16819 20488
rect 16761 20479 16819 20485
rect 16942 20476 16948 20488
rect 17000 20476 17006 20528
rect 20162 20516 20168 20528
rect 18630 20488 20168 20516
rect 13630 20448 13636 20460
rect 13688 20457 13694 20460
rect 13228 20420 13400 20448
rect 13598 20420 13636 20448
rect 13228 20408 13234 20420
rect 13630 20408 13636 20420
rect 13688 20411 13698 20457
rect 13688 20408 13694 20411
rect 17034 20408 17040 20460
rect 17092 20448 17098 20460
rect 17129 20451 17187 20457
rect 17129 20448 17141 20451
rect 17092 20420 17141 20448
rect 17092 20408 17098 20420
rect 17129 20417 17141 20420
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 16117 20383 16175 20389
rect 16117 20380 16129 20383
rect 12912 20352 16129 20380
rect 16117 20349 16129 20352
rect 16163 20349 16175 20383
rect 16117 20343 16175 20349
rect 17402 20340 17408 20392
rect 17460 20340 17466 20392
rect 18414 20340 18420 20392
rect 18472 20380 18478 20392
rect 18708 20380 18736 20488
rect 20162 20476 20168 20488
rect 20220 20476 20226 20528
rect 20548 20516 20576 20556
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20680 20556 21097 20584
rect 20680 20544 20686 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 22370 20544 22376 20596
rect 22428 20544 22434 20596
rect 23106 20544 23112 20596
rect 23164 20544 23170 20596
rect 21726 20516 21732 20528
rect 20548 20488 21732 20516
rect 21726 20476 21732 20488
rect 21784 20476 21790 20528
rect 24210 20476 24216 20528
rect 24268 20476 24274 20528
rect 25314 20476 25320 20528
rect 25372 20516 25378 20528
rect 25590 20516 25596 20528
rect 25372 20488 25596 20516
rect 25372 20476 25378 20488
rect 25590 20476 25596 20488
rect 25648 20476 25654 20528
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 19797 20451 19855 20457
rect 19797 20448 19809 20451
rect 19392 20420 19809 20448
rect 19392 20408 19398 20420
rect 19797 20417 19809 20420
rect 19843 20417 19855 20451
rect 19797 20411 19855 20417
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 19935 20420 20116 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 18472 20352 18736 20380
rect 18472 20340 18478 20352
rect 19426 20340 19432 20392
rect 19484 20380 19490 20392
rect 19981 20383 20039 20389
rect 19981 20380 19993 20383
rect 19484 20352 19993 20380
rect 19484 20340 19490 20352
rect 19981 20349 19993 20352
rect 20027 20349 20039 20383
rect 20088 20380 20116 20420
rect 20898 20408 20904 20460
rect 20956 20448 20962 20460
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20956 20420 21005 20448
rect 20956 20408 20962 20420
rect 20993 20417 21005 20420
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 21174 20408 21180 20460
rect 21232 20448 21238 20460
rect 22002 20448 22008 20460
rect 21232 20420 22008 20448
rect 21232 20408 21238 20420
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 23477 20451 23535 20457
rect 23477 20448 23489 20451
rect 23348 20420 23489 20448
rect 23348 20408 23354 20420
rect 23477 20417 23489 20420
rect 23523 20417 23535 20451
rect 23477 20411 23535 20417
rect 21082 20380 21088 20392
rect 20088 20352 21088 20380
rect 19981 20343 20039 20349
rect 21082 20340 21088 20352
rect 21140 20340 21146 20392
rect 21266 20340 21272 20392
rect 21324 20340 21330 20392
rect 21910 20340 21916 20392
rect 21968 20380 21974 20392
rect 22465 20383 22523 20389
rect 21968 20352 22094 20380
rect 21968 20340 21974 20352
rect 17126 20312 17132 20324
rect 12544 20284 13768 20312
rect 13538 20244 13544 20256
rect 12406 20216 13544 20244
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 13740 20244 13768 20284
rect 15304 20284 17132 20312
rect 15304 20244 15332 20284
rect 17126 20272 17132 20284
rect 17184 20272 17190 20324
rect 20162 20272 20168 20324
rect 20220 20312 20226 20324
rect 21284 20312 21312 20340
rect 20220 20284 21312 20312
rect 22066 20312 22094 20352
rect 22465 20349 22477 20383
rect 22511 20349 22523 20383
rect 22465 20343 22523 20349
rect 22480 20312 22508 20343
rect 22646 20340 22652 20392
rect 22704 20340 22710 20392
rect 23750 20340 23756 20392
rect 23808 20340 23814 20392
rect 22066 20284 23612 20312
rect 20220 20272 20226 20284
rect 23584 20256 23612 20284
rect 13740 20216 15332 20244
rect 18506 20204 18512 20256
rect 18564 20244 18570 20256
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18564 20216 18889 20244
rect 18564 20204 18570 20216
rect 18877 20213 18889 20216
rect 18923 20244 18935 20247
rect 18966 20244 18972 20256
rect 18923 20216 18972 20244
rect 18923 20213 18935 20216
rect 18877 20207 18935 20213
rect 18966 20204 18972 20216
rect 19024 20204 19030 20256
rect 19334 20204 19340 20256
rect 19392 20204 19398 20256
rect 19429 20247 19487 20253
rect 19429 20213 19441 20247
rect 19475 20244 19487 20247
rect 19610 20244 19616 20256
rect 19475 20216 19616 20244
rect 19475 20213 19487 20216
rect 19429 20207 19487 20213
rect 19610 20204 19616 20216
rect 19668 20204 19674 20256
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 20625 20247 20683 20253
rect 20625 20244 20637 20247
rect 20128 20216 20637 20244
rect 20128 20204 20134 20216
rect 20625 20213 20637 20216
rect 20671 20213 20683 20247
rect 20625 20207 20683 20213
rect 21266 20204 21272 20256
rect 21324 20244 21330 20256
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 21324 20216 22017 20244
rect 21324 20204 21330 20216
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 22005 20207 22063 20213
rect 23566 20204 23572 20256
rect 23624 20204 23630 20256
rect 25130 20204 25136 20256
rect 25188 20244 25194 20256
rect 25225 20247 25283 20253
rect 25225 20244 25237 20247
rect 25188 20216 25237 20244
rect 25188 20204 25194 20216
rect 25225 20213 25237 20216
rect 25271 20213 25283 20247
rect 25225 20207 25283 20213
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 3878 20000 3884 20052
rect 3936 20040 3942 20052
rect 3973 20043 4031 20049
rect 3973 20040 3985 20043
rect 3936 20012 3985 20040
rect 3936 20000 3942 20012
rect 3973 20009 3985 20012
rect 4019 20009 4031 20043
rect 7466 20040 7472 20052
rect 3973 20003 4031 20009
rect 4080 20012 7472 20040
rect 2774 19864 2780 19916
rect 2832 19864 2838 19916
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19836 2283 19839
rect 4080 19836 4108 20012
rect 7466 20000 7472 20012
rect 7524 20000 7530 20052
rect 7650 20000 7656 20052
rect 7708 20040 7714 20052
rect 9398 20040 9404 20052
rect 7708 20012 9404 20040
rect 7708 20000 7714 20012
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 9508 20012 9720 20040
rect 4154 19932 4160 19984
rect 4212 19972 4218 19984
rect 4338 19972 4344 19984
rect 4212 19944 4344 19972
rect 4212 19932 4218 19944
rect 4338 19932 4344 19944
rect 4396 19932 4402 19984
rect 9508 19972 9536 20012
rect 4632 19944 9536 19972
rect 9692 19972 9720 20012
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 16117 20043 16175 20049
rect 16117 20040 16129 20043
rect 10008 20012 16129 20040
rect 10008 20000 10014 20012
rect 16117 20009 16129 20012
rect 16163 20009 16175 20043
rect 16117 20003 16175 20009
rect 17126 20000 17132 20052
rect 17184 20040 17190 20052
rect 17773 20043 17831 20049
rect 17773 20040 17785 20043
rect 17184 20012 17785 20040
rect 17184 20000 17190 20012
rect 17773 20009 17785 20012
rect 17819 20009 17831 20043
rect 17773 20003 17831 20009
rect 21818 20000 21824 20052
rect 21876 20040 21882 20052
rect 21876 20012 22232 20040
rect 21876 20000 21882 20012
rect 13265 19975 13323 19981
rect 9692 19944 11652 19972
rect 2271 19808 4108 19836
rect 4157 19839 4215 19845
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4522 19836 4528 19848
rect 4203 19808 4528 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 4632 19845 4660 19944
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 8662 19904 8668 19916
rect 5684 19876 8668 19904
rect 5684 19864 5690 19876
rect 8662 19864 8668 19876
rect 8720 19864 8726 19916
rect 9677 19907 9735 19913
rect 9677 19873 9689 19907
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19836 5779 19839
rect 6730 19836 6736 19848
rect 5767 19808 6736 19836
rect 5767 19805 5779 19808
rect 5721 19799 5779 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 6822 19796 6828 19848
rect 6880 19796 6886 19848
rect 7469 19839 7527 19845
rect 7469 19805 7481 19839
rect 7515 19836 7527 19839
rect 7929 19839 7987 19845
rect 7929 19836 7941 19839
rect 7515 19808 7941 19836
rect 7515 19805 7527 19808
rect 7469 19799 7527 19805
rect 7929 19805 7941 19808
rect 7975 19805 7987 19839
rect 9692 19836 9720 19867
rect 10870 19864 10876 19916
rect 10928 19864 10934 19916
rect 11624 19904 11652 19944
rect 13265 19941 13277 19975
rect 13311 19972 13323 19975
rect 13446 19972 13452 19984
rect 13311 19944 13452 19972
rect 13311 19941 13323 19944
rect 13265 19935 13323 19941
rect 13280 19904 13308 19935
rect 13446 19932 13452 19944
rect 13504 19932 13510 19984
rect 13722 19932 13728 19984
rect 13780 19932 13786 19984
rect 13906 19932 13912 19984
rect 13964 19972 13970 19984
rect 15102 19972 15108 19984
rect 13964 19944 15108 19972
rect 13964 19932 13970 19944
rect 15102 19932 15108 19944
rect 15160 19932 15166 19984
rect 19429 19975 19487 19981
rect 19429 19972 19441 19975
rect 15304 19944 19441 19972
rect 15010 19904 15016 19916
rect 11624 19876 13308 19904
rect 14200 19876 15016 19904
rect 10686 19836 10692 19848
rect 7929 19799 7987 19805
rect 8496 19808 10692 19836
rect 1765 19771 1823 19777
rect 1765 19737 1777 19771
rect 1811 19768 1823 19771
rect 1811 19740 2774 19768
rect 1811 19737 1823 19740
rect 1765 19731 1823 19737
rect 2746 19700 2774 19740
rect 3970 19728 3976 19780
rect 4028 19768 4034 19780
rect 8496 19768 8524 19808
rect 10686 19796 10692 19808
rect 10744 19796 10750 19848
rect 11514 19796 11520 19848
rect 11572 19796 11578 19848
rect 13354 19796 13360 19848
rect 13412 19836 13418 19848
rect 14200 19836 14228 19876
rect 15010 19864 15016 19876
rect 15068 19864 15074 19916
rect 14734 19836 14740 19848
rect 13412 19808 14228 19836
rect 14292 19808 14740 19836
rect 13412 19796 13418 19808
rect 4028 19740 8524 19768
rect 8573 19771 8631 19777
rect 4028 19728 4034 19740
rect 8573 19737 8585 19771
rect 8619 19768 8631 19771
rect 11793 19771 11851 19777
rect 11793 19768 11805 19771
rect 8619 19740 11805 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 11793 19737 11805 19740
rect 11839 19737 11851 19771
rect 13814 19768 13820 19780
rect 13018 19740 13820 19768
rect 11793 19731 11851 19737
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 14292 19768 14320 19808
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 15304 19845 15332 19944
rect 19429 19941 19441 19944
rect 19475 19941 19487 19975
rect 22204 19972 22232 20012
rect 22278 20000 22284 20052
rect 22336 20040 22342 20052
rect 23198 20040 23204 20052
rect 22336 20012 23204 20040
rect 22336 20000 22342 20012
rect 23198 20000 23204 20012
rect 23256 20000 23262 20052
rect 22370 19972 22376 19984
rect 22204 19944 22376 19972
rect 19429 19935 19487 19941
rect 22370 19932 22376 19944
rect 22428 19932 22434 19984
rect 23106 19932 23112 19984
rect 23164 19972 23170 19984
rect 23474 19972 23480 19984
rect 23164 19944 23480 19972
rect 23164 19932 23170 19944
rect 23474 19932 23480 19944
rect 23532 19972 23538 19984
rect 23532 19944 23704 19972
rect 23532 19932 23538 19944
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19805 15347 19839
rect 15488 19836 15516 19867
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 15620 19876 16681 19904
rect 15620 19864 15626 19876
rect 16669 19873 16681 19876
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 17126 19904 17132 19916
rect 16816 19876 17132 19904
rect 16816 19864 16822 19876
rect 17126 19864 17132 19876
rect 17184 19904 17190 19916
rect 17405 19907 17463 19913
rect 17405 19904 17417 19907
rect 17184 19876 17417 19904
rect 17184 19864 17190 19876
rect 17405 19873 17417 19876
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 18322 19864 18328 19916
rect 18380 19864 18386 19916
rect 19058 19864 19064 19916
rect 19116 19904 19122 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19116 19876 19993 19904
rect 19116 19864 19122 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19904 20959 19907
rect 23290 19904 23296 19916
rect 20947 19876 23296 19904
rect 20947 19873 20959 19876
rect 20901 19867 20959 19873
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 23676 19913 23704 19944
rect 23661 19907 23719 19913
rect 23661 19873 23673 19907
rect 23707 19873 23719 19907
rect 23661 19867 23719 19873
rect 24394 19864 24400 19916
rect 24452 19904 24458 19916
rect 25133 19907 25191 19913
rect 25133 19904 25145 19907
rect 24452 19876 25145 19904
rect 24452 19864 24458 19876
rect 25133 19873 25145 19876
rect 25179 19873 25191 19907
rect 25133 19867 25191 19873
rect 16022 19836 16028 19848
rect 15488 19808 16028 19836
rect 15289 19799 15347 19805
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 16482 19796 16488 19848
rect 16540 19836 16546 19848
rect 16577 19839 16635 19845
rect 16577 19836 16589 19839
rect 16540 19808 16589 19836
rect 16540 19796 16546 19808
rect 16577 19805 16589 19808
rect 16623 19805 16635 19839
rect 16577 19799 16635 19805
rect 17218 19796 17224 19848
rect 17276 19836 17282 19848
rect 17313 19839 17371 19845
rect 17313 19836 17325 19839
rect 17276 19808 17325 19836
rect 17276 19796 17282 19808
rect 17313 19805 17325 19808
rect 17359 19836 17371 19839
rect 17586 19836 17592 19848
rect 17359 19808 17592 19836
rect 17359 19805 17371 19808
rect 17313 19799 17371 19805
rect 17586 19796 17592 19808
rect 17644 19836 17650 19848
rect 18233 19839 18291 19845
rect 18233 19836 18245 19839
rect 17644 19808 18245 19836
rect 17644 19796 17650 19808
rect 18233 19805 18245 19808
rect 18279 19805 18291 19839
rect 18233 19799 18291 19805
rect 18874 19796 18880 19848
rect 18932 19836 18938 19848
rect 20530 19836 20536 19848
rect 18932 19808 20536 19836
rect 18932 19796 18938 19808
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 22462 19796 22468 19848
rect 22520 19836 22526 19848
rect 22922 19836 22928 19848
rect 22520 19808 22928 19836
rect 22520 19796 22526 19808
rect 22922 19796 22928 19808
rect 22980 19836 22986 19848
rect 24121 19839 24179 19845
rect 24121 19836 24133 19839
rect 22980 19808 24133 19836
rect 22980 19796 22986 19808
rect 24121 19805 24133 19808
rect 24167 19805 24179 19839
rect 24121 19799 24179 19805
rect 13924 19740 14320 19768
rect 4522 19700 4528 19712
rect 2746 19672 4528 19700
rect 4522 19660 4528 19672
rect 4580 19660 4586 19712
rect 5261 19703 5319 19709
rect 5261 19669 5273 19703
rect 5307 19700 5319 19703
rect 5350 19700 5356 19712
rect 5307 19672 5356 19700
rect 5307 19669 5319 19672
rect 5261 19663 5319 19669
rect 5350 19660 5356 19672
rect 5408 19660 5414 19712
rect 5718 19660 5724 19712
rect 5776 19700 5782 19712
rect 6365 19703 6423 19709
rect 6365 19700 6377 19703
rect 5776 19672 6377 19700
rect 5776 19660 5782 19672
rect 6365 19669 6377 19672
rect 6411 19669 6423 19703
rect 6365 19663 6423 19669
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 9125 19703 9183 19709
rect 9125 19700 9137 19703
rect 8444 19672 9137 19700
rect 8444 19660 8450 19672
rect 9125 19669 9137 19672
rect 9171 19669 9183 19703
rect 9125 19663 9183 19669
rect 9214 19660 9220 19712
rect 9272 19700 9278 19712
rect 9493 19703 9551 19709
rect 9493 19700 9505 19703
rect 9272 19672 9505 19700
rect 9272 19660 9278 19672
rect 9493 19669 9505 19672
rect 9539 19669 9551 19703
rect 9493 19663 9551 19669
rect 9585 19703 9643 19709
rect 9585 19669 9597 19703
rect 9631 19700 9643 19703
rect 9950 19700 9956 19712
rect 9631 19672 9956 19700
rect 9631 19669 9643 19672
rect 9585 19663 9643 19669
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 10318 19660 10324 19712
rect 10376 19660 10382 19712
rect 10410 19660 10416 19712
rect 10468 19700 10474 19712
rect 10689 19703 10747 19709
rect 10689 19700 10701 19703
rect 10468 19672 10701 19700
rect 10468 19660 10474 19672
rect 10689 19669 10701 19672
rect 10735 19669 10747 19703
rect 10689 19663 10747 19669
rect 10781 19703 10839 19709
rect 10781 19669 10793 19703
rect 10827 19700 10839 19703
rect 13924 19700 13952 19740
rect 14366 19728 14372 19780
rect 14424 19768 14430 19780
rect 15381 19771 15439 19777
rect 15381 19768 15393 19771
rect 14424 19740 15393 19768
rect 14424 19728 14430 19740
rect 15381 19737 15393 19740
rect 15427 19737 15439 19771
rect 18506 19768 18512 19780
rect 15381 19731 15439 19737
rect 16408 19740 18512 19768
rect 10827 19672 13952 19700
rect 10827 19669 10839 19672
rect 10781 19663 10839 19669
rect 13998 19660 14004 19712
rect 14056 19700 14062 19712
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 14056 19672 14289 19700
rect 14056 19660 14062 19672
rect 14277 19669 14289 19672
rect 14323 19669 14335 19703
rect 14277 19663 14335 19669
rect 14918 19660 14924 19712
rect 14976 19660 14982 19712
rect 15010 19660 15016 19712
rect 15068 19700 15074 19712
rect 16408 19700 16436 19740
rect 18506 19728 18512 19740
rect 18564 19728 18570 19780
rect 19889 19771 19947 19777
rect 19889 19768 19901 19771
rect 18800 19740 19901 19768
rect 15068 19672 16436 19700
rect 15068 19660 15074 19672
rect 16482 19660 16488 19712
rect 16540 19660 16546 19712
rect 17586 19660 17592 19712
rect 17644 19700 17650 19712
rect 18141 19703 18199 19709
rect 18141 19700 18153 19703
rect 17644 19672 18153 19700
rect 17644 19660 17650 19672
rect 18141 19669 18153 19672
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 18690 19660 18696 19712
rect 18748 19700 18754 19712
rect 18800 19709 18828 19740
rect 19889 19737 19901 19740
rect 19935 19737 19947 19771
rect 19889 19731 19947 19737
rect 20809 19771 20867 19777
rect 20809 19737 20821 19771
rect 20855 19768 20867 19771
rect 21174 19768 21180 19780
rect 20855 19740 21180 19768
rect 20855 19737 20867 19740
rect 20809 19731 20867 19737
rect 21174 19728 21180 19740
rect 21232 19728 21238 19780
rect 25041 19771 25099 19777
rect 25041 19768 25053 19771
rect 21560 19740 21666 19768
rect 23124 19740 25053 19768
rect 18785 19703 18843 19709
rect 18785 19700 18797 19703
rect 18748 19672 18797 19700
rect 18748 19660 18754 19672
rect 18785 19669 18797 19672
rect 18831 19669 18843 19703
rect 18785 19663 18843 19669
rect 18966 19660 18972 19712
rect 19024 19660 19030 19712
rect 19337 19703 19395 19709
rect 19337 19669 19349 19703
rect 19383 19700 19395 19703
rect 19518 19700 19524 19712
rect 19383 19672 19524 19700
rect 19383 19669 19395 19672
rect 19337 19663 19395 19669
rect 19518 19660 19524 19672
rect 19576 19700 19582 19712
rect 19797 19703 19855 19709
rect 19797 19700 19809 19703
rect 19576 19672 19809 19700
rect 19576 19660 19582 19672
rect 19797 19669 19809 19672
rect 19843 19700 19855 19703
rect 20257 19703 20315 19709
rect 20257 19700 20269 19703
rect 19843 19672 20269 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 20257 19669 20269 19672
rect 20303 19669 20315 19703
rect 20257 19663 20315 19669
rect 20438 19660 20444 19712
rect 20496 19660 20502 19712
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 21450 19700 21456 19712
rect 20772 19672 21456 19700
rect 20772 19660 20778 19672
rect 21450 19660 21456 19672
rect 21508 19700 21514 19712
rect 21560 19700 21588 19740
rect 21508 19672 21588 19700
rect 22649 19703 22707 19709
rect 21508 19660 21514 19672
rect 22649 19669 22661 19703
rect 22695 19700 22707 19703
rect 23014 19700 23020 19712
rect 22695 19672 23020 19700
rect 22695 19669 22707 19672
rect 22649 19663 22707 19669
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 23124 19709 23152 19740
rect 25041 19737 25053 19740
rect 25087 19737 25099 19771
rect 25041 19731 25099 19737
rect 23109 19703 23167 19709
rect 23109 19669 23121 19703
rect 23155 19669 23167 19703
rect 23109 19663 23167 19669
rect 23198 19660 23204 19712
rect 23256 19700 23262 19712
rect 23477 19703 23535 19709
rect 23477 19700 23489 19703
rect 23256 19672 23489 19700
rect 23256 19660 23262 19672
rect 23477 19669 23489 19672
rect 23523 19669 23535 19703
rect 23477 19663 23535 19669
rect 23569 19703 23627 19709
rect 23569 19669 23581 19703
rect 23615 19700 23627 19703
rect 23750 19700 23756 19712
rect 23615 19672 23756 19700
rect 23615 19669 23627 19672
rect 23569 19663 23627 19669
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 24578 19660 24584 19712
rect 24636 19660 24642 19712
rect 24949 19703 25007 19709
rect 24949 19669 24961 19703
rect 24995 19700 25007 19703
rect 25314 19700 25320 19712
rect 24995 19672 25320 19700
rect 24995 19669 25007 19672
rect 24949 19663 25007 19669
rect 25314 19660 25320 19672
rect 25372 19660 25378 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 3605 19499 3663 19505
rect 3605 19465 3617 19499
rect 3651 19496 3663 19499
rect 4062 19496 4068 19508
rect 3651 19468 4068 19496
rect 3651 19465 3663 19468
rect 3605 19459 3663 19465
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 5626 19496 5632 19508
rect 4172 19468 5632 19496
rect 1486 19388 1492 19440
rect 1544 19428 1550 19440
rect 4172 19428 4200 19468
rect 5626 19456 5632 19468
rect 5684 19456 5690 19508
rect 5994 19456 6000 19508
rect 6052 19456 6058 19508
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 7377 19499 7435 19505
rect 7377 19496 7389 19499
rect 6788 19468 7389 19496
rect 6788 19456 6794 19468
rect 7377 19465 7389 19468
rect 7423 19465 7435 19499
rect 7377 19459 7435 19465
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 7524 19468 10548 19496
rect 7524 19456 7530 19468
rect 6270 19428 6276 19440
rect 1544 19400 4200 19428
rect 4264 19400 6276 19428
rect 1544 19388 1550 19400
rect 1946 19320 1952 19372
rect 2004 19320 2010 19372
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19360 3847 19363
rect 4154 19360 4160 19372
rect 3835 19332 4160 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 4264 19369 4292 19400
rect 6270 19388 6276 19400
rect 6328 19388 6334 19440
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 8481 19431 8539 19437
rect 8481 19428 8493 19431
rect 6972 19400 8493 19428
rect 6972 19388 6978 19400
rect 8481 19397 8493 19400
rect 8527 19397 8539 19431
rect 10520 19428 10548 19468
rect 10686 19456 10692 19508
rect 10744 19456 10750 19508
rect 11514 19456 11520 19508
rect 11572 19496 11578 19508
rect 14274 19496 14280 19508
rect 11572 19468 14280 19496
rect 11572 19456 11578 19468
rect 12069 19431 12127 19437
rect 12069 19428 12081 19431
rect 10520 19400 12081 19428
rect 8481 19391 8539 19397
rect 12069 19397 12081 19400
rect 12115 19397 12127 19431
rect 12069 19391 12127 19397
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 5350 19320 5356 19372
rect 5408 19320 5414 19372
rect 6638 19320 6644 19372
rect 6696 19360 6702 19372
rect 6733 19363 6791 19369
rect 6733 19360 6745 19363
rect 6696 19332 6745 19360
rect 6696 19320 6702 19332
rect 6733 19329 6745 19332
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 7650 19360 7656 19372
rect 7524 19332 7656 19360
rect 7524 19320 7530 19332
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 7834 19320 7840 19372
rect 7892 19320 7898 19372
rect 8938 19320 8944 19372
rect 8996 19320 9002 19372
rect 10318 19320 10324 19372
rect 10376 19320 10382 19372
rect 11333 19363 11391 19369
rect 11333 19329 11345 19363
rect 11379 19360 11391 19363
rect 11882 19360 11888 19372
rect 11379 19332 11888 19360
rect 11379 19329 11391 19332
rect 11333 19323 11391 19329
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 12544 19369 12572 19468
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 14734 19456 14740 19508
rect 14792 19456 14798 19508
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 15102 19496 15108 19508
rect 14884 19468 15108 19496
rect 14884 19456 14890 19468
rect 15102 19456 15108 19468
rect 15160 19496 15166 19508
rect 15197 19499 15255 19505
rect 15197 19496 15209 19499
rect 15160 19468 15209 19496
rect 15160 19456 15166 19468
rect 15197 19465 15209 19468
rect 15243 19465 15255 19499
rect 15197 19459 15255 19465
rect 17678 19456 17684 19508
rect 17736 19496 17742 19508
rect 17736 19468 18736 19496
rect 17736 19456 17742 19468
rect 12802 19388 12808 19440
rect 12860 19388 12866 19440
rect 16942 19428 16948 19440
rect 15028 19400 16948 19428
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19329 12587 19363
rect 12529 19323 12587 19329
rect 13906 19320 13912 19372
rect 13964 19320 13970 19372
rect 15028 19360 15056 19400
rect 16942 19388 16948 19400
rect 17000 19388 17006 19440
rect 18708 19428 18736 19468
rect 19610 19456 19616 19508
rect 19668 19456 19674 19508
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 20990 19496 20996 19508
rect 20947 19468 20996 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21358 19456 21364 19508
rect 21416 19496 21422 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21416 19468 22017 19496
rect 21416 19456 21422 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22373 19499 22431 19505
rect 22373 19465 22385 19499
rect 22419 19496 22431 19499
rect 22554 19496 22560 19508
rect 22419 19468 22560 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 22554 19456 22560 19468
rect 22612 19456 22618 19508
rect 25041 19499 25099 19505
rect 25041 19465 25053 19499
rect 25087 19496 25099 19499
rect 25222 19496 25228 19508
rect 25087 19468 25228 19496
rect 25087 19465 25099 19468
rect 25041 19459 25099 19465
rect 25222 19456 25228 19468
rect 25280 19496 25286 19508
rect 26510 19496 26516 19508
rect 25280 19468 26516 19496
rect 25280 19456 25286 19468
rect 26510 19456 26516 19468
rect 26568 19456 26574 19508
rect 19705 19431 19763 19437
rect 19705 19428 19717 19431
rect 18708 19400 19717 19428
rect 19705 19397 19717 19400
rect 19751 19397 19763 19431
rect 19705 19391 19763 19397
rect 21450 19388 21456 19440
rect 21508 19428 21514 19440
rect 21508 19400 24058 19428
rect 21508 19388 21514 19400
rect 14016 19332 15056 19360
rect 1578 19252 1584 19304
rect 1636 19292 1642 19304
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 1636 19264 2237 19292
rect 1636 19252 1642 19264
rect 2225 19261 2237 19264
rect 2271 19261 2283 19295
rect 2225 19255 2283 19261
rect 2590 19252 2596 19304
rect 2648 19292 2654 19304
rect 4522 19292 4528 19304
rect 2648 19264 4528 19292
rect 2648 19252 2654 19264
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 4893 19295 4951 19301
rect 4893 19261 4905 19295
rect 4939 19292 4951 19295
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 4939 19264 9229 19292
rect 4939 19261 4951 19264
rect 4893 19255 4951 19261
rect 9217 19261 9229 19264
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 11112 19264 11161 19292
rect 11112 19252 11118 19264
rect 11149 19261 11161 19264
rect 11195 19292 11207 19295
rect 12250 19292 12256 19304
rect 11195 19264 12256 19292
rect 11195 19261 11207 19264
rect 11149 19255 11207 19261
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 13354 19292 13360 19304
rect 12544 19264 13360 19292
rect 4154 19184 4160 19236
rect 4212 19224 4218 19236
rect 5258 19224 5264 19236
rect 4212 19196 5264 19224
rect 4212 19184 4218 19196
rect 5258 19184 5264 19196
rect 5316 19224 5322 19236
rect 6365 19227 6423 19233
rect 6365 19224 6377 19227
rect 5316 19196 6377 19224
rect 5316 19184 5322 19196
rect 6365 19193 6377 19196
rect 6411 19193 6423 19227
rect 6365 19187 6423 19193
rect 7006 19184 7012 19236
rect 7064 19224 7070 19236
rect 8754 19224 8760 19236
rect 7064 19196 8760 19224
rect 7064 19184 7070 19196
rect 8754 19184 8760 19196
rect 8812 19184 8818 19236
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 12544 19156 12572 19264
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13446 19252 13452 19304
rect 13504 19292 13510 19304
rect 14016 19292 14044 19332
rect 15102 19320 15108 19372
rect 15160 19320 15166 19372
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 15436 19332 16129 19360
rect 15436 19320 15442 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 17034 19320 17040 19372
rect 17092 19320 17098 19372
rect 20714 19360 20720 19372
rect 18446 19332 20720 19360
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 21082 19360 21088 19372
rect 20855 19332 21088 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21634 19320 21640 19372
rect 21692 19360 21698 19372
rect 22278 19360 22284 19372
rect 21692 19332 22284 19360
rect 21692 19320 21698 19332
rect 22278 19320 22284 19332
rect 22336 19320 22342 19372
rect 22465 19363 22523 19369
rect 22465 19329 22477 19363
rect 22511 19329 22523 19363
rect 23106 19360 23112 19372
rect 22465 19323 22523 19329
rect 22572 19332 23112 19360
rect 13504 19264 14044 19292
rect 13504 19252 13510 19264
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 15289 19295 15347 19301
rect 15289 19292 15301 19295
rect 14148 19264 15301 19292
rect 14148 19252 14154 19264
rect 15289 19261 15301 19264
rect 15335 19261 15347 19295
rect 17313 19295 17371 19301
rect 17313 19292 17325 19295
rect 15289 19255 15347 19261
rect 15396 19264 17325 19292
rect 15396 19224 15424 19264
rect 17313 19261 17325 19264
rect 17359 19261 17371 19295
rect 19797 19295 19855 19301
rect 19797 19292 19809 19295
rect 17313 19255 17371 19261
rect 18800 19264 19809 19292
rect 13832 19196 15424 19224
rect 16132 19196 17080 19224
rect 7340 19128 12572 19156
rect 7340 19116 7346 19128
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 13832 19156 13860 19196
rect 13412 19128 13860 19156
rect 14277 19159 14335 19165
rect 13412 19116 13418 19128
rect 14277 19125 14289 19159
rect 14323 19156 14335 19159
rect 14458 19156 14464 19168
rect 14323 19128 14464 19156
rect 14323 19125 14335 19128
rect 14277 19119 14335 19125
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 15010 19116 15016 19168
rect 15068 19156 15074 19168
rect 16132 19156 16160 19196
rect 15068 19128 16160 19156
rect 15068 19116 15074 19128
rect 16206 19116 16212 19168
rect 16264 19116 16270 19168
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 16666 19156 16672 19168
rect 16448 19128 16672 19156
rect 16448 19116 16454 19128
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 16758 19116 16764 19168
rect 16816 19116 16822 19168
rect 17052 19156 17080 19196
rect 18800 19165 18828 19264
rect 19797 19261 19809 19264
rect 19843 19261 19855 19295
rect 19797 19255 19855 19261
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20956 19264 21005 19292
rect 20956 19252 20962 19264
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 19978 19184 19984 19236
rect 20036 19224 20042 19236
rect 22480 19224 22508 19323
rect 22572 19304 22600 19332
rect 23106 19320 23112 19332
rect 23164 19320 23170 19372
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 22554 19252 22560 19304
rect 22612 19252 22618 19304
rect 22646 19252 22652 19304
rect 22704 19252 22710 19304
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 23934 19292 23940 19304
rect 23615 19264 23940 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 23934 19252 23940 19264
rect 23992 19252 23998 19304
rect 24762 19252 24768 19304
rect 24820 19292 24826 19304
rect 25222 19292 25228 19304
rect 24820 19264 25228 19292
rect 24820 19252 24826 19264
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 22922 19224 22928 19236
rect 20036 19196 22094 19224
rect 22480 19196 22928 19224
rect 20036 19184 20042 19196
rect 18785 19159 18843 19165
rect 18785 19156 18797 19159
rect 17052 19128 18797 19156
rect 18785 19125 18797 19128
rect 18831 19125 18843 19159
rect 18785 19119 18843 19125
rect 19242 19116 19248 19168
rect 19300 19116 19306 19168
rect 20438 19116 20444 19168
rect 20496 19116 20502 19168
rect 20806 19116 20812 19168
rect 20864 19156 20870 19168
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 20864 19128 21465 19156
rect 20864 19116 20870 19128
rect 21453 19125 21465 19128
rect 21499 19156 21511 19159
rect 21634 19156 21640 19168
rect 21499 19128 21640 19156
rect 21499 19125 21511 19128
rect 21453 19119 21511 19125
rect 21634 19116 21640 19128
rect 21692 19116 21698 19168
rect 22066 19156 22094 19196
rect 22922 19184 22928 19196
rect 22980 19184 22986 19236
rect 25409 19227 25467 19233
rect 25409 19224 25421 19227
rect 24596 19196 25421 19224
rect 24596 19156 24624 19196
rect 25409 19193 25421 19196
rect 25455 19193 25467 19227
rect 25409 19187 25467 19193
rect 22066 19128 24624 19156
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 4798 18912 4804 18964
rect 4856 18952 4862 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 4856 18924 9229 18952
rect 4856 18912 4862 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 9217 18915 9275 18921
rect 9490 18912 9496 18964
rect 9548 18952 9554 18964
rect 12342 18952 12348 18964
rect 9548 18924 12348 18952
rect 9548 18912 9554 18924
rect 12342 18912 12348 18924
rect 12400 18952 12406 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 12400 18924 12449 18952
rect 12400 18912 12406 18924
rect 12437 18921 12449 18924
rect 12483 18921 12495 18955
rect 14277 18955 14335 18961
rect 12437 18915 12495 18921
rect 12544 18924 13860 18952
rect 12066 18884 12072 18896
rect 7944 18856 12072 18884
rect 1670 18708 1676 18760
rect 1728 18708 1734 18760
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18748 2835 18751
rect 3970 18748 3976 18760
rect 2823 18720 3976 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 4614 18708 4620 18760
rect 4672 18708 4678 18760
rect 5718 18708 5724 18760
rect 5776 18708 5782 18760
rect 6362 18708 6368 18760
rect 6420 18748 6426 18760
rect 6638 18748 6644 18760
rect 6420 18720 6644 18748
rect 6420 18708 6426 18720
rect 6638 18708 6644 18720
rect 6696 18708 6702 18760
rect 6822 18708 6828 18760
rect 6880 18708 6886 18760
rect 7944 18757 7972 18856
rect 12066 18844 12072 18856
rect 12124 18844 12130 18896
rect 12250 18844 12256 18896
rect 12308 18884 12314 18896
rect 12544 18884 12572 18924
rect 12308 18856 12572 18884
rect 12308 18844 12314 18856
rect 12986 18844 12992 18896
rect 13044 18844 13050 18896
rect 13170 18844 13176 18896
rect 13228 18884 13234 18896
rect 13722 18884 13728 18896
rect 13228 18856 13728 18884
rect 13228 18844 13234 18856
rect 13722 18844 13728 18856
rect 13780 18844 13786 18896
rect 13832 18884 13860 18924
rect 14277 18921 14289 18955
rect 14323 18952 14335 18955
rect 14366 18952 14372 18964
rect 14323 18924 14372 18952
rect 14323 18921 14335 18924
rect 14277 18915 14335 18921
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 19058 18952 19064 18964
rect 15672 18924 19064 18952
rect 15562 18884 15568 18896
rect 13832 18856 15568 18884
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 9306 18776 9312 18828
rect 9364 18816 9370 18828
rect 9769 18819 9827 18825
rect 9769 18816 9781 18819
rect 9364 18788 9781 18816
rect 9364 18776 9370 18788
rect 9769 18785 9781 18788
rect 9815 18785 9827 18819
rect 9769 18779 9827 18785
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 12618 18816 12624 18828
rect 11020 18788 12624 18816
rect 11020 18776 11026 18788
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 13188 18788 13400 18816
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 10134 18708 10140 18760
rect 10192 18748 10198 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 10192 18720 10425 18748
rect 10192 18708 10198 18720
rect 10413 18717 10425 18720
rect 10459 18748 10471 18751
rect 12250 18748 12256 18760
rect 10459 18720 12256 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 12713 18751 12771 18757
rect 12713 18717 12725 18751
rect 12759 18748 12771 18751
rect 13078 18748 13084 18760
rect 12759 18720 13084 18748
rect 12759 18717 12771 18720
rect 12713 18711 12771 18717
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 5626 18680 5632 18692
rect 3988 18652 5632 18680
rect 2222 18572 2228 18624
rect 2280 18612 2286 18624
rect 2317 18615 2375 18621
rect 2317 18612 2329 18615
rect 2280 18584 2329 18612
rect 2280 18572 2286 18584
rect 2317 18581 2329 18584
rect 2363 18581 2375 18615
rect 2317 18575 2375 18581
rect 3418 18572 3424 18624
rect 3476 18572 3482 18624
rect 3988 18621 4016 18652
rect 5626 18640 5632 18652
rect 5684 18640 5690 18692
rect 5994 18640 6000 18692
rect 6052 18680 6058 18692
rect 9490 18680 9496 18692
rect 6052 18652 9496 18680
rect 6052 18640 6058 18652
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 9585 18683 9643 18689
rect 9585 18649 9597 18683
rect 9631 18680 9643 18683
rect 13188 18680 13216 18788
rect 13372 18748 13400 18788
rect 13446 18776 13452 18828
rect 13504 18776 13510 18828
rect 13630 18776 13636 18828
rect 13688 18776 13694 18828
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 14921 18819 14979 18825
rect 14921 18816 14933 18819
rect 13872 18788 14933 18816
rect 13872 18776 13878 18788
rect 14921 18785 14933 18788
rect 14967 18816 14979 18819
rect 15672 18816 15700 18924
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 23658 18952 23664 18964
rect 19944 18924 23664 18952
rect 19944 18912 19950 18924
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 17313 18887 17371 18893
rect 17313 18853 17325 18887
rect 17359 18884 17371 18887
rect 17586 18884 17592 18896
rect 17359 18856 17592 18884
rect 17359 18853 17371 18856
rect 17313 18847 17371 18853
rect 17586 18844 17592 18856
rect 17644 18844 17650 18896
rect 18049 18887 18107 18893
rect 18049 18853 18061 18887
rect 18095 18884 18107 18887
rect 19334 18884 19340 18896
rect 18095 18856 19340 18884
rect 18095 18853 18107 18856
rect 18049 18847 18107 18853
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 21634 18844 21640 18896
rect 21692 18884 21698 18896
rect 21910 18884 21916 18896
rect 21692 18856 21916 18884
rect 21692 18844 21698 18856
rect 21910 18844 21916 18856
rect 21968 18844 21974 18896
rect 22646 18844 22652 18896
rect 22704 18884 22710 18896
rect 23382 18884 23388 18896
rect 22704 18856 23388 18884
rect 22704 18844 22710 18856
rect 23382 18844 23388 18856
rect 23440 18844 23446 18896
rect 23937 18887 23995 18893
rect 23937 18853 23949 18887
rect 23983 18884 23995 18887
rect 26602 18884 26608 18896
rect 23983 18856 26608 18884
rect 23983 18853 23995 18856
rect 23937 18847 23995 18853
rect 26602 18844 26608 18856
rect 26660 18844 26666 18896
rect 14967 18788 15700 18816
rect 15841 18819 15899 18825
rect 14967 18785 14979 18788
rect 14921 18779 14979 18785
rect 15841 18785 15853 18819
rect 15887 18816 15899 18819
rect 16298 18816 16304 18828
rect 15887 18788 16304 18816
rect 15887 18785 15899 18788
rect 15841 18779 15899 18785
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 16908 18788 17448 18816
rect 16908 18776 16914 18788
rect 13998 18748 14004 18760
rect 13372 18720 14004 18748
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 14274 18708 14280 18760
rect 14332 18748 14338 18760
rect 15565 18751 15623 18757
rect 15565 18748 15577 18751
rect 14332 18720 15577 18748
rect 14332 18708 14338 18720
rect 15565 18717 15577 18720
rect 15611 18717 15623 18751
rect 17420 18748 17448 18788
rect 17494 18776 17500 18828
rect 17552 18816 17558 18828
rect 18601 18819 18659 18825
rect 18601 18816 18613 18819
rect 17552 18788 18613 18816
rect 17552 18776 17558 18788
rect 18601 18785 18613 18788
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 20254 18776 20260 18828
rect 20312 18776 20318 18828
rect 20530 18776 20536 18828
rect 20588 18776 20594 18828
rect 20622 18776 20628 18828
rect 20680 18816 20686 18828
rect 23109 18819 23167 18825
rect 20680 18788 21772 18816
rect 20680 18776 20686 18788
rect 18782 18748 18788 18760
rect 17420 18720 18788 18748
rect 15565 18711 15623 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 21744 18748 21772 18788
rect 23109 18785 23121 18819
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 22738 18748 22744 18760
rect 9631 18652 13216 18680
rect 9631 18649 9643 18652
rect 9585 18643 9643 18649
rect 13354 18640 13360 18692
rect 13412 18640 13418 18692
rect 14737 18683 14795 18689
rect 14737 18649 14749 18683
rect 14783 18680 14795 18683
rect 14826 18680 14832 18692
rect 14783 18652 14832 18680
rect 14783 18649 14795 18652
rect 14737 18643 14795 18649
rect 14826 18640 14832 18652
rect 14884 18640 14890 18692
rect 16574 18640 16580 18692
rect 16632 18640 16638 18692
rect 19150 18680 19156 18692
rect 17144 18652 19156 18680
rect 3973 18615 4031 18621
rect 3973 18581 3985 18615
rect 4019 18581 4031 18615
rect 3973 18575 4031 18581
rect 5258 18572 5264 18624
rect 5316 18572 5322 18624
rect 5810 18572 5816 18624
rect 5868 18612 5874 18624
rect 6178 18612 6184 18624
rect 5868 18584 6184 18612
rect 5868 18572 5874 18584
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 6362 18572 6368 18624
rect 6420 18572 6426 18624
rect 7006 18572 7012 18624
rect 7064 18612 7070 18624
rect 7469 18615 7527 18621
rect 7469 18612 7481 18615
rect 7064 18584 7481 18612
rect 7064 18572 7070 18584
rect 7469 18581 7481 18584
rect 7515 18581 7527 18615
rect 7469 18575 7527 18581
rect 7834 18572 7840 18624
rect 7892 18612 7898 18624
rect 8573 18615 8631 18621
rect 8573 18612 8585 18615
rect 7892 18584 8585 18612
rect 7892 18572 7898 18584
rect 8573 18581 8585 18584
rect 8619 18581 8631 18615
rect 8573 18575 8631 18581
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 11330 18612 11336 18624
rect 9723 18584 11336 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 12342 18572 12348 18624
rect 12400 18612 12406 18624
rect 14645 18615 14703 18621
rect 14645 18612 14657 18615
rect 12400 18584 14657 18612
rect 12400 18572 12406 18584
rect 14645 18581 14657 18584
rect 14691 18612 14703 18615
rect 16666 18612 16672 18624
rect 14691 18584 16672 18612
rect 14691 18581 14703 18584
rect 14645 18575 14703 18581
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 16850 18572 16856 18624
rect 16908 18612 16914 18624
rect 17144 18612 17172 18652
rect 19150 18640 19156 18652
rect 19208 18640 19214 18692
rect 20806 18680 20812 18692
rect 19628 18652 20812 18680
rect 16908 18584 17172 18612
rect 16908 18572 16914 18584
rect 17586 18572 17592 18624
rect 17644 18572 17650 18624
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 18414 18612 18420 18624
rect 17828 18584 18420 18612
rect 17828 18572 17834 18584
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 18506 18572 18512 18624
rect 18564 18572 18570 18624
rect 18782 18572 18788 18624
rect 18840 18612 18846 18624
rect 19628 18612 19656 18652
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 18840 18584 19656 18612
rect 18840 18572 18846 18584
rect 19702 18572 19708 18624
rect 19760 18572 19766 18624
rect 21450 18572 21456 18624
rect 21508 18612 21514 18624
rect 21652 18612 21680 18734
rect 21744 18720 22744 18748
rect 22738 18708 22744 18720
rect 22796 18708 22802 18760
rect 22830 18708 22836 18760
rect 22888 18748 22894 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22888 18720 22937 18748
rect 22888 18708 22894 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 23124 18748 23152 18779
rect 25038 18776 25044 18828
rect 25096 18776 25102 18828
rect 25130 18776 25136 18828
rect 25188 18776 25194 18828
rect 25314 18748 25320 18760
rect 23124 18720 25320 18748
rect 22925 18711 22983 18717
rect 25314 18708 25320 18720
rect 25372 18708 25378 18760
rect 22186 18640 22192 18692
rect 22244 18680 22250 18692
rect 23753 18683 23811 18689
rect 22244 18652 22876 18680
rect 22244 18640 22250 18652
rect 21508 18584 21680 18612
rect 21508 18572 21514 18584
rect 21910 18572 21916 18624
rect 21968 18612 21974 18624
rect 22005 18615 22063 18621
rect 22005 18612 22017 18615
rect 21968 18584 22017 18612
rect 21968 18572 21974 18584
rect 22005 18581 22017 18584
rect 22051 18581 22063 18615
rect 22005 18575 22063 18581
rect 22465 18615 22523 18621
rect 22465 18581 22477 18615
rect 22511 18612 22523 18615
rect 22646 18612 22652 18624
rect 22511 18584 22652 18612
rect 22511 18581 22523 18584
rect 22465 18575 22523 18581
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 22848 18621 22876 18652
rect 23753 18649 23765 18683
rect 23799 18680 23811 18683
rect 24670 18680 24676 18692
rect 23799 18652 24676 18680
rect 23799 18649 23811 18652
rect 23753 18643 23811 18649
rect 24670 18640 24676 18652
rect 24728 18640 24734 18692
rect 22833 18615 22891 18621
rect 22833 18581 22845 18615
rect 22879 18581 22891 18615
rect 22833 18575 22891 18581
rect 24578 18572 24584 18624
rect 24636 18572 24642 18624
rect 24946 18572 24952 18624
rect 25004 18572 25010 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 3789 18411 3847 18417
rect 3789 18408 3801 18411
rect 1728 18380 3801 18408
rect 1728 18368 1734 18380
rect 3789 18377 3801 18380
rect 3835 18377 3847 18411
rect 3789 18371 3847 18377
rect 5994 18368 6000 18420
rect 6052 18368 6058 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 6236 18380 6377 18408
rect 6236 18368 6242 18380
rect 6365 18377 6377 18380
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 6822 18368 6828 18420
rect 6880 18408 6886 18420
rect 10689 18411 10747 18417
rect 10689 18408 10701 18411
rect 6880 18380 10701 18408
rect 6880 18368 6886 18380
rect 10689 18377 10701 18380
rect 10735 18408 10747 18411
rect 14090 18408 14096 18420
rect 10735 18380 14096 18408
rect 10735 18377 10747 18380
rect 10689 18371 10747 18377
rect 14090 18368 14096 18380
rect 14148 18368 14154 18420
rect 14274 18368 14280 18420
rect 14332 18368 14338 18420
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 15013 18411 15071 18417
rect 15013 18408 15025 18411
rect 14884 18380 15025 18408
rect 14884 18368 14890 18380
rect 15013 18377 15025 18380
rect 15059 18377 15071 18411
rect 15013 18371 15071 18377
rect 15289 18411 15347 18417
rect 15289 18377 15301 18411
rect 15335 18408 15347 18411
rect 16025 18411 16083 18417
rect 16025 18408 16037 18411
rect 15335 18380 16037 18408
rect 15335 18377 15347 18380
rect 15289 18371 15347 18377
rect 16025 18377 16037 18380
rect 16071 18408 16083 18411
rect 16114 18408 16120 18420
rect 16071 18380 16120 18408
rect 16071 18377 16083 18380
rect 16025 18371 16083 18377
rect 16114 18368 16120 18380
rect 16172 18368 16178 18420
rect 16666 18368 16672 18420
rect 16724 18368 16730 18420
rect 18340 18380 20392 18408
rect 18340 18352 18368 18380
rect 4893 18343 4951 18349
rect 4893 18340 4905 18343
rect 2056 18312 4905 18340
rect 2056 18281 2084 18312
rect 4893 18309 4905 18312
rect 4939 18309 4951 18343
rect 4893 18303 4951 18309
rect 5258 18300 5264 18352
rect 5316 18340 5322 18352
rect 9217 18343 9275 18349
rect 9217 18340 9229 18343
rect 5316 18312 9229 18340
rect 5316 18300 5322 18312
rect 9217 18309 9229 18312
rect 9263 18309 9275 18343
rect 9217 18303 9275 18309
rect 12250 18300 12256 18352
rect 12308 18340 12314 18352
rect 12989 18343 13047 18349
rect 12989 18340 13001 18343
rect 12308 18312 13001 18340
rect 12308 18300 12314 18312
rect 12989 18309 13001 18312
rect 13035 18340 13047 18343
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 13035 18312 18245 18340
rect 13035 18309 13047 18312
rect 12989 18303 13047 18309
rect 18233 18309 18245 18312
rect 18279 18340 18291 18343
rect 18322 18340 18328 18352
rect 18279 18312 18328 18340
rect 18279 18309 18291 18312
rect 18233 18303 18291 18309
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 18874 18340 18880 18352
rect 18472 18312 18880 18340
rect 18472 18300 18478 18312
rect 18874 18300 18880 18312
rect 18932 18300 18938 18352
rect 19981 18343 20039 18349
rect 19981 18309 19993 18343
rect 20027 18340 20039 18343
rect 20254 18340 20260 18352
rect 20027 18312 20260 18340
rect 20027 18309 20039 18312
rect 19981 18303 20039 18309
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 20364 18340 20392 18380
rect 20530 18368 20536 18420
rect 20588 18408 20594 18420
rect 20588 18380 22416 18408
rect 20588 18368 20594 18380
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 20364 18312 22017 18340
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22388 18340 22416 18380
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 23290 18408 23296 18420
rect 22520 18380 23296 18408
rect 22520 18368 22526 18380
rect 23290 18368 23296 18380
rect 23348 18368 23354 18420
rect 24857 18411 24915 18417
rect 24857 18377 24869 18411
rect 24903 18408 24915 18411
rect 25866 18408 25872 18420
rect 24903 18380 25872 18408
rect 24903 18377 24915 18380
rect 24857 18371 24915 18377
rect 25866 18368 25872 18380
rect 25924 18368 25930 18420
rect 22388 18312 24256 18340
rect 22005 18303 22063 18309
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 3145 18275 3203 18281
rect 3145 18241 3157 18275
rect 3191 18272 3203 18275
rect 3878 18272 3884 18284
rect 3191 18244 3884 18272
rect 3191 18241 3203 18244
rect 3145 18235 3203 18241
rect 3878 18232 3884 18244
rect 3936 18232 3942 18284
rect 4246 18232 4252 18284
rect 4304 18232 4310 18284
rect 5350 18232 5356 18284
rect 5408 18232 5414 18284
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 6914 18272 6920 18284
rect 6779 18244 6920 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7300 18244 7512 18272
rect 2685 18207 2743 18213
rect 2685 18173 2697 18207
rect 2731 18204 2743 18207
rect 7300 18204 7328 18244
rect 2731 18176 7328 18204
rect 2731 18173 2743 18176
rect 2685 18167 2743 18173
rect 7374 18164 7380 18216
rect 7432 18164 7438 18216
rect 7484 18204 7512 18244
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 8938 18232 8944 18284
rect 8996 18232 9002 18284
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 10502 18272 10508 18284
rect 10376 18244 10508 18272
rect 10376 18232 10382 18244
rect 10502 18232 10508 18244
rect 10560 18232 10566 18284
rect 11146 18232 11152 18284
rect 11204 18272 11210 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 11204 18244 12173 18272
rect 11204 18232 11210 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 13078 18232 13084 18284
rect 13136 18272 13142 18284
rect 13814 18272 13820 18284
rect 13136 18244 13820 18272
rect 13136 18232 13142 18244
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 14240 18244 15945 18272
rect 14240 18232 14246 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 17126 18272 17132 18284
rect 15933 18235 15991 18241
rect 16021 18244 17132 18272
rect 7484 18176 10272 18204
rect 6914 18096 6920 18148
rect 6972 18136 6978 18148
rect 7392 18136 7420 18164
rect 6972 18108 7420 18136
rect 10244 18136 10272 18176
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 11241 18207 11299 18213
rect 11241 18204 11253 18207
rect 11112 18176 11253 18204
rect 11112 18164 11118 18176
rect 11241 18173 11253 18176
rect 11287 18173 11299 18207
rect 11790 18204 11796 18216
rect 11241 18167 11299 18173
rect 11348 18176 11796 18204
rect 11348 18136 11376 18176
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 10244 18108 11376 18136
rect 12268 18136 12296 18167
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 13262 18204 13268 18216
rect 12676 18176 13268 18204
rect 12676 18164 12682 18176
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 15654 18204 15660 18216
rect 13504 18176 15660 18204
rect 13504 18164 13510 18176
rect 15654 18164 15660 18176
rect 15712 18164 15718 18216
rect 15746 18164 15752 18216
rect 15804 18204 15810 18216
rect 16021 18204 16049 18244
rect 17126 18232 17132 18244
rect 17184 18272 17190 18284
rect 17405 18275 17463 18281
rect 17405 18272 17417 18275
rect 17184 18244 17417 18272
rect 17184 18232 17190 18244
rect 17405 18241 17417 18244
rect 17451 18241 17463 18275
rect 17405 18235 17463 18241
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 20530 18272 20536 18284
rect 19484 18244 20536 18272
rect 19484 18232 19490 18244
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 20806 18232 20812 18284
rect 20864 18232 20870 18284
rect 20901 18275 20959 18281
rect 20901 18241 20913 18275
rect 20947 18272 20959 18275
rect 21082 18272 21088 18284
rect 20947 18244 21088 18272
rect 20947 18241 20959 18244
rect 20901 18235 20959 18241
rect 21082 18232 21088 18244
rect 21140 18272 21146 18284
rect 24228 18281 24256 18312
rect 25314 18300 25320 18352
rect 25372 18300 25378 18352
rect 21453 18275 21511 18281
rect 21453 18272 21465 18275
rect 21140 18244 21465 18272
rect 21140 18232 21146 18244
rect 21453 18241 21465 18244
rect 21499 18241 21511 18275
rect 21453 18235 21511 18241
rect 24213 18275 24271 18281
rect 24213 18241 24225 18275
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 25590 18232 25596 18284
rect 25648 18272 25654 18284
rect 25866 18272 25872 18284
rect 25648 18244 25872 18272
rect 25648 18232 25654 18244
rect 25866 18232 25872 18244
rect 25924 18232 25930 18284
rect 15804 18176 16049 18204
rect 15804 18164 15810 18176
rect 16114 18164 16120 18216
rect 16172 18164 16178 18216
rect 16482 18164 16488 18216
rect 16540 18204 16546 18216
rect 17497 18207 17555 18213
rect 17497 18204 17509 18207
rect 16540 18176 17509 18204
rect 16540 18164 16546 18176
rect 17497 18173 17509 18176
rect 17543 18204 17555 18207
rect 17586 18204 17592 18216
rect 17543 18176 17592 18204
rect 17543 18173 17555 18176
rect 17497 18167 17555 18173
rect 17586 18164 17592 18176
rect 17644 18164 17650 18216
rect 17681 18207 17739 18213
rect 17681 18173 17693 18207
rect 17727 18204 17739 18207
rect 17770 18204 17776 18216
rect 17727 18176 17776 18204
rect 17727 18173 17739 18176
rect 17681 18167 17739 18173
rect 17770 18164 17776 18176
rect 17828 18164 17834 18216
rect 17862 18164 17868 18216
rect 17920 18204 17926 18216
rect 20714 18204 20720 18216
rect 17920 18176 20720 18204
rect 17920 18164 17926 18176
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 20993 18207 21051 18213
rect 20993 18173 21005 18207
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 15565 18139 15623 18145
rect 15565 18136 15577 18139
rect 12268 18108 15577 18136
rect 6972 18096 6978 18108
rect 15565 18105 15577 18108
rect 15611 18105 15623 18139
rect 15565 18099 15623 18105
rect 16390 18096 16396 18148
rect 16448 18136 16454 18148
rect 16448 18108 19104 18136
rect 16448 18096 16454 18108
rect 1670 18028 1676 18080
rect 1728 18028 1734 18080
rect 7374 18028 7380 18080
rect 7432 18028 7438 18080
rect 8478 18028 8484 18080
rect 8536 18028 8542 18080
rect 8662 18028 8668 18080
rect 8720 18068 8726 18080
rect 9306 18068 9312 18080
rect 8720 18040 9312 18068
rect 8720 18028 8726 18040
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 11149 18071 11207 18077
rect 11149 18037 11161 18071
rect 11195 18068 11207 18071
rect 11514 18068 11520 18080
rect 11195 18040 11520 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 11790 18028 11796 18080
rect 11848 18028 11854 18080
rect 12250 18028 12256 18080
rect 12308 18068 12314 18080
rect 13170 18068 13176 18080
rect 12308 18040 13176 18068
rect 12308 18028 12314 18040
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 14642 18068 14648 18080
rect 13964 18040 14648 18068
rect 13964 18028 13970 18040
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 16482 18068 16488 18080
rect 15712 18040 16488 18068
rect 15712 18028 15718 18040
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 17037 18071 17095 18077
rect 17037 18037 17049 18071
rect 17083 18068 17095 18071
rect 18414 18068 18420 18080
rect 17083 18040 18420 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 19076 18068 19104 18108
rect 19150 18096 19156 18148
rect 19208 18136 19214 18148
rect 21008 18136 21036 18167
rect 19208 18108 21036 18136
rect 19208 18096 19214 18108
rect 24762 18096 24768 18148
rect 24820 18136 24826 18148
rect 25133 18139 25191 18145
rect 25133 18136 25145 18139
rect 24820 18108 25145 18136
rect 24820 18096 24826 18108
rect 25133 18105 25145 18108
rect 25179 18105 25191 18139
rect 25133 18099 25191 18105
rect 19518 18068 19524 18080
rect 19076 18040 19524 18068
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 20441 18071 20499 18077
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 20622 18068 20628 18080
rect 20487 18040 20628 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 22922 18028 22928 18080
rect 22980 18068 22986 18080
rect 24394 18068 24400 18080
rect 22980 18040 24400 18068
rect 22980 18028 22986 18040
rect 24394 18028 24400 18040
rect 24452 18028 24458 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 2363 17836 4568 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 3970 17756 3976 17808
rect 4028 17756 4034 17808
rect 4540 17796 4568 17836
rect 4614 17824 4620 17876
rect 4672 17864 4678 17876
rect 5261 17867 5319 17873
rect 5261 17864 5273 17867
rect 4672 17836 5273 17864
rect 4672 17824 4678 17836
rect 5261 17833 5273 17836
rect 5307 17833 5319 17867
rect 5261 17827 5319 17833
rect 5350 17824 5356 17876
rect 5408 17864 5414 17876
rect 6365 17867 6423 17873
rect 6365 17864 6377 17867
rect 5408 17836 6377 17864
rect 5408 17824 5414 17836
rect 6365 17833 6377 17836
rect 6411 17833 6423 17867
rect 6914 17864 6920 17876
rect 6365 17827 6423 17833
rect 6472 17836 6920 17864
rect 6472 17796 6500 17836
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7432 17836 10824 17864
rect 7432 17824 7438 17836
rect 4540 17768 6500 17796
rect 6730 17756 6736 17808
rect 6788 17796 6794 17808
rect 6788 17768 7972 17796
rect 6788 17756 6794 17768
rect 3418 17688 3424 17740
rect 3476 17728 3482 17740
rect 7944 17728 7972 17768
rect 8202 17756 8208 17808
rect 8260 17796 8266 17808
rect 9122 17796 9128 17808
rect 8260 17768 9128 17796
rect 8260 17756 8266 17768
rect 9122 17756 9128 17768
rect 9180 17756 9186 17808
rect 10796 17796 10824 17836
rect 11238 17824 11244 17876
rect 11296 17824 11302 17876
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 12342 17864 12348 17876
rect 12124 17836 12348 17864
rect 12124 17824 12130 17836
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13449 17867 13507 17873
rect 13449 17864 13461 17867
rect 12492 17836 13461 17864
rect 12492 17824 12498 17836
rect 13449 17833 13461 17836
rect 13495 17833 13507 17867
rect 13449 17827 13507 17833
rect 13538 17824 13544 17876
rect 13596 17864 13602 17876
rect 13909 17867 13967 17873
rect 13909 17864 13921 17867
rect 13596 17836 13921 17864
rect 13596 17824 13602 17836
rect 13909 17833 13921 17836
rect 13955 17864 13967 17867
rect 15746 17864 15752 17876
rect 13955 17836 15752 17864
rect 13955 17833 13967 17836
rect 13909 17827 13967 17833
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 16574 17864 16580 17876
rect 15896 17836 16580 17864
rect 15896 17824 15902 17836
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 17129 17867 17187 17873
rect 17129 17864 17141 17867
rect 17000 17836 17141 17864
rect 17000 17824 17006 17836
rect 17129 17833 17141 17836
rect 17175 17833 17187 17867
rect 17129 17827 17187 17833
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17402 17864 17408 17876
rect 17276 17836 17408 17864
rect 17276 17824 17282 17836
rect 17402 17824 17408 17836
rect 17460 17824 17466 17876
rect 17586 17824 17592 17876
rect 17644 17864 17650 17876
rect 17644 17836 24624 17864
rect 17644 17824 17650 17836
rect 16669 17799 16727 17805
rect 10796 17768 11836 17796
rect 8294 17728 8300 17740
rect 3476 17700 4660 17728
rect 7944 17700 8300 17728
rect 3476 17688 3482 17700
rect 1670 17620 1676 17672
rect 1728 17620 1734 17672
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17660 2835 17663
rect 3786 17660 3792 17672
rect 2823 17632 3792 17660
rect 2823 17629 2835 17632
rect 2777 17623 2835 17629
rect 3786 17620 3792 17632
rect 3844 17620 3850 17672
rect 4632 17669 4660 17700
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 8573 17731 8631 17737
rect 8573 17697 8585 17731
rect 8619 17728 8631 17731
rect 8846 17728 8852 17740
rect 8619 17700 8852 17728
rect 8619 17697 8631 17700
rect 8573 17691 8631 17697
rect 8846 17688 8852 17700
rect 8904 17688 8910 17740
rect 8938 17688 8944 17740
rect 8996 17728 9002 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 8996 17700 9505 17728
rect 8996 17688 9002 17700
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 4617 17663 4675 17669
rect 4617 17629 4629 17663
rect 4663 17629 4675 17663
rect 4617 17623 4675 17629
rect 3418 17552 3424 17604
rect 3476 17552 3482 17604
rect 4172 17592 4200 17623
rect 5718 17620 5724 17672
rect 5776 17620 5782 17672
rect 6178 17660 6184 17672
rect 5828 17632 6184 17660
rect 5828 17592 5856 17632
rect 6178 17620 6184 17632
rect 6236 17620 6242 17672
rect 6825 17663 6883 17669
rect 6825 17629 6837 17663
rect 6871 17660 6883 17663
rect 7650 17660 7656 17672
rect 6871 17632 7656 17660
rect 6871 17629 6883 17632
rect 6825 17623 6883 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 8662 17660 8668 17672
rect 7975 17632 8668 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 9048 17648 9137 17660
rect 9030 17596 9036 17648
rect 9088 17632 9137 17648
rect 9088 17596 9094 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9125 17623 9183 17629
rect 4172 17564 5856 17592
rect 9232 17536 9260 17700
rect 9493 17697 9505 17700
rect 9539 17728 9551 17731
rect 11698 17728 11704 17740
rect 9539 17700 11704 17728
rect 9539 17697 9551 17700
rect 9493 17691 9551 17697
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11808 17728 11836 17768
rect 16669 17765 16681 17799
rect 16715 17796 16727 17799
rect 19426 17796 19432 17808
rect 16715 17768 19432 17796
rect 16715 17765 16727 17768
rect 16669 17759 16727 17765
rect 19426 17756 19432 17768
rect 19484 17756 19490 17808
rect 22094 17756 22100 17808
rect 22152 17756 22158 17808
rect 22186 17756 22192 17808
rect 22244 17796 22250 17808
rect 22465 17799 22523 17805
rect 22465 17796 22477 17799
rect 22244 17768 22477 17796
rect 22244 17756 22250 17768
rect 22465 17765 22477 17768
rect 22511 17765 22523 17799
rect 22465 17759 22523 17765
rect 22830 17756 22836 17808
rect 22888 17756 22894 17808
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11808 17700 11989 17728
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12066 17688 12072 17740
rect 12124 17728 12130 17740
rect 12434 17728 12440 17740
rect 12124 17700 12440 17728
rect 12124 17688 12130 17700
rect 12434 17688 12440 17700
rect 12492 17688 12498 17740
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 14182 17728 14188 17740
rect 12676 17700 14188 17728
rect 12676 17688 12682 17700
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 14921 17731 14979 17737
rect 14921 17728 14933 17731
rect 14332 17700 14933 17728
rect 14332 17688 14338 17700
rect 14921 17697 14933 17700
rect 14967 17697 14979 17731
rect 14921 17691 14979 17697
rect 15197 17731 15255 17737
rect 15197 17697 15209 17731
rect 15243 17728 15255 17731
rect 15286 17728 15292 17740
rect 15243 17700 15292 17728
rect 15243 17697 15255 17700
rect 15197 17691 15255 17697
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 16758 17688 16764 17740
rect 16816 17728 16822 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 16816 17700 17693 17728
rect 16816 17688 16822 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 18325 17731 18383 17737
rect 18325 17697 18337 17731
rect 18371 17728 18383 17731
rect 18598 17728 18604 17740
rect 18371 17700 18604 17728
rect 18371 17697 18383 17700
rect 18325 17691 18383 17697
rect 18598 17688 18604 17700
rect 18656 17688 18662 17740
rect 18874 17688 18880 17740
rect 18932 17688 18938 17740
rect 21634 17728 21640 17740
rect 19536 17700 21640 17728
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 14734 17660 14740 17672
rect 13688 17632 14740 17660
rect 13688 17620 13694 17632
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 16592 17632 17724 17660
rect 9769 17595 9827 17601
rect 9769 17592 9781 17595
rect 9646 17564 9781 17592
rect 9646 17536 9674 17564
rect 9769 17561 9781 17564
rect 9815 17561 9827 17595
rect 9769 17555 9827 17561
rect 10318 17552 10324 17604
rect 10376 17552 10382 17604
rect 12066 17592 12072 17604
rect 11164 17564 12072 17592
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 5902 17524 5908 17536
rect 2096 17496 5908 17524
rect 2096 17484 2102 17496
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 7466 17484 7472 17536
rect 7524 17484 7530 17536
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 8941 17527 8999 17533
rect 8941 17524 8953 17527
rect 8628 17496 8953 17524
rect 8628 17484 8634 17496
rect 8941 17493 8953 17496
rect 8987 17493 8999 17527
rect 8941 17487 8999 17493
rect 9214 17484 9220 17536
rect 9272 17484 9278 17536
rect 9582 17484 9588 17536
rect 9640 17496 9674 17536
rect 9640 17484 9646 17496
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 11164 17524 11192 17564
rect 12066 17552 12072 17564
rect 12124 17552 12130 17604
rect 13262 17592 13268 17604
rect 13202 17564 13268 17592
rect 13262 17552 13268 17564
rect 13320 17552 13326 17604
rect 13354 17552 13360 17604
rect 13412 17592 13418 17604
rect 14277 17595 14335 17601
rect 14277 17592 14289 17595
rect 13412 17564 14289 17592
rect 13412 17552 13418 17564
rect 14277 17561 14289 17564
rect 14323 17561 14335 17595
rect 14277 17555 14335 17561
rect 15838 17552 15844 17604
rect 15896 17552 15902 17604
rect 10560 17496 11192 17524
rect 10560 17484 10566 17496
rect 11238 17484 11244 17536
rect 11296 17524 11302 17536
rect 16592 17524 16620 17632
rect 16666 17552 16672 17604
rect 16724 17592 16730 17604
rect 17589 17595 17647 17601
rect 17589 17592 17601 17595
rect 16724 17564 17601 17592
rect 16724 17552 16730 17564
rect 17589 17561 17601 17564
rect 17635 17561 17647 17595
rect 17589 17555 17647 17561
rect 11296 17496 16620 17524
rect 11296 17484 11302 17496
rect 16942 17484 16948 17536
rect 17000 17524 17006 17536
rect 17497 17527 17555 17533
rect 17497 17524 17509 17527
rect 17000 17496 17509 17524
rect 17000 17484 17006 17496
rect 17497 17493 17509 17496
rect 17543 17493 17555 17527
rect 17696 17524 17724 17632
rect 19058 17620 19064 17672
rect 19116 17660 19122 17672
rect 19536 17669 19564 17700
rect 21634 17688 21640 17700
rect 21692 17688 21698 17740
rect 22112 17728 22140 17756
rect 22925 17731 22983 17737
rect 22925 17728 22937 17731
rect 22112 17700 22937 17728
rect 22925 17697 22937 17700
rect 22971 17697 22983 17731
rect 22925 17691 22983 17697
rect 23937 17731 23995 17737
rect 23937 17697 23949 17731
rect 23983 17728 23995 17731
rect 24026 17728 24032 17740
rect 23983 17700 24032 17728
rect 23983 17697 23995 17700
rect 23937 17691 23995 17697
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 19521 17663 19579 17669
rect 19521 17660 19533 17663
rect 19116 17632 19533 17660
rect 19116 17620 19122 17632
rect 19521 17629 19533 17632
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 19978 17620 19984 17672
rect 20036 17620 20042 17672
rect 20714 17620 20720 17672
rect 20772 17620 20778 17672
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 24486 17660 24492 17672
rect 23799 17632 24492 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 24486 17620 24492 17632
rect 24544 17620 24550 17672
rect 24596 17669 24624 17836
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17629 24639 17663
rect 24581 17623 24639 17629
rect 18414 17552 18420 17604
rect 18472 17592 18478 17604
rect 20732 17592 20760 17620
rect 18472 17564 20760 17592
rect 18472 17552 18478 17564
rect 20990 17552 20996 17604
rect 21048 17552 21054 17604
rect 21450 17552 21456 17604
rect 21508 17552 21514 17604
rect 23661 17595 23719 17601
rect 23661 17561 23673 17595
rect 23707 17592 23719 17595
rect 23842 17592 23848 17604
rect 23707 17564 23848 17592
rect 23707 17561 23719 17564
rect 23661 17555 23719 17561
rect 23842 17552 23848 17564
rect 23900 17552 23906 17604
rect 22278 17524 22284 17536
rect 17696 17496 22284 17524
rect 17497 17487 17555 17493
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 23290 17484 23296 17536
rect 23348 17484 23354 17536
rect 24946 17484 24952 17536
rect 25004 17524 25010 17536
rect 25225 17527 25283 17533
rect 25225 17524 25237 17527
rect 25004 17496 25237 17524
rect 25004 17484 25010 17496
rect 25225 17493 25237 17496
rect 25271 17493 25283 17527
rect 25225 17487 25283 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 2682 17280 2688 17332
rect 2740 17280 2746 17332
rect 3786 17280 3792 17332
rect 3844 17280 3850 17332
rect 6454 17280 6460 17332
rect 6512 17320 6518 17332
rect 7282 17320 7288 17332
rect 6512 17292 7288 17320
rect 6512 17280 6518 17292
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 7374 17280 7380 17332
rect 7432 17280 7438 17332
rect 7650 17280 7656 17332
rect 7708 17280 7714 17332
rect 8757 17323 8815 17329
rect 8757 17289 8769 17323
rect 8803 17320 8815 17323
rect 8803 17292 10824 17320
rect 8803 17289 8815 17292
rect 8757 17283 8815 17289
rect 1765 17255 1823 17261
rect 1765 17221 1777 17255
rect 1811 17252 1823 17255
rect 4893 17255 4951 17261
rect 1811 17224 3188 17252
rect 1811 17221 1823 17224
rect 1765 17215 1823 17221
rect 3160 17193 3188 17224
rect 4893 17221 4905 17255
rect 4939 17252 4951 17255
rect 6730 17252 6736 17264
rect 4939 17224 6736 17252
rect 4939 17221 4951 17224
rect 4893 17215 4951 17221
rect 6730 17212 6736 17224
rect 6788 17212 6794 17264
rect 7392 17252 7420 17280
rect 7208 17224 7420 17252
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17153 2099 17187
rect 2041 17147 2099 17153
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17184 3203 17187
rect 3418 17184 3424 17196
rect 3191 17156 3424 17184
rect 3191 17153 3203 17156
rect 3145 17147 3203 17153
rect 2056 17116 2084 17147
rect 3418 17144 3424 17156
rect 3476 17144 3482 17196
rect 4246 17144 4252 17196
rect 4304 17144 4310 17196
rect 5350 17144 5356 17196
rect 5408 17144 5414 17196
rect 7006 17144 7012 17196
rect 7064 17144 7070 17196
rect 7208 17128 7236 17224
rect 7466 17212 7472 17264
rect 7524 17252 7530 17264
rect 9493 17255 9551 17261
rect 9493 17252 9505 17255
rect 7524 17224 9505 17252
rect 7524 17212 7530 17224
rect 9493 17221 9505 17224
rect 9539 17221 9551 17255
rect 9493 17215 9551 17221
rect 10502 17212 10508 17264
rect 10560 17212 10566 17264
rect 10796 17252 10824 17292
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 14642 17320 14648 17332
rect 11388 17292 14648 17320
rect 11388 17280 11394 17292
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17289 14795 17323
rect 14737 17283 14795 17289
rect 12805 17255 12863 17261
rect 12805 17252 12817 17255
rect 10796 17224 12817 17252
rect 12805 17221 12817 17224
rect 12851 17221 12863 17255
rect 12805 17215 12863 17221
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 14752 17252 14780 17283
rect 15470 17280 15476 17332
rect 15528 17280 15534 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 15620 17292 20024 17320
rect 15620 17280 15626 17292
rect 15488 17252 15516 17280
rect 14240 17224 14780 17252
rect 15120 17224 15516 17252
rect 15841 17255 15899 17261
rect 14240 17212 14246 17224
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17184 8171 17187
rect 8478 17184 8484 17196
rect 8159 17156 8484 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 9214 17144 9220 17196
rect 9272 17144 9278 17196
rect 11882 17144 11888 17196
rect 11940 17144 11946 17196
rect 14090 17184 14096 17196
rect 13938 17156 14096 17184
rect 14090 17144 14096 17156
rect 14148 17184 14154 17196
rect 14921 17187 14979 17193
rect 14148 17156 14872 17184
rect 14148 17144 14154 17156
rect 5902 17116 5908 17128
rect 2056 17088 5908 17116
rect 5902 17076 5908 17088
rect 5960 17076 5966 17128
rect 7190 17076 7196 17128
rect 7248 17076 7254 17128
rect 8680 17088 9352 17116
rect 5626 17008 5632 17060
rect 5684 17048 5690 17060
rect 7834 17048 7840 17060
rect 5684 17020 7840 17048
rect 5684 17008 5690 17020
rect 7834 17008 7840 17020
rect 7892 17008 7898 17060
rect 8110 17008 8116 17060
rect 8168 17048 8174 17060
rect 8680 17048 8708 17088
rect 8168 17020 8708 17048
rect 8168 17008 8174 17020
rect 5994 16940 6000 16992
rect 6052 16940 6058 16992
rect 6730 16940 6736 16992
rect 6788 16980 6794 16992
rect 9214 16980 9220 16992
rect 6788 16952 9220 16980
rect 6788 16940 6794 16952
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 9324 16980 9352 17088
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 9548 17088 11652 17116
rect 9548 17076 9554 17088
rect 10686 17008 10692 17060
rect 10744 17048 10750 17060
rect 11238 17048 11244 17060
rect 10744 17020 11244 17048
rect 10744 17008 10750 17020
rect 11238 17008 11244 17020
rect 11296 17008 11302 17060
rect 10594 16980 10600 16992
rect 9324 16952 10600 16980
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 10962 16940 10968 16992
rect 11020 16940 11026 16992
rect 11624 16980 11652 17088
rect 11698 17076 11704 17128
rect 11756 17116 11762 17128
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 11756 17088 12541 17116
rect 11756 17076 11762 17088
rect 12529 17085 12541 17088
rect 12575 17085 12587 17119
rect 13354 17116 13360 17128
rect 12529 17079 12587 17085
rect 12636 17088 13360 17116
rect 12066 17008 12072 17060
rect 12124 17008 12130 17060
rect 12434 17008 12440 17060
rect 12492 17048 12498 17060
rect 12636 17048 12664 17088
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 13446 17076 13452 17128
rect 13504 17116 13510 17128
rect 14844 17116 14872 17156
rect 14921 17153 14933 17187
rect 14967 17184 14979 17187
rect 15120 17184 15148 17224
rect 15841 17221 15853 17255
rect 15887 17252 15899 17255
rect 16485 17255 16543 17261
rect 16485 17252 16497 17255
rect 15887 17224 16497 17252
rect 15887 17221 15899 17224
rect 15841 17215 15899 17221
rect 16485 17221 16497 17224
rect 16531 17252 16543 17255
rect 16666 17252 16672 17264
rect 16531 17224 16672 17252
rect 16531 17221 16543 17224
rect 16485 17215 16543 17221
rect 16666 17212 16672 17224
rect 16724 17212 16730 17264
rect 17221 17255 17279 17261
rect 17221 17221 17233 17255
rect 17267 17252 17279 17255
rect 18598 17252 18604 17264
rect 17267 17224 18604 17252
rect 17267 17221 17279 17224
rect 17221 17215 17279 17221
rect 18598 17212 18604 17224
rect 18656 17212 18662 17264
rect 18690 17212 18696 17264
rect 18748 17212 18754 17264
rect 19996 17252 20024 17292
rect 20162 17280 20168 17332
rect 20220 17280 20226 17332
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 21269 17323 21327 17329
rect 21269 17320 21281 17323
rect 20864 17292 21281 17320
rect 20864 17280 20870 17292
rect 21269 17289 21281 17292
rect 21315 17289 21327 17323
rect 21269 17283 21327 17289
rect 22066 17292 23888 17320
rect 19996 17224 20668 17252
rect 14967 17156 15148 17184
rect 14967 17153 14979 17156
rect 14921 17147 14979 17153
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 15528 17156 15761 17184
rect 15528 17144 15534 17156
rect 15749 17153 15761 17156
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 16022 17144 16028 17196
rect 16080 17184 16086 17196
rect 17586 17184 17592 17196
rect 16080 17156 17592 17184
rect 16080 17144 16086 17156
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 18414 17144 18420 17196
rect 18472 17144 18478 17196
rect 19794 17144 19800 17196
rect 19852 17144 19858 17196
rect 20640 17193 20668 17224
rect 21450 17212 21456 17264
rect 21508 17252 21514 17264
rect 22066 17252 22094 17292
rect 21508 17224 22094 17252
rect 21508 17212 21514 17224
rect 23860 17196 23888 17292
rect 26234 17212 26240 17264
rect 26292 17252 26298 17264
rect 26786 17252 26792 17264
rect 26292 17224 26792 17252
rect 26292 17212 26298 17224
rect 26786 17212 26792 17224
rect 26844 17212 26850 17264
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 22462 17184 22468 17196
rect 20772 17156 22468 17184
rect 20772 17144 20778 17156
rect 22462 17144 22468 17156
rect 22520 17144 22526 17196
rect 23842 17144 23848 17196
rect 23900 17144 23906 17196
rect 24673 17187 24731 17193
rect 24673 17153 24685 17187
rect 24719 17184 24731 17187
rect 24762 17184 24768 17196
rect 24719 17156 24768 17184
rect 24719 17153 24731 17156
rect 24673 17147 24731 17153
rect 24762 17144 24768 17156
rect 24820 17144 24826 17196
rect 15838 17116 15844 17128
rect 13504 17088 14780 17116
rect 14844 17088 15844 17116
rect 13504 17076 13510 17088
rect 12492 17020 12664 17048
rect 14752 17048 14780 17088
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 15933 17119 15991 17125
rect 15933 17085 15945 17119
rect 15979 17085 15991 17119
rect 15933 17079 15991 17085
rect 15948 17048 15976 17079
rect 16206 17076 16212 17128
rect 16264 17116 16270 17128
rect 16850 17116 16856 17128
rect 16264 17088 16856 17116
rect 16264 17076 16270 17088
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 17052 17088 17325 17116
rect 14752 17020 15976 17048
rect 12492 17008 12498 17020
rect 13998 16980 14004 16992
rect 11624 16952 14004 16980
rect 13998 16940 14004 16952
rect 14056 16980 14062 16992
rect 14277 16983 14335 16989
rect 14277 16980 14289 16983
rect 14056 16952 14289 16980
rect 14056 16940 14062 16952
rect 14277 16949 14289 16952
rect 14323 16949 14335 16983
rect 14277 16943 14335 16949
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 15381 16983 15439 16989
rect 15381 16980 15393 16983
rect 14700 16952 15393 16980
rect 14700 16940 14706 16952
rect 15381 16949 15393 16952
rect 15427 16949 15439 16983
rect 15381 16943 15439 16949
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 16724 16952 16865 16980
rect 16724 16940 16730 16952
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 17052 16980 17080 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17405 17119 17463 17125
rect 17405 17085 17417 17119
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 17126 17008 17132 17060
rect 17184 17048 17190 17060
rect 17420 17048 17448 17079
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 18012 17088 18153 17116
rect 18012 17076 18018 17088
rect 18141 17085 18153 17088
rect 18187 17116 18199 17119
rect 19058 17116 19064 17128
rect 18187 17088 19064 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 19058 17076 19064 17088
rect 19116 17076 19122 17128
rect 19812 17116 19840 17144
rect 21450 17116 21456 17128
rect 19812 17088 21456 17116
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 22741 17119 22799 17125
rect 22741 17116 22753 17119
rect 22152 17088 22753 17116
rect 22152 17076 22158 17088
rect 22741 17085 22753 17088
rect 22787 17085 22799 17119
rect 22741 17079 22799 17085
rect 22830 17076 22836 17128
rect 22888 17116 22894 17128
rect 24026 17116 24032 17128
rect 22888 17088 24032 17116
rect 22888 17076 22894 17088
rect 24026 17076 24032 17088
rect 24084 17116 24090 17128
rect 24213 17119 24271 17125
rect 24213 17116 24225 17119
rect 24084 17088 24225 17116
rect 24084 17076 24090 17088
rect 24213 17085 24225 17088
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 17184 17020 17448 17048
rect 17184 17008 17190 17020
rect 20530 17008 20536 17060
rect 20588 17048 20594 17060
rect 25317 17051 25375 17057
rect 25317 17048 25329 17051
rect 20588 17020 22600 17048
rect 20588 17008 20594 17020
rect 17402 16980 17408 16992
rect 17052 16952 17408 16980
rect 16853 16943 16911 16949
rect 17402 16940 17408 16952
rect 17460 16980 17466 16992
rect 17865 16983 17923 16989
rect 17865 16980 17877 16983
rect 17460 16952 17877 16980
rect 17460 16940 17466 16952
rect 17865 16949 17877 16952
rect 17911 16980 17923 16983
rect 21450 16980 21456 16992
rect 17911 16952 21456 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 21450 16940 21456 16952
rect 21508 16980 21514 16992
rect 21545 16983 21603 16989
rect 21545 16980 21557 16983
rect 21508 16952 21557 16980
rect 21508 16940 21514 16952
rect 21545 16949 21557 16952
rect 21591 16949 21603 16983
rect 21545 16943 21603 16949
rect 22002 16940 22008 16992
rect 22060 16940 22066 16992
rect 22094 16940 22100 16992
rect 22152 16940 22158 16992
rect 22572 16980 22600 17020
rect 23768 17020 25329 17048
rect 23768 16980 23796 17020
rect 25317 17017 25329 17020
rect 25363 17017 25375 17051
rect 25317 17011 25375 17017
rect 22572 16952 23796 16980
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 4617 16779 4675 16785
rect 4617 16776 4629 16779
rect 4580 16748 4629 16776
rect 4580 16736 4586 16748
rect 4617 16745 4629 16748
rect 4663 16745 4675 16779
rect 4617 16739 4675 16745
rect 9030 16736 9036 16788
rect 9088 16776 9094 16788
rect 9088 16748 9168 16776
rect 9088 16736 9094 16748
rect 8846 16708 8852 16720
rect 6840 16680 8852 16708
rect 4062 16600 4068 16652
rect 4120 16600 4126 16652
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 2682 16572 2688 16584
rect 1719 16544 2688 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 2682 16532 2688 16544
rect 2740 16532 2746 16584
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16572 2835 16575
rect 3510 16572 3516 16584
rect 2823 16544 3516 16572
rect 2823 16541 2835 16544
rect 2777 16535 2835 16541
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16541 4031 16575
rect 4080 16572 4108 16600
rect 4430 16572 4436 16584
rect 4080 16544 4436 16572
rect 3973 16535 4031 16541
rect 3988 16504 4016 16535
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 5258 16532 5264 16584
rect 5316 16532 5322 16584
rect 5721 16575 5779 16581
rect 5721 16541 5733 16575
rect 5767 16572 5779 16575
rect 6178 16572 6184 16584
rect 5767 16544 6184 16572
rect 5767 16541 5779 16544
rect 5721 16535 5779 16541
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 6270 16532 6276 16584
rect 6328 16572 6334 16584
rect 6840 16581 6868 16680
rect 8846 16668 8852 16680
rect 8904 16668 8910 16720
rect 9140 16708 9168 16748
rect 9490 16736 9496 16788
rect 9548 16776 9554 16788
rect 23198 16776 23204 16788
rect 9548 16748 23204 16776
rect 9548 16736 9554 16748
rect 23198 16736 23204 16748
rect 23256 16736 23262 16788
rect 9674 16708 9680 16720
rect 9140 16680 9680 16708
rect 9674 16668 9680 16680
rect 9732 16668 9738 16720
rect 11256 16680 11468 16708
rect 8662 16640 8668 16652
rect 8266 16612 8668 16640
rect 6365 16575 6423 16581
rect 6365 16572 6377 16575
rect 6328 16544 6377 16572
rect 6328 16532 6334 16544
rect 6365 16541 6377 16544
rect 6411 16541 6423 16575
rect 6365 16535 6423 16541
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16572 7987 16575
rect 8266 16572 8294 16612
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 8754 16600 8760 16652
rect 8812 16600 8818 16652
rect 11256 16649 11284 16680
rect 9033 16643 9091 16649
rect 9033 16609 9045 16643
rect 9079 16640 9091 16643
rect 11241 16643 11299 16649
rect 9079 16612 11192 16640
rect 9079 16609 9091 16612
rect 9033 16603 9091 16609
rect 7975 16544 8294 16572
rect 7975 16541 7987 16544
rect 7929 16535 7987 16541
rect 2746 16476 4016 16504
rect 2314 16396 2320 16448
rect 2372 16396 2378 16448
rect 2406 16396 2412 16448
rect 2464 16436 2470 16448
rect 2746 16436 2774 16476
rect 4062 16464 4068 16516
rect 4120 16504 4126 16516
rect 5166 16504 5172 16516
rect 4120 16476 5172 16504
rect 4120 16464 4126 16476
rect 5166 16464 5172 16476
rect 5224 16464 5230 16516
rect 7098 16464 7104 16516
rect 7156 16504 7162 16516
rect 8110 16504 8116 16516
rect 7156 16476 8116 16504
rect 7156 16464 7162 16476
rect 8110 16464 8116 16476
rect 8168 16464 8174 16516
rect 8202 16464 8208 16516
rect 8260 16504 8266 16516
rect 8478 16504 8484 16516
rect 8260 16476 8484 16504
rect 8260 16464 8266 16476
rect 8478 16464 8484 16476
rect 8536 16464 8542 16516
rect 8772 16504 8800 16600
rect 9674 16532 9680 16584
rect 9732 16532 9738 16584
rect 11164 16572 11192 16612
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 11330 16600 11336 16652
rect 11388 16600 11394 16652
rect 11440 16640 11468 16680
rect 13998 16668 14004 16720
rect 14056 16708 14062 16720
rect 14056 16680 14412 16708
rect 14056 16668 14062 16680
rect 13722 16640 13728 16652
rect 11440 16612 13728 16640
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 14090 16640 14096 16652
rect 13832 16612 14096 16640
rect 11164 16544 11652 16572
rect 9125 16507 9183 16513
rect 9125 16504 9137 16507
rect 8772 16476 9137 16504
rect 9125 16473 9137 16476
rect 9171 16473 9183 16507
rect 9125 16467 9183 16473
rect 9214 16464 9220 16516
rect 9272 16504 9278 16516
rect 11624 16504 11652 16544
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11756 16544 11989 16572
rect 11756 16532 11762 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13832 16572 13860 16612
rect 14090 16600 14096 16612
rect 14148 16600 14154 16652
rect 14274 16600 14280 16652
rect 14332 16600 14338 16652
rect 14384 16640 14412 16680
rect 16022 16668 16028 16720
rect 16080 16668 16086 16720
rect 16114 16668 16120 16720
rect 16172 16708 16178 16720
rect 16298 16708 16304 16720
rect 16172 16680 16304 16708
rect 16172 16668 16178 16680
rect 16298 16668 16304 16680
rect 16356 16668 16362 16720
rect 21542 16668 21548 16720
rect 21600 16708 21606 16720
rect 22186 16708 22192 16720
rect 21600 16680 22192 16708
rect 21600 16668 21606 16680
rect 22186 16668 22192 16680
rect 22244 16668 22250 16720
rect 23658 16708 23664 16720
rect 23584 16680 23664 16708
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 14384 16612 14565 16640
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 16850 16600 16856 16652
rect 16908 16640 16914 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 16908 16612 17141 16640
rect 16908 16600 16914 16612
rect 17129 16609 17141 16612
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 17862 16640 17868 16652
rect 17451 16612 17868 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 18414 16600 18420 16652
rect 18472 16640 18478 16652
rect 18782 16640 18788 16652
rect 18472 16612 18788 16640
rect 18472 16600 18478 16612
rect 18782 16600 18788 16612
rect 18840 16600 18846 16652
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 22278 16640 22284 16652
rect 19475 16612 22284 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16640 22615 16643
rect 23584 16640 23612 16680
rect 23658 16668 23664 16680
rect 23716 16668 23722 16720
rect 22603 16612 23612 16640
rect 22603 16609 22615 16612
rect 22557 16603 22615 16609
rect 24762 16600 24768 16652
rect 24820 16640 24826 16652
rect 25682 16640 25688 16652
rect 24820 16612 25688 16640
rect 24820 16600 24826 16612
rect 25682 16600 25688 16612
rect 25740 16600 25746 16652
rect 13412 16544 13860 16572
rect 16669 16575 16727 16581
rect 13412 16532 13418 16544
rect 16669 16541 16681 16575
rect 16715 16572 16727 16575
rect 16942 16572 16948 16584
rect 16715 16544 16948 16572
rect 16715 16541 16727 16544
rect 16669 16535 16727 16541
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 21821 16575 21879 16581
rect 21821 16541 21833 16575
rect 21867 16572 21879 16575
rect 22002 16572 22008 16584
rect 21867 16544 22008 16572
rect 21867 16541 21879 16544
rect 21821 16535 21879 16541
rect 22002 16532 22008 16544
rect 22060 16532 22066 16584
rect 23934 16532 23940 16584
rect 23992 16572 23998 16584
rect 24581 16575 24639 16581
rect 24581 16572 24593 16575
rect 23992 16544 24593 16572
rect 23992 16532 23998 16544
rect 24581 16541 24593 16544
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 11882 16504 11888 16516
rect 9272 16476 9444 16504
rect 11624 16476 11888 16504
rect 9272 16464 9278 16476
rect 2464 16408 2774 16436
rect 3421 16439 3479 16445
rect 2464 16396 2470 16408
rect 3421 16405 3433 16439
rect 3467 16436 3479 16439
rect 4890 16436 4896 16448
rect 3467 16408 4896 16436
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 4890 16396 4896 16408
rect 4948 16396 4954 16448
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 5077 16439 5135 16445
rect 5077 16436 5089 16439
rect 5040 16408 5089 16436
rect 5040 16396 5046 16408
rect 5077 16405 5089 16408
rect 5123 16405 5135 16439
rect 5077 16399 5135 16405
rect 7469 16439 7527 16445
rect 7469 16405 7481 16439
rect 7515 16436 7527 16439
rect 8294 16436 8300 16448
rect 7515 16408 8300 16436
rect 7515 16405 7527 16408
rect 7469 16399 7527 16405
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 8570 16396 8576 16448
rect 8628 16396 8634 16448
rect 9416 16445 9444 16476
rect 11882 16464 11888 16476
rect 11940 16464 11946 16516
rect 12250 16464 12256 16516
rect 12308 16464 12314 16516
rect 15838 16504 15844 16516
rect 15778 16476 15844 16504
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 17678 16504 17684 16516
rect 15948 16476 17684 16504
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16436 9459 16439
rect 9490 16436 9496 16448
rect 9447 16408 9496 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 10321 16439 10379 16445
rect 10321 16405 10333 16439
rect 10367 16436 10379 16439
rect 10502 16436 10508 16448
rect 10367 16408 10508 16436
rect 10367 16405 10379 16408
rect 10321 16399 10379 16405
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 10594 16396 10600 16448
rect 10652 16436 10658 16448
rect 10781 16439 10839 16445
rect 10781 16436 10793 16439
rect 10652 16408 10793 16436
rect 10652 16396 10658 16408
rect 10781 16405 10793 16408
rect 10827 16405 10839 16439
rect 10781 16399 10839 16405
rect 11146 16396 11152 16448
rect 11204 16396 11210 16448
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 12216 16408 13737 16436
rect 12216 16396 12222 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 14642 16396 14648 16448
rect 14700 16436 14706 16448
rect 15948 16436 15976 16476
rect 17678 16464 17684 16476
rect 17736 16464 17742 16516
rect 18630 16476 19656 16504
rect 14700 16408 15976 16436
rect 16485 16439 16543 16445
rect 14700 16396 14706 16408
rect 16485 16405 16497 16439
rect 16531 16436 16543 16439
rect 18782 16436 18788 16448
rect 16531 16408 18788 16436
rect 16531 16405 16543 16408
rect 16485 16399 16543 16405
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 18874 16396 18880 16448
rect 18932 16396 18938 16448
rect 19628 16436 19656 16476
rect 19702 16464 19708 16516
rect 19760 16464 19766 16516
rect 23842 16504 23848 16516
rect 20088 16476 20194 16504
rect 23782 16476 23848 16504
rect 19794 16436 19800 16448
rect 19628 16408 19800 16436
rect 19794 16396 19800 16408
rect 19852 16436 19858 16448
rect 20088 16436 20116 16476
rect 23842 16464 23848 16476
rect 23900 16464 23906 16516
rect 19852 16408 20116 16436
rect 19852 16396 19858 16408
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 21048 16408 21189 16436
rect 21048 16396 21054 16408
rect 21177 16405 21189 16408
rect 21223 16405 21235 16439
rect 21177 16399 21235 16405
rect 21637 16439 21695 16445
rect 21637 16405 21649 16439
rect 21683 16436 21695 16439
rect 21726 16436 21732 16448
rect 21683 16408 21732 16436
rect 21683 16405 21695 16408
rect 21637 16399 21695 16405
rect 21726 16396 21732 16408
rect 21784 16396 21790 16448
rect 22186 16396 22192 16448
rect 22244 16436 22250 16448
rect 22738 16436 22744 16448
rect 22244 16408 22744 16436
rect 22244 16396 22250 16408
rect 22738 16396 22744 16408
rect 22796 16396 22802 16448
rect 24026 16396 24032 16448
rect 24084 16396 24090 16448
rect 24210 16396 24216 16448
rect 24268 16436 24274 16448
rect 25225 16439 25283 16445
rect 25225 16436 25237 16439
rect 24268 16408 25237 16436
rect 24268 16396 24274 16408
rect 25225 16405 25237 16408
rect 25271 16405 25283 16439
rect 25225 16399 25283 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 1578 16192 1584 16244
rect 1636 16192 1642 16244
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4893 16235 4951 16241
rect 4893 16232 4905 16235
rect 4304 16204 4905 16232
rect 4304 16192 4310 16204
rect 4893 16201 4905 16204
rect 4939 16201 4951 16235
rect 4893 16195 4951 16201
rect 5258 16192 5264 16244
rect 5316 16232 5322 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5316 16204 6009 16232
rect 5316 16192 5322 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 6546 16192 6552 16244
rect 6604 16192 6610 16244
rect 7837 16235 7895 16241
rect 7837 16232 7849 16235
rect 6840 16204 7849 16232
rect 1596 16096 1624 16192
rect 2682 16124 2688 16176
rect 2740 16164 2746 16176
rect 5166 16164 5172 16176
rect 2740 16136 5172 16164
rect 2740 16124 2746 16136
rect 5166 16124 5172 16136
rect 5224 16124 5230 16176
rect 5718 16124 5724 16176
rect 5776 16164 5782 16176
rect 6840 16164 6868 16204
rect 7837 16201 7849 16204
rect 7883 16201 7895 16235
rect 7837 16195 7895 16201
rect 7926 16192 7932 16244
rect 7984 16232 7990 16244
rect 8662 16232 8668 16244
rect 7984 16204 8668 16232
rect 7984 16192 7990 16204
rect 8662 16192 8668 16204
rect 8720 16192 8726 16244
rect 8938 16192 8944 16244
rect 8996 16232 9002 16244
rect 10594 16232 10600 16244
rect 8996 16204 10600 16232
rect 8996 16192 9002 16204
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 11149 16235 11207 16241
rect 11149 16201 11161 16235
rect 11195 16232 11207 16235
rect 12250 16232 12256 16244
rect 11195 16204 12256 16232
rect 11195 16201 11207 16204
rect 11149 16195 11207 16201
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 13446 16192 13452 16244
rect 13504 16192 13510 16244
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 15381 16235 15439 16241
rect 15381 16232 15393 16235
rect 13780 16204 15393 16232
rect 13780 16192 13786 16204
rect 15381 16201 15393 16204
rect 15427 16201 15439 16235
rect 15381 16195 15439 16201
rect 18322 16192 18328 16244
rect 18380 16192 18386 16244
rect 18782 16192 18788 16244
rect 18840 16232 18846 16244
rect 19613 16235 19671 16241
rect 19613 16232 19625 16235
rect 18840 16204 19625 16232
rect 18840 16192 18846 16204
rect 19613 16201 19625 16204
rect 19659 16201 19671 16235
rect 19613 16195 19671 16201
rect 20254 16192 20260 16244
rect 20312 16232 20318 16244
rect 20806 16232 20812 16244
rect 20312 16204 20812 16232
rect 20312 16192 20318 16204
rect 20806 16192 20812 16204
rect 20864 16232 20870 16244
rect 21174 16232 21180 16244
rect 20864 16204 21180 16232
rect 20864 16192 20870 16204
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 21450 16192 21456 16244
rect 21508 16232 21514 16244
rect 21726 16232 21732 16244
rect 21508 16204 21732 16232
rect 21508 16192 21514 16204
rect 21726 16192 21732 16204
rect 21784 16192 21790 16244
rect 22296 16204 23152 16232
rect 10962 16164 10968 16176
rect 5776 16136 6868 16164
rect 7208 16136 10968 16164
rect 5776 16124 5782 16136
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 1596 16068 2053 16096
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 2041 16059 2099 16065
rect 2746 16068 3157 16096
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 16028 1823 16031
rect 2746 16028 2774 16068
rect 3145 16065 3157 16068
rect 3191 16096 3203 16099
rect 3326 16096 3332 16108
rect 3191 16068 3332 16096
rect 3191 16065 3203 16068
rect 3145 16059 3203 16065
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16065 4307 16099
rect 4249 16059 4307 16065
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16096 5411 16099
rect 6454 16096 6460 16108
rect 5399 16068 6460 16096
rect 5399 16065 5411 16068
rect 5353 16059 5411 16065
rect 1811 16000 2774 16028
rect 4264 16028 4292 16059
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 6730 16056 6736 16108
rect 6788 16056 6794 16108
rect 6822 16056 6828 16108
rect 6880 16096 6886 16108
rect 7208 16105 7236 16136
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 11882 16124 11888 16176
rect 11940 16164 11946 16176
rect 11940 16136 12466 16164
rect 11940 16124 11946 16136
rect 13354 16124 13360 16176
rect 13412 16164 13418 16176
rect 13906 16164 13912 16176
rect 13412 16136 13912 16164
rect 13412 16124 13418 16136
rect 13906 16124 13912 16136
rect 13964 16124 13970 16176
rect 14826 16124 14832 16176
rect 14884 16164 14890 16176
rect 15013 16167 15071 16173
rect 15013 16164 15025 16167
rect 14884 16136 15025 16164
rect 14884 16124 14890 16136
rect 15013 16133 15025 16136
rect 15059 16164 15071 16167
rect 15841 16167 15899 16173
rect 15841 16164 15853 16167
rect 15059 16136 15853 16164
rect 15059 16133 15071 16136
rect 15013 16127 15071 16133
rect 15841 16133 15853 16136
rect 15887 16133 15899 16167
rect 16298 16164 16304 16176
rect 15841 16127 15899 16133
rect 15948 16136 16304 16164
rect 7193 16099 7251 16105
rect 6880 16068 7144 16096
rect 6880 16056 6886 16068
rect 7006 16028 7012 16040
rect 4264 16000 7012 16028
rect 1811 15997 1823 16000
rect 1765 15991 1823 15997
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7116 16028 7144 16068
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 8294 16056 8300 16108
rect 8352 16056 8358 16108
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16096 8999 16099
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 8987 16068 9413 16096
rect 8987 16065 8999 16068
rect 8941 16059 8999 16065
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 10134 16096 10140 16108
rect 9732 16068 10140 16096
rect 9732 16056 9738 16068
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 10502 16056 10508 16108
rect 10560 16056 10566 16108
rect 11698 16056 11704 16108
rect 11756 16056 11762 16108
rect 13538 16056 13544 16108
rect 13596 16096 13602 16108
rect 13814 16096 13820 16108
rect 13596 16068 13820 16096
rect 13596 16056 13602 16068
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16096 14335 16099
rect 14918 16096 14924 16108
rect 14323 16068 14924 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 14918 16056 14924 16068
rect 14976 16056 14982 16108
rect 15746 16056 15752 16108
rect 15804 16056 15810 16108
rect 15948 16096 15976 16136
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 18414 16124 18420 16176
rect 18472 16164 18478 16176
rect 19518 16164 19524 16176
rect 18472 16136 19524 16164
rect 18472 16124 18478 16136
rect 19518 16124 19524 16136
rect 19576 16124 19582 16176
rect 19702 16124 19708 16176
rect 19760 16164 19766 16176
rect 22296 16164 22324 16204
rect 19760 16136 22324 16164
rect 22373 16167 22431 16173
rect 19760 16124 19766 16136
rect 22373 16133 22385 16167
rect 22419 16164 22431 16167
rect 22554 16164 22560 16176
rect 22419 16136 22560 16164
rect 22419 16133 22431 16136
rect 22373 16127 22431 16133
rect 22554 16124 22560 16136
rect 22612 16164 22618 16176
rect 23017 16167 23075 16173
rect 23017 16164 23029 16167
rect 22612 16136 23029 16164
rect 22612 16124 22618 16136
rect 23017 16133 23029 16136
rect 23063 16133 23075 16167
rect 23124 16164 23152 16204
rect 23474 16192 23480 16244
rect 23532 16232 23538 16244
rect 23845 16235 23903 16241
rect 23845 16232 23857 16235
rect 23532 16204 23857 16232
rect 23532 16192 23538 16204
rect 23845 16201 23857 16204
rect 23891 16201 23903 16235
rect 23845 16195 23903 16201
rect 25682 16164 25688 16176
rect 23124 16136 25688 16164
rect 23017 16127 23075 16133
rect 25682 16124 25688 16136
rect 25740 16124 25746 16176
rect 15856 16068 15976 16096
rect 17037 16099 17095 16105
rect 9490 16028 9496 16040
rect 7116 16000 9496 16028
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 11146 15988 11152 16040
rect 11204 16028 11210 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 11204 16000 11989 16028
rect 11204 15988 11210 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 14090 16028 14096 16040
rect 12400 16000 14096 16028
rect 12400 15988 12406 16000
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 14369 16031 14427 16037
rect 14369 15997 14381 16031
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 15102 16028 15108 16040
rect 14599 16000 15108 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 2685 15963 2743 15969
rect 2685 15929 2697 15963
rect 2731 15960 2743 15963
rect 5626 15960 5632 15972
rect 2731 15932 5632 15960
rect 2731 15929 2743 15932
rect 2685 15923 2743 15929
rect 5626 15920 5632 15932
rect 5684 15920 5690 15972
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 7190 15960 7196 15972
rect 6788 15932 7196 15960
rect 6788 15920 6794 15932
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 8754 15920 8760 15972
rect 8812 15960 8818 15972
rect 14384 15960 14412 15991
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 15856 15960 15884 16068
rect 17037 16065 17049 16099
rect 17083 16096 17095 16099
rect 19058 16096 19064 16108
rect 17083 16068 19064 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 19168 16068 20269 16096
rect 15930 15988 15936 16040
rect 15988 15988 15994 16040
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 19168 16028 19196 16068
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 16448 16000 19196 16028
rect 16448 15988 16454 16000
rect 19610 15988 19616 16040
rect 19668 16028 19674 16040
rect 19705 16031 19763 16037
rect 19705 16028 19717 16031
rect 19668 16000 19717 16028
rect 19668 15988 19674 16000
rect 19705 15997 19717 16000
rect 19751 15997 19763 16031
rect 19705 15991 19763 15997
rect 19797 16031 19855 16037
rect 19797 15997 19809 16031
rect 19843 15997 19855 16031
rect 20272 16028 20300 16059
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 21453 16099 21511 16105
rect 21453 16096 21465 16099
rect 20864 16068 21465 16096
rect 20864 16056 20870 16068
rect 21453 16065 21465 16068
rect 21499 16065 21511 16099
rect 21453 16059 21511 16065
rect 22465 16099 22523 16105
rect 22465 16065 22477 16099
rect 22511 16096 22523 16099
rect 22738 16096 22744 16108
rect 22511 16068 22744 16096
rect 22511 16065 22523 16068
rect 22465 16059 22523 16065
rect 22738 16056 22744 16068
rect 22796 16056 22802 16108
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16096 23811 16099
rect 24118 16096 24124 16108
rect 23799 16068 24124 16096
rect 23799 16065 23811 16068
rect 23753 16059 23811 16065
rect 24118 16056 24124 16068
rect 24176 16056 24182 16108
rect 24578 16056 24584 16108
rect 24636 16056 24642 16108
rect 20901 16031 20959 16037
rect 20901 16028 20913 16031
rect 20272 16000 20913 16028
rect 19797 15991 19855 15997
rect 20901 15997 20913 16000
rect 20947 15997 20959 16031
rect 20901 15991 20959 15997
rect 8812 15932 11836 15960
rect 8812 15920 8818 15932
rect 3789 15895 3847 15901
rect 3789 15861 3801 15895
rect 3835 15892 3847 15895
rect 3878 15892 3884 15904
rect 3835 15864 3884 15892
rect 3835 15861 3847 15864
rect 3789 15855 3847 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 4890 15852 4896 15904
rect 4948 15892 4954 15904
rect 7466 15892 7472 15904
rect 4948 15864 7472 15892
rect 4948 15852 4954 15864
rect 7466 15852 7472 15864
rect 7524 15852 7530 15904
rect 7926 15852 7932 15904
rect 7984 15892 7990 15904
rect 9950 15892 9956 15904
rect 7984 15864 9956 15892
rect 7984 15852 7990 15864
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10045 15895 10103 15901
rect 10045 15861 10057 15895
rect 10091 15892 10103 15895
rect 10410 15892 10416 15904
rect 10091 15864 10416 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 11808 15892 11836 15932
rect 13832 15932 14320 15960
rect 14384 15932 15884 15960
rect 13832 15892 13860 15932
rect 11808 15864 13860 15892
rect 13906 15852 13912 15904
rect 13964 15852 13970 15904
rect 14292 15892 14320 15932
rect 16298 15920 16304 15972
rect 16356 15960 16362 15972
rect 19245 15963 19303 15969
rect 19245 15960 19257 15963
rect 16356 15932 19257 15960
rect 16356 15920 16362 15932
rect 19245 15929 19257 15932
rect 19291 15929 19303 15963
rect 19245 15923 19303 15929
rect 16393 15895 16451 15901
rect 16393 15892 16405 15895
rect 14292 15864 16405 15892
rect 16393 15861 16405 15864
rect 16439 15892 16451 15895
rect 16482 15892 16488 15904
rect 16439 15864 16488 15892
rect 16439 15861 16451 15864
rect 16393 15855 16451 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 16761 15895 16819 15901
rect 16761 15861 16773 15895
rect 16807 15892 16819 15895
rect 16942 15892 16948 15904
rect 16807 15864 16948 15892
rect 16807 15861 16819 15864
rect 16761 15855 16819 15861
rect 16942 15852 16948 15864
rect 17000 15852 17006 15904
rect 17034 15852 17040 15904
rect 17092 15892 17098 15904
rect 19812 15892 19840 15991
rect 21082 15988 21088 16040
rect 21140 15988 21146 16040
rect 21174 15988 21180 16040
rect 21232 16028 21238 16040
rect 21910 16028 21916 16040
rect 21232 16000 21916 16028
rect 21232 15988 21238 16000
rect 21910 15988 21916 16000
rect 21968 16028 21974 16040
rect 22557 16031 22615 16037
rect 21968 16000 22324 16028
rect 21968 15988 21974 16000
rect 20441 15963 20499 15969
rect 20441 15929 20453 15963
rect 20487 15960 20499 15963
rect 22296 15960 22324 16000
rect 22557 15997 22569 16031
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 22572 15960 22600 15991
rect 24026 15988 24032 16040
rect 24084 16028 24090 16040
rect 24302 16028 24308 16040
rect 24084 16000 24308 16028
rect 24084 15988 24090 16000
rect 24302 15988 24308 16000
rect 24360 15988 24366 16040
rect 23658 15960 23664 15972
rect 20487 15932 22232 15960
rect 22296 15932 22600 15960
rect 22664 15932 23664 15960
rect 20487 15929 20499 15932
rect 20441 15923 20499 15929
rect 17092 15864 19840 15892
rect 17092 15852 17098 15864
rect 22002 15852 22008 15904
rect 22060 15852 22066 15904
rect 22204 15892 22232 15932
rect 22664 15892 22692 15932
rect 23658 15920 23664 15932
rect 23716 15920 23722 15972
rect 22204 15864 22692 15892
rect 23382 15852 23388 15904
rect 23440 15852 23446 15904
rect 25222 15852 25228 15904
rect 25280 15852 25286 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 3973 15691 4031 15697
rect 3973 15657 3985 15691
rect 4019 15688 4031 15691
rect 4154 15688 4160 15700
rect 4019 15660 4160 15688
rect 4019 15657 4031 15660
rect 3973 15651 4031 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 6365 15691 6423 15697
rect 6365 15657 6377 15691
rect 6411 15688 6423 15691
rect 7558 15688 7564 15700
rect 6411 15660 7564 15688
rect 6411 15657 6423 15660
rect 6365 15651 6423 15657
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 10410 15648 10416 15700
rect 10468 15688 10474 15700
rect 10578 15691 10636 15697
rect 10578 15688 10590 15691
rect 10468 15660 10590 15688
rect 10468 15648 10474 15660
rect 10578 15657 10590 15660
rect 10624 15657 10636 15691
rect 13722 15688 13728 15700
rect 10578 15651 10636 15657
rect 13556 15660 13728 15688
rect 2130 15580 2136 15632
rect 2188 15580 2194 15632
rect 2590 15580 2596 15632
rect 2648 15580 2654 15632
rect 7190 15580 7196 15632
rect 7248 15620 7254 15632
rect 9674 15620 9680 15632
rect 7248 15592 9680 15620
rect 7248 15580 7254 15592
rect 9674 15580 9680 15592
rect 9732 15580 9738 15632
rect 11698 15580 11704 15632
rect 11756 15580 11762 15632
rect 12250 15580 12256 15632
rect 12308 15620 12314 15632
rect 12710 15620 12716 15632
rect 12308 15592 12716 15620
rect 12308 15580 12314 15592
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 13556 15620 13584 15660
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 13814 15648 13820 15700
rect 13872 15648 13878 15700
rect 14550 15688 14556 15700
rect 13924 15660 14556 15688
rect 12820 15592 13584 15620
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15552 1639 15555
rect 2608 15552 2636 15580
rect 1627 15524 4200 15552
rect 1627 15521 1639 15524
rect 1581 15515 1639 15521
rect 2590 15444 2596 15496
rect 2648 15444 2654 15496
rect 4172 15493 4200 15524
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 7742 15552 7748 15564
rect 4304 15524 7748 15552
rect 4304 15512 4310 15524
rect 7742 15512 7748 15524
rect 7800 15512 7806 15564
rect 9122 15552 9128 15564
rect 8496 15524 9128 15552
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 1486 15376 1492 15428
rect 1544 15416 1550 15428
rect 1949 15419 2007 15425
rect 1949 15416 1961 15419
rect 1544 15388 1961 15416
rect 1544 15376 1550 15388
rect 1949 15385 1961 15388
rect 1995 15385 2007 15419
rect 2884 15416 2912 15447
rect 4614 15444 4620 15496
rect 4672 15444 4678 15496
rect 5718 15444 5724 15496
rect 5776 15444 5782 15496
rect 5994 15444 6000 15496
rect 6052 15484 6058 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6052 15456 6837 15484
rect 6052 15444 6058 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8496 15484 8524 15524
rect 9122 15512 9128 15524
rect 9180 15552 9186 15564
rect 10321 15555 10379 15561
rect 9180 15524 9996 15552
rect 9180 15512 9186 15524
rect 7975 15456 8524 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 9217 15487 9275 15493
rect 9217 15484 9229 15487
rect 8628 15456 9229 15484
rect 8628 15444 8634 15456
rect 9217 15453 9229 15456
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 4706 15416 4712 15428
rect 2884 15388 4712 15416
rect 1949 15379 2007 15385
rect 4706 15376 4712 15388
rect 4764 15376 4770 15428
rect 7469 15419 7527 15425
rect 7469 15385 7481 15419
rect 7515 15416 7527 15419
rect 8662 15416 8668 15428
rect 7515 15388 8668 15416
rect 7515 15385 7527 15388
rect 7469 15379 7527 15385
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 9968 15416 9996 15524
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 10594 15552 10600 15564
rect 10367 15524 10600 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 10594 15512 10600 15524
rect 10652 15552 10658 15564
rect 11716 15552 11744 15580
rect 10652 15524 11744 15552
rect 10652 15512 10658 15524
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12820 15484 12848 15592
rect 13630 15580 13636 15632
rect 13688 15620 13694 15632
rect 13924 15620 13952 15660
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 14734 15648 14740 15700
rect 14792 15688 14798 15700
rect 16025 15691 16083 15697
rect 16025 15688 16037 15691
rect 14792 15660 16037 15688
rect 14792 15648 14798 15660
rect 16025 15657 16037 15660
rect 16071 15657 16083 15691
rect 16025 15651 16083 15657
rect 16574 15648 16580 15700
rect 16632 15648 16638 15700
rect 17586 15688 17592 15700
rect 17052 15660 17592 15688
rect 13688 15592 13952 15620
rect 13688 15580 13694 15592
rect 16482 15580 16488 15632
rect 16540 15620 16546 15632
rect 17052 15620 17080 15660
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 18693 15691 18751 15697
rect 18693 15657 18705 15691
rect 18739 15688 18751 15691
rect 20898 15688 20904 15700
rect 18739 15660 20904 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 20898 15648 20904 15660
rect 20956 15688 20962 15700
rect 21450 15688 21456 15700
rect 20956 15660 21456 15688
rect 20956 15648 20962 15660
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 22370 15648 22376 15700
rect 22428 15688 22434 15700
rect 23014 15688 23020 15700
rect 22428 15660 23020 15688
rect 22428 15648 22434 15660
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 23753 15691 23811 15697
rect 23753 15657 23765 15691
rect 23799 15688 23811 15691
rect 24578 15688 24584 15700
rect 23799 15660 24584 15688
rect 23799 15657 23811 15660
rect 23753 15651 23811 15657
rect 24578 15648 24584 15660
rect 24636 15648 24642 15700
rect 16540 15592 17080 15620
rect 16540 15580 16546 15592
rect 18874 15580 18880 15632
rect 18932 15620 18938 15632
rect 23934 15620 23940 15632
rect 18932 15592 23940 15620
rect 18932 15580 18938 15592
rect 13173 15555 13231 15561
rect 13173 15521 13185 15555
rect 13219 15552 13231 15555
rect 13814 15552 13820 15564
rect 13219 15524 13820 15552
rect 13219 15521 13231 15524
rect 13173 15515 13231 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 14274 15512 14280 15564
rect 14332 15552 14338 15564
rect 14332 15524 16988 15552
rect 14332 15512 14338 15524
rect 16960 15496 16988 15524
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 19337 15555 19395 15561
rect 19337 15521 19349 15555
rect 19383 15552 19395 15555
rect 19610 15552 19616 15564
rect 19383 15524 19616 15552
rect 19383 15521 19395 15524
rect 19337 15515 19395 15521
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 19978 15512 19984 15564
rect 20036 15512 20042 15564
rect 20070 15512 20076 15564
rect 20128 15512 20134 15564
rect 20180 15561 20208 15592
rect 23934 15580 23940 15592
rect 23992 15580 23998 15632
rect 20165 15555 20223 15561
rect 20165 15521 20177 15555
rect 20211 15521 20223 15555
rect 20165 15515 20223 15521
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 21361 15555 21419 15561
rect 21361 15521 21373 15555
rect 21407 15521 21419 15555
rect 21361 15515 21419 15521
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 12216 15456 12848 15484
rect 12912 15456 13737 15484
rect 12216 15444 12222 15456
rect 11882 15416 11888 15428
rect 9968 15388 10640 15416
rect 11822 15388 11888 15416
rect 4430 15308 4436 15360
rect 4488 15348 4494 15360
rect 4890 15348 4896 15360
rect 4488 15320 4896 15348
rect 4488 15308 4494 15320
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 5258 15308 5264 15360
rect 5316 15308 5322 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 7926 15348 7932 15360
rect 7616 15320 7932 15348
rect 7616 15308 7622 15320
rect 7926 15308 7932 15320
rect 7984 15308 7990 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 8573 15351 8631 15357
rect 8573 15348 8585 15351
rect 8352 15320 8585 15348
rect 8352 15308 8358 15320
rect 8573 15317 8585 15320
rect 8619 15317 8631 15351
rect 8573 15311 8631 15317
rect 9861 15351 9919 15357
rect 9861 15317 9873 15351
rect 9907 15348 9919 15351
rect 10502 15348 10508 15360
rect 9907 15320 10508 15348
rect 9907 15317 9919 15320
rect 9861 15311 9919 15317
rect 10502 15308 10508 15320
rect 10560 15308 10566 15360
rect 10612 15348 10640 15388
rect 11882 15376 11888 15388
rect 11940 15376 11946 15428
rect 11974 15376 11980 15428
rect 12032 15416 12038 15428
rect 12912 15416 12940 15456
rect 13725 15453 13737 15456
rect 13771 15484 13783 15487
rect 14090 15484 14096 15496
rect 13771 15456 14096 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 16298 15484 16304 15496
rect 15686 15456 16304 15484
rect 16298 15444 16304 15456
rect 16356 15484 16362 15496
rect 16356 15456 16896 15484
rect 16356 15444 16362 15456
rect 12032 15388 12940 15416
rect 12989 15419 13047 15425
rect 12032 15376 12038 15388
rect 12989 15385 13001 15419
rect 13035 15416 13047 15419
rect 13035 15388 14504 15416
rect 13035 15385 13047 15388
rect 12989 15379 13047 15385
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 10612 15320 12081 15348
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12069 15311 12127 15317
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 12529 15351 12587 15357
rect 12529 15348 12541 15351
rect 12492 15320 12541 15348
rect 12492 15308 12498 15320
rect 12529 15317 12541 15320
rect 12575 15317 12587 15351
rect 12529 15311 12587 15317
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 12768 15320 12909 15348
rect 12768 15308 12774 15320
rect 12897 15317 12909 15320
rect 12943 15317 12955 15351
rect 12897 15311 12955 15317
rect 13722 15308 13728 15360
rect 13780 15348 13786 15360
rect 14366 15348 14372 15360
rect 13780 15320 14372 15348
rect 13780 15308 13786 15320
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 14476 15348 14504 15388
rect 14550 15376 14556 15428
rect 14608 15376 14614 15428
rect 16666 15416 16672 15428
rect 15856 15388 16672 15416
rect 15856 15348 15884 15388
rect 16666 15376 16672 15388
rect 16724 15376 16730 15428
rect 16868 15416 16896 15456
rect 16942 15444 16948 15496
rect 17000 15444 17006 15496
rect 19996 15484 20024 15512
rect 18984 15456 20024 15484
rect 20717 15487 20775 15493
rect 17678 15416 17684 15428
rect 16868 15388 17684 15416
rect 14476 15320 15884 15348
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 16172 15320 16313 15348
rect 16172 15308 16178 15320
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 17604 15348 17632 15388
rect 17678 15376 17684 15388
rect 17736 15376 17742 15428
rect 18984 15348 19012 15456
rect 20717 15453 20729 15487
rect 20763 15484 20775 15487
rect 20806 15484 20812 15496
rect 20763 15456 20812 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 20806 15444 20812 15456
rect 20864 15484 20870 15496
rect 21177 15487 21235 15493
rect 21177 15484 21189 15487
rect 20864 15456 21189 15484
rect 20864 15444 20870 15456
rect 21177 15453 21189 15456
rect 21223 15453 21235 15487
rect 21376 15484 21404 15515
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 21508 15524 24624 15552
rect 21508 15512 21514 15524
rect 21177 15447 21235 15453
rect 21284 15456 21404 15484
rect 19426 15376 19432 15428
rect 19484 15416 19490 15428
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 19484 15388 19993 15416
rect 19484 15376 19490 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 20162 15376 20168 15428
rect 20220 15416 20226 15428
rect 20220 15388 20944 15416
rect 20220 15376 20226 15388
rect 17604 15320 19012 15348
rect 16301 15311 16359 15317
rect 19058 15308 19064 15360
rect 19116 15308 19122 15360
rect 19610 15308 19616 15360
rect 19668 15308 19674 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 20809 15351 20867 15357
rect 20809 15348 20821 15351
rect 19852 15320 20821 15348
rect 19852 15308 19858 15320
rect 20809 15317 20821 15320
rect 20855 15317 20867 15351
rect 20916 15348 20944 15388
rect 20990 15376 20996 15428
rect 21048 15416 21054 15428
rect 21284 15416 21312 15456
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22462 15484 22468 15496
rect 22244 15456 22468 15484
rect 22244 15444 22250 15456
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 23109 15487 23167 15493
rect 23109 15453 23121 15487
rect 23155 15484 23167 15487
rect 24210 15484 24216 15496
rect 23155 15456 24216 15484
rect 23155 15453 23167 15456
rect 23109 15447 23167 15453
rect 24210 15444 24216 15456
rect 24268 15444 24274 15496
rect 24596 15493 24624 15524
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 21048 15388 21312 15416
rect 21048 15376 21054 15388
rect 25774 15376 25780 15428
rect 25832 15416 25838 15428
rect 26418 15416 26424 15428
rect 25832 15388 26424 15416
rect 25832 15376 25838 15388
rect 26418 15376 26424 15388
rect 26476 15376 26482 15428
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 20916 15320 22661 15348
rect 20809 15311 20867 15317
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 22649 15311 22707 15317
rect 24118 15308 24124 15360
rect 24176 15308 24182 15360
rect 25225 15351 25283 15357
rect 25225 15317 25237 15351
rect 25271 15348 25283 15351
rect 25498 15348 25504 15360
rect 25271 15320 25504 15348
rect 25271 15317 25283 15320
rect 25225 15311 25283 15317
rect 25498 15308 25504 15320
rect 25556 15308 25562 15360
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 2590 15104 2596 15156
rect 2648 15144 2654 15156
rect 4893 15147 4951 15153
rect 4893 15144 4905 15147
rect 2648 15116 4905 15144
rect 2648 15104 2654 15116
rect 4893 15113 4905 15116
rect 4939 15113 4951 15147
rect 4893 15107 4951 15113
rect 5902 15104 5908 15156
rect 5960 15144 5966 15156
rect 5997 15147 6055 15153
rect 5997 15144 6009 15147
rect 5960 15116 6009 15144
rect 5960 15104 5966 15116
rect 5997 15113 6009 15116
rect 6043 15113 6055 15147
rect 5997 15107 6055 15113
rect 6270 15104 6276 15156
rect 6328 15144 6334 15156
rect 7282 15144 7288 15156
rect 6328 15116 7288 15144
rect 6328 15104 6334 15116
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7708 15116 7849 15144
rect 7708 15104 7714 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 13814 15144 13820 15156
rect 7837 15107 7895 15113
rect 9416 15116 13820 15144
rect 1854 15036 1860 15088
rect 1912 15076 1918 15088
rect 2130 15076 2136 15088
rect 1912 15048 2136 15076
rect 1912 15036 1918 15048
rect 2130 15036 2136 15048
rect 2188 15036 2194 15088
rect 2222 15036 2228 15088
rect 2280 15076 2286 15088
rect 2280 15048 7236 15076
rect 2280 15036 2286 15048
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 15008 3203 15011
rect 4154 15008 4160 15020
rect 3191 14980 4160 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 1946 14940 1952 14952
rect 1903 14912 1952 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 2133 14943 2191 14949
rect 2133 14909 2145 14943
rect 2179 14940 2191 14943
rect 3786 14940 3792 14952
rect 2179 14912 3792 14940
rect 2179 14909 2191 14912
rect 2133 14903 2191 14909
rect 3786 14900 3792 14912
rect 3844 14900 3850 14952
rect 1670 14832 1676 14884
rect 1728 14872 1734 14884
rect 4264 14872 4292 14971
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 5353 15011 5411 15017
rect 5353 15008 5365 15011
rect 4580 14980 5365 15008
rect 4580 14968 4586 14980
rect 5353 14977 5365 14980
rect 5399 15008 5411 15011
rect 5442 15008 5448 15020
rect 5399 14980 5448 15008
rect 5399 14977 5411 14980
rect 5353 14971 5411 14977
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 7208 15017 7236 15048
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 15008 8355 15011
rect 8570 15008 8576 15020
rect 8343 14980 8576 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 6748 14940 6776 14971
rect 8570 14968 8576 14980
rect 8628 14968 8634 15020
rect 9416 15017 9444 15116
rect 13814 15104 13820 15116
rect 13872 15144 13878 15156
rect 14461 15147 14519 15153
rect 14461 15144 14473 15147
rect 13872 15116 14473 15144
rect 13872 15104 13878 15116
rect 14461 15113 14473 15116
rect 14507 15113 14519 15147
rect 14461 15107 14519 15113
rect 15562 15104 15568 15156
rect 15620 15104 15626 15156
rect 17954 15144 17960 15156
rect 15672 15116 17960 15144
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 10870 15076 10876 15088
rect 10008 15048 10876 15076
rect 10008 15036 10014 15048
rect 10870 15036 10876 15048
rect 10928 15036 10934 15088
rect 11146 15036 11152 15088
rect 11204 15036 11210 15088
rect 12158 15036 12164 15088
rect 12216 15036 12222 15088
rect 13262 15076 13268 15088
rect 12728 15048 13268 15076
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 15008 11851 15011
rect 12526 15008 12532 15020
rect 11839 14980 12532 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 12526 14968 12532 14980
rect 12584 15008 12590 15020
rect 12728 15008 12756 15048
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 13446 15036 13452 15088
rect 13504 15036 13510 15088
rect 12584 14980 12756 15008
rect 12584 14968 12590 14980
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 14792 14980 14933 15008
rect 14792 14968 14798 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 9030 14940 9036 14952
rect 6748 14912 9036 14940
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9490 14900 9496 14952
rect 9548 14940 9554 14952
rect 11238 14940 11244 14952
rect 9548 14912 11244 14940
rect 9548 14900 9554 14912
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14940 12771 14943
rect 12989 14943 13047 14949
rect 12759 14912 12848 14940
rect 12759 14909 12771 14912
rect 12713 14903 12771 14909
rect 7742 14872 7748 14884
rect 1728 14844 4292 14872
rect 6472 14844 7748 14872
rect 1728 14832 1734 14844
rect 1854 14764 1860 14816
rect 1912 14804 1918 14816
rect 3510 14804 3516 14816
rect 1912 14776 3516 14804
rect 1912 14764 1918 14776
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 3789 14807 3847 14813
rect 3789 14773 3801 14807
rect 3835 14804 3847 14807
rect 6472 14804 6500 14844
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 9214 14832 9220 14884
rect 9272 14872 9278 14884
rect 12158 14872 12164 14884
rect 9272 14844 12164 14872
rect 9272 14832 9278 14844
rect 12158 14832 12164 14844
rect 12216 14832 12222 14884
rect 3835 14776 6500 14804
rect 6549 14807 6607 14813
rect 3835 14773 3847 14776
rect 3789 14767 3847 14773
rect 6549 14773 6561 14807
rect 6595 14804 6607 14807
rect 7558 14804 7564 14816
rect 6595 14776 7564 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 8941 14807 8999 14813
rect 8941 14773 8953 14807
rect 8987 14804 8999 14807
rect 9674 14804 9680 14816
rect 8987 14776 9680 14804
rect 8987 14773 8999 14776
rect 8941 14767 8999 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 10045 14807 10103 14813
rect 10045 14773 10057 14807
rect 10091 14804 10103 14807
rect 10870 14804 10876 14816
rect 10091 14776 10876 14804
rect 10091 14773 10103 14776
rect 10045 14767 10103 14773
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 12820 14804 12848 14912
rect 12989 14909 13001 14943
rect 13035 14940 13047 14943
rect 14826 14940 14832 14952
rect 13035 14912 14832 14940
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 14090 14832 14096 14884
rect 14148 14872 14154 14884
rect 15672 14872 15700 15116
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 25130 15144 25136 15156
rect 19628 15116 25136 15144
rect 16114 15036 16120 15088
rect 16172 15036 16178 15088
rect 17034 15076 17040 15088
rect 16224 15048 17040 15076
rect 14148 14844 15700 14872
rect 14148 14832 14154 14844
rect 14274 14804 14280 14816
rect 12820 14776 14280 14804
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 16224 14804 16252 15048
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 17678 15036 17684 15088
rect 17736 15036 17742 15088
rect 19628 15085 19656 15116
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 19613 15079 19671 15085
rect 19613 15045 19625 15079
rect 19659 15045 19671 15079
rect 19613 15039 19671 15045
rect 20070 15036 20076 15088
rect 20128 15036 20134 15088
rect 21450 15036 21456 15088
rect 21508 15036 21514 15088
rect 22370 15036 22376 15088
rect 22428 15076 22434 15088
rect 23017 15079 23075 15085
rect 23017 15076 23029 15079
rect 22428 15048 23029 15076
rect 22428 15036 22434 15048
rect 23017 15045 23029 15048
rect 23063 15045 23075 15079
rect 23017 15039 23075 15045
rect 23566 15036 23572 15088
rect 23624 15036 23630 15088
rect 21542 14968 21548 15020
rect 21600 15008 21606 15020
rect 22097 15011 22155 15017
rect 22097 15008 22109 15011
rect 21600 14980 22109 15008
rect 21600 14968 21606 14980
rect 22097 14977 22109 14980
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 22278 14968 22284 15020
rect 22336 15008 22342 15020
rect 22741 15011 22799 15017
rect 22741 15008 22753 15011
rect 22336 14980 22753 15008
rect 22336 14968 22342 14980
rect 22741 14977 22753 14980
rect 22787 14977 22799 15011
rect 22741 14971 22799 14977
rect 25133 15011 25191 15017
rect 25133 14977 25145 15011
rect 25179 15008 25191 15011
rect 25590 15008 25596 15020
rect 25179 14980 25596 15008
rect 25179 14977 25191 14980
rect 25133 14971 25191 14977
rect 25590 14968 25596 14980
rect 25648 14968 25654 15020
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 17218 14940 17224 14952
rect 17175 14912 17224 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 16301 14875 16359 14881
rect 16301 14841 16313 14875
rect 16347 14872 16359 14875
rect 16482 14872 16488 14884
rect 16347 14844 16488 14872
rect 16347 14841 16359 14844
rect 16301 14835 16359 14841
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 16868 14816 16896 14903
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 19334 14940 19340 14952
rect 18156 14912 19340 14940
rect 14792 14776 16252 14804
rect 14792 14764 14798 14776
rect 16574 14764 16580 14816
rect 16632 14804 16638 14816
rect 16850 14804 16856 14816
rect 16632 14776 16856 14804
rect 16632 14764 16638 14776
rect 16850 14764 16856 14776
rect 16908 14804 16914 14816
rect 18156 14804 18184 14912
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 22646 14940 22652 14952
rect 19444 14912 22652 14940
rect 18874 14832 18880 14884
rect 18932 14872 18938 14884
rect 19061 14875 19119 14881
rect 19061 14872 19073 14875
rect 18932 14844 19073 14872
rect 18932 14832 18938 14844
rect 19061 14841 19073 14844
rect 19107 14872 19119 14875
rect 19444 14872 19472 14912
rect 22646 14900 22652 14912
rect 22704 14900 22710 14952
rect 23382 14940 23388 14952
rect 22756 14912 23388 14940
rect 22756 14884 22784 14912
rect 23382 14900 23388 14912
rect 23440 14900 23446 14952
rect 24394 14900 24400 14952
rect 24452 14940 24458 14952
rect 24489 14943 24547 14949
rect 24489 14940 24501 14943
rect 24452 14912 24501 14940
rect 24452 14900 24458 14912
rect 24489 14909 24501 14912
rect 24535 14909 24547 14943
rect 24489 14903 24547 14909
rect 19107 14844 19472 14872
rect 21085 14875 21143 14881
rect 19107 14841 19119 14844
rect 19061 14835 19119 14841
rect 21085 14841 21097 14875
rect 21131 14872 21143 14875
rect 22281 14875 22339 14881
rect 21131 14844 22094 14872
rect 21131 14841 21143 14844
rect 21085 14835 21143 14841
rect 16908 14776 18184 14804
rect 18601 14807 18659 14813
rect 16908 14764 16914 14776
rect 18601 14773 18613 14807
rect 18647 14804 18659 14807
rect 20714 14804 20720 14816
rect 18647 14776 20720 14804
rect 18647 14773 18659 14776
rect 18601 14767 18659 14773
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 21542 14764 21548 14816
rect 21600 14764 21606 14816
rect 22066 14804 22094 14844
rect 22281 14841 22293 14875
rect 22327 14872 22339 14875
rect 22462 14872 22468 14884
rect 22327 14844 22468 14872
rect 22327 14841 22339 14844
rect 22281 14835 22339 14841
rect 22462 14832 22468 14844
rect 22520 14832 22526 14884
rect 22738 14832 22744 14884
rect 22796 14832 22802 14884
rect 23014 14804 23020 14816
rect 22066 14776 23020 14804
rect 23014 14764 23020 14776
rect 23072 14804 23078 14816
rect 24578 14804 24584 14816
rect 23072 14776 24584 14804
rect 23072 14764 23078 14776
rect 24578 14764 24584 14776
rect 24636 14764 24642 14816
rect 25038 14764 25044 14816
rect 25096 14804 25102 14816
rect 25225 14807 25283 14813
rect 25225 14804 25237 14807
rect 25096 14776 25237 14804
rect 25096 14764 25102 14776
rect 25225 14773 25237 14776
rect 25271 14773 25283 14807
rect 25225 14767 25283 14773
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 3970 14600 3976 14612
rect 2148 14572 3976 14600
rect 1578 14356 1584 14408
rect 1636 14356 1642 14408
rect 2148 14405 2176 14572
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 5776 14572 7481 14600
rect 5776 14560 5782 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 7469 14563 7527 14569
rect 8570 14560 8576 14612
rect 8628 14560 8634 14612
rect 9030 14560 9036 14612
rect 9088 14560 9094 14612
rect 9214 14560 9220 14612
rect 9272 14560 9278 14612
rect 9508 14572 11928 14600
rect 5258 14492 5264 14544
rect 5316 14532 5322 14544
rect 5316 14504 6868 14532
rect 5316 14492 5322 14504
rect 2314 14424 2320 14476
rect 2372 14464 2378 14476
rect 2372 14436 5764 14464
rect 2372 14424 2378 14436
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 2682 14396 2688 14408
rect 2639 14368 2688 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 4062 14396 4068 14408
rect 2915 14368 4068 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4430 14396 4436 14408
rect 4203 14368 4436 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 4614 14356 4620 14408
rect 4672 14356 4678 14408
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 5736 14405 5764 14436
rect 6362 14424 6368 14476
rect 6420 14424 6426 14476
rect 6840 14405 6868 14504
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 8938 14464 8944 14476
rect 7340 14436 8944 14464
rect 7340 14424 7346 14436
rect 8938 14424 8944 14436
rect 8996 14424 9002 14476
rect 5261 14399 5319 14405
rect 5261 14396 5273 14399
rect 5224 14368 5273 14396
rect 5224 14356 5230 14368
rect 5261 14365 5273 14368
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14365 5779 14399
rect 5721 14359 5779 14365
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 8294 14396 8300 14408
rect 7975 14368 8300 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 9508 14405 9536 14572
rect 9674 14492 9680 14544
rect 9732 14532 9738 14544
rect 11900 14532 11928 14572
rect 12158 14560 12164 14612
rect 12216 14600 12222 14612
rect 12216 14572 12480 14600
rect 12216 14560 12222 14572
rect 12342 14532 12348 14544
rect 9732 14504 10732 14532
rect 11900 14504 12348 14532
rect 9732 14492 9738 14504
rect 10594 14424 10600 14476
rect 10652 14424 10658 14476
rect 10704 14464 10732 14504
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 12452 14532 12480 14572
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 12621 14603 12679 14609
rect 12621 14600 12633 14603
rect 12584 14572 12633 14600
rect 12584 14560 12590 14572
rect 12621 14569 12633 14572
rect 12667 14569 12679 14603
rect 12621 14563 12679 14569
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 15746 14600 15752 14612
rect 13596 14572 15752 14600
rect 13596 14560 13602 14572
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 16022 14560 16028 14612
rect 16080 14600 16086 14612
rect 16758 14600 16764 14612
rect 16080 14572 16764 14600
rect 16080 14560 16086 14572
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 17770 14600 17776 14612
rect 17460 14572 17776 14600
rect 17460 14560 17466 14572
rect 17770 14560 17776 14572
rect 17828 14600 17834 14612
rect 18233 14603 18291 14609
rect 18233 14600 18245 14603
rect 17828 14572 18245 14600
rect 17828 14560 17834 14572
rect 18233 14569 18245 14572
rect 18279 14569 18291 14603
rect 18233 14563 18291 14569
rect 18598 14560 18604 14612
rect 18656 14600 18662 14612
rect 18693 14603 18751 14609
rect 18693 14600 18705 14603
rect 18656 14572 18705 14600
rect 18656 14560 18662 14572
rect 18693 14569 18705 14572
rect 18739 14569 18751 14603
rect 18693 14563 18751 14569
rect 21910 14560 21916 14612
rect 21968 14600 21974 14612
rect 22094 14600 22100 14612
rect 21968 14572 22100 14600
rect 21968 14560 21974 14572
rect 22094 14560 22100 14572
rect 22152 14560 22158 14612
rect 22278 14560 22284 14612
rect 22336 14560 22342 14612
rect 12452 14504 14412 14532
rect 10873 14467 10931 14473
rect 10873 14464 10885 14467
rect 10704 14436 10885 14464
rect 10873 14433 10885 14436
rect 10919 14433 10931 14467
rect 10873 14427 10931 14433
rect 10962 14424 10968 14476
rect 11020 14464 11026 14476
rect 14090 14464 14096 14476
rect 11020 14436 14096 14464
rect 11020 14424 11026 14436
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14384 14464 14412 14504
rect 15856 14504 16620 14532
rect 15194 14464 15200 14476
rect 14384 14436 15200 14464
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 12250 14396 12256 14408
rect 11940 14368 12256 14396
rect 11940 14356 11946 14368
rect 12250 14356 12256 14368
rect 12308 14396 12314 14408
rect 13081 14399 13139 14405
rect 12308 14368 13032 14396
rect 12308 14356 12314 14368
rect 1596 14328 1624 14356
rect 2314 14328 2320 14340
rect 1596 14300 2320 14328
rect 2314 14288 2320 14300
rect 2372 14288 2378 14340
rect 3510 14288 3516 14340
rect 3568 14328 3574 14340
rect 5810 14328 5816 14340
rect 3568 14300 5816 14328
rect 3568 14288 3574 14300
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 6546 14288 6552 14340
rect 6604 14328 6610 14340
rect 12710 14328 12716 14340
rect 6604 14300 10272 14328
rect 6604 14288 6610 14300
rect 1578 14220 1584 14272
rect 1636 14260 1642 14272
rect 1949 14263 2007 14269
rect 1949 14260 1961 14263
rect 1636 14232 1961 14260
rect 1636 14220 1642 14232
rect 1949 14229 1961 14232
rect 1995 14229 2007 14263
rect 1949 14223 2007 14229
rect 3970 14220 3976 14272
rect 4028 14220 4034 14272
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 8938 14260 8944 14272
rect 7892 14232 8944 14260
rect 7892 14220 7898 14232
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 10137 14263 10195 14269
rect 10137 14260 10149 14263
rect 9272 14232 10149 14260
rect 9272 14220 9278 14232
rect 10137 14229 10149 14232
rect 10183 14229 10195 14263
rect 10244 14260 10272 14300
rect 12176 14300 12716 14328
rect 12176 14260 12204 14300
rect 12710 14288 12716 14300
rect 12768 14288 12774 14340
rect 13004 14328 13032 14368
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13170 14396 13176 14408
rect 13127 14368 13176 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 13354 14328 13360 14340
rect 13004 14300 13360 14328
rect 13354 14288 13360 14300
rect 13412 14288 13418 14340
rect 13725 14331 13783 14337
rect 13725 14297 13737 14331
rect 13771 14328 13783 14331
rect 14553 14331 14611 14337
rect 14553 14328 14565 14331
rect 13771 14300 14565 14328
rect 13771 14297 13783 14300
rect 13725 14291 13783 14297
rect 14553 14297 14565 14300
rect 14599 14297 14611 14331
rect 14553 14291 14611 14297
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 15010 14328 15016 14340
rect 14700 14300 15016 14328
rect 14700 14288 14706 14300
rect 15010 14288 15016 14300
rect 15068 14288 15074 14340
rect 10244 14232 12204 14260
rect 10137 14223 10195 14229
rect 14090 14220 14096 14272
rect 14148 14260 14154 14272
rect 15856 14260 15884 14504
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 16206 14464 16212 14476
rect 15988 14436 16212 14464
rect 15988 14424 15994 14436
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16485 14467 16543 14473
rect 16485 14433 16497 14467
rect 16531 14433 16543 14467
rect 16592 14464 16620 14504
rect 17862 14492 17868 14544
rect 17920 14532 17926 14544
rect 21450 14532 21456 14544
rect 17920 14504 21456 14532
rect 17920 14492 17926 14504
rect 21450 14492 21456 14504
rect 21508 14492 21514 14544
rect 19794 14464 19800 14476
rect 16592 14436 19800 14464
rect 16485 14427 16543 14433
rect 16500 14328 16528 14427
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 20073 14467 20131 14473
rect 20073 14433 20085 14467
rect 20119 14464 20131 14467
rect 20714 14464 20720 14476
rect 20119 14436 20720 14464
rect 20119 14433 20131 14436
rect 20073 14427 20131 14433
rect 20714 14424 20720 14436
rect 20772 14464 20778 14476
rect 22002 14464 22008 14476
rect 20772 14436 22008 14464
rect 20772 14424 20778 14436
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 23477 14467 23535 14473
rect 23477 14464 23489 14467
rect 23440 14436 23489 14464
rect 23440 14424 23446 14436
rect 23477 14433 23489 14436
rect 23523 14433 23535 14467
rect 23477 14427 23535 14433
rect 23569 14467 23627 14473
rect 23569 14433 23581 14467
rect 23615 14433 23627 14467
rect 23569 14427 23627 14433
rect 18874 14356 18880 14408
rect 18932 14356 18938 14408
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20438 14396 20444 14408
rect 19935 14368 20444 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 22830 14356 22836 14408
rect 22888 14396 22894 14408
rect 23584 14396 23612 14427
rect 24026 14424 24032 14476
rect 24084 14464 24090 14476
rect 25133 14467 25191 14473
rect 25133 14464 25145 14467
rect 24084 14436 25145 14464
rect 24084 14424 24090 14436
rect 25133 14433 25145 14436
rect 25179 14433 25191 14467
rect 25133 14427 25191 14433
rect 22888 14368 23612 14396
rect 25041 14399 25099 14405
rect 22888 14356 22894 14368
rect 25041 14365 25053 14399
rect 25087 14396 25099 14399
rect 25406 14396 25412 14408
rect 25087 14368 25412 14396
rect 25087 14365 25099 14368
rect 25041 14359 25099 14365
rect 25406 14356 25412 14368
rect 25464 14356 25470 14408
rect 16761 14331 16819 14337
rect 16500 14300 16620 14328
rect 16592 14272 16620 14300
rect 16761 14297 16773 14331
rect 16807 14297 16819 14331
rect 16761 14291 16819 14297
rect 14148 14232 15884 14260
rect 14148 14220 14154 14232
rect 16574 14220 16580 14272
rect 16632 14220 16638 14272
rect 16776 14260 16804 14291
rect 17034 14288 17040 14340
rect 17092 14328 17098 14340
rect 17092 14300 17250 14328
rect 17092 14288 17098 14300
rect 18322 14288 18328 14340
rect 18380 14328 18386 14340
rect 20809 14331 20867 14337
rect 20809 14328 20821 14331
rect 18380 14300 20821 14328
rect 18380 14288 18386 14300
rect 20809 14297 20821 14300
rect 20855 14297 20867 14331
rect 24029 14331 24087 14337
rect 24029 14328 24041 14331
rect 20809 14291 20867 14297
rect 23400 14300 24041 14328
rect 23400 14272 23428 14300
rect 24029 14297 24041 14300
rect 24075 14297 24087 14331
rect 24029 14291 24087 14297
rect 24486 14288 24492 14340
rect 24544 14328 24550 14340
rect 25314 14328 25320 14340
rect 24544 14300 25320 14328
rect 24544 14288 24550 14300
rect 25314 14288 25320 14300
rect 25372 14288 25378 14340
rect 17770 14260 17776 14272
rect 16776 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 18472 14232 19441 14260
rect 18472 14220 18478 14232
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19429 14223 19487 14229
rect 19794 14220 19800 14272
rect 19852 14220 19858 14272
rect 20438 14220 20444 14272
rect 20496 14260 20502 14272
rect 21910 14260 21916 14272
rect 20496 14232 21916 14260
rect 20496 14220 20502 14232
rect 21910 14220 21916 14232
rect 21968 14220 21974 14272
rect 23014 14220 23020 14272
rect 23072 14220 23078 14272
rect 23382 14220 23388 14272
rect 23440 14220 23446 14272
rect 24118 14220 24124 14272
rect 24176 14260 24182 14272
rect 24581 14263 24639 14269
rect 24581 14260 24593 14263
rect 24176 14232 24593 14260
rect 24176 14220 24182 14232
rect 24581 14229 24593 14232
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 24762 14220 24768 14272
rect 24820 14260 24826 14272
rect 24949 14263 25007 14269
rect 24949 14260 24961 14263
rect 24820 14232 24961 14260
rect 24820 14220 24826 14232
rect 24949 14229 24961 14232
rect 24995 14229 25007 14263
rect 24949 14223 25007 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 1302 14016 1308 14068
rect 1360 14056 1366 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 1360 14028 2789 14056
rect 1360 14016 1366 14028
rect 2777 14025 2789 14028
rect 2823 14025 2835 14059
rect 2777 14019 2835 14025
rect 2866 14016 2872 14068
rect 2924 14016 2930 14068
rect 4706 14016 4712 14068
rect 4764 14016 4770 14068
rect 6546 14016 6552 14068
rect 6604 14016 6610 14068
rect 8294 14056 8300 14068
rect 6656 14028 8300 14056
rect 3145 13991 3203 13997
rect 3145 13957 3157 13991
rect 3191 13988 3203 13991
rect 4154 13988 4160 14000
rect 3191 13960 4160 13988
rect 3191 13957 3203 13960
rect 3145 13951 3203 13957
rect 4154 13948 4160 13960
rect 4212 13988 4218 14000
rect 6656 13988 6684 14028
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 10594 14056 10600 14068
rect 9508 14028 10600 14056
rect 9122 13988 9128 14000
rect 4212 13960 6684 13988
rect 7208 13960 9128 13988
rect 4212 13948 4218 13960
rect 1578 13880 1584 13932
rect 1636 13880 1642 13932
rect 1854 13880 1860 13932
rect 1912 13880 1918 13932
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13920 3479 13923
rect 3467 13892 4844 13920
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 3694 13812 3700 13864
rect 3752 13812 3758 13864
rect 4816 13852 4844 13892
rect 4890 13880 4896 13932
rect 4948 13880 4954 13932
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 7208 13929 7236 13960
rect 9122 13948 9128 13960
rect 9180 13948 9186 14000
rect 9508 13988 9536 14028
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 11149 14059 11207 14065
rect 11149 14056 11161 14059
rect 11020 14028 11161 14056
rect 11020 14016 11026 14028
rect 11149 14025 11161 14028
rect 11195 14056 11207 14059
rect 11238 14056 11244 14068
rect 11195 14028 11244 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 13170 14016 13176 14068
rect 13228 14016 13234 14068
rect 13722 14056 13728 14068
rect 13556 14028 13728 14056
rect 9416 13960 9536 13988
rect 7193 13923 7251 13929
rect 7193 13889 7205 13923
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13920 8355 13923
rect 9214 13920 9220 13932
rect 8343 13892 9220 13920
rect 8343 13889 8355 13892
rect 8297 13883 8355 13889
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9416 13929 9444 13960
rect 10410 13948 10416 14000
rect 10468 13948 10474 14000
rect 12618 13988 12624 14000
rect 10980 13960 12624 13988
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 5718 13852 5724 13864
rect 4816 13824 5724 13852
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6362 13852 6368 13864
rect 6043 13824 6368 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6362 13812 6368 13824
rect 6420 13812 6426 13864
rect 7834 13812 7840 13864
rect 7892 13812 7898 13864
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13852 8999 13855
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 8987 13824 9689 13852
rect 8987 13821 8999 13824
rect 8941 13815 8999 13821
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 10318 13812 10324 13864
rect 10376 13852 10382 13864
rect 10980 13852 11008 13960
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 11146 13880 11152 13932
rect 11204 13920 11210 13932
rect 11885 13923 11943 13929
rect 11885 13920 11897 13923
rect 11204 13892 11897 13920
rect 11204 13880 11210 13892
rect 11885 13889 11897 13892
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 12069 13923 12127 13929
rect 12069 13889 12081 13923
rect 12115 13920 12127 13923
rect 12342 13920 12348 13932
rect 12115 13892 12348 13920
rect 12115 13889 12127 13892
rect 12069 13883 12127 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 12526 13880 12532 13932
rect 12584 13880 12590 13932
rect 10376 13824 11008 13852
rect 10376 13812 10382 13824
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 13556 13852 13584 14028
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 14274 14016 14280 14068
rect 14332 14016 14338 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 14608 14028 17509 14056
rect 14608 14016 14614 14028
rect 17497 14025 17509 14028
rect 17543 14025 17555 14059
rect 17497 14019 17555 14025
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 18598 14056 18604 14068
rect 17920 14028 18604 14056
rect 17920 14016 17926 14028
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19392 14028 19533 14056
rect 19392 14016 19398 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20346 14016 20352 14068
rect 20404 14016 20410 14068
rect 20717 14059 20775 14065
rect 20717 14025 20729 14059
rect 20763 14056 20775 14059
rect 21818 14056 21824 14068
rect 20763 14028 21824 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 24026 14016 24032 14068
rect 24084 14056 24090 14068
rect 24210 14056 24216 14068
rect 24084 14028 24216 14056
rect 24084 14016 24090 14028
rect 24210 14016 24216 14028
rect 24268 14016 24274 14068
rect 25130 14016 25136 14068
rect 25188 14016 25194 14068
rect 14292 13988 14320 14016
rect 13648 13960 14320 13988
rect 13648 13929 13676 13960
rect 15654 13948 15660 14000
rect 15712 13988 15718 14000
rect 18233 13991 18291 13997
rect 18233 13988 18245 13991
rect 15712 13960 18245 13988
rect 15712 13948 15718 13960
rect 18233 13957 18245 13960
rect 18279 13988 18291 13991
rect 18322 13988 18328 14000
rect 18279 13960 18328 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18322 13948 18328 13960
rect 18380 13948 18386 14000
rect 21177 13991 21235 13997
rect 21177 13957 21189 13991
rect 21223 13988 21235 13991
rect 21358 13988 21364 14000
rect 21223 13960 21364 13988
rect 21223 13957 21235 13960
rect 21177 13951 21235 13957
rect 21358 13948 21364 13960
rect 21416 13948 21422 14000
rect 21910 13948 21916 14000
rect 21968 13988 21974 14000
rect 21968 13960 22324 13988
rect 21968 13948 21974 13960
rect 22296 13932 22324 13960
rect 23566 13948 23572 14000
rect 23624 13948 23630 14000
rect 13633 13923 13691 13929
rect 13633 13889 13645 13923
rect 13679 13889 13691 13923
rect 13633 13883 13691 13889
rect 15010 13880 15016 13932
rect 15068 13920 15074 13932
rect 15841 13923 15899 13929
rect 15068 13892 15516 13920
rect 15068 13880 15074 13892
rect 11480 13824 13584 13852
rect 11480 13812 11486 13824
rect 14550 13812 14556 13864
rect 14608 13852 14614 13864
rect 15102 13852 15108 13864
rect 14608 13824 15108 13852
rect 14608 13812 14614 13824
rect 15102 13812 15108 13824
rect 15160 13852 15166 13864
rect 15381 13855 15439 13861
rect 15381 13852 15393 13855
rect 15160 13824 15393 13852
rect 15160 13812 15166 13824
rect 15381 13821 15393 13824
rect 15427 13821 15439 13855
rect 15488 13852 15516 13892
rect 15841 13889 15853 13923
rect 15887 13920 15899 13923
rect 16298 13920 16304 13932
rect 15887 13892 16304 13920
rect 15887 13889 15899 13892
rect 15841 13883 15899 13889
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 16632 13892 16865 13920
rect 16632 13880 16638 13892
rect 16853 13889 16865 13892
rect 16899 13889 16911 13923
rect 20714 13920 20720 13932
rect 16853 13883 16911 13889
rect 18340 13892 20720 13920
rect 18340 13864 18368 13892
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 22066 13892 22232 13920
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 15488 13824 16037 13852
rect 15381 13815 15439 13821
rect 16025 13821 16037 13824
rect 16071 13852 16083 13855
rect 17034 13852 17040 13864
rect 16071 13824 17040 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17678 13812 17684 13864
rect 17736 13852 17742 13864
rect 18322 13852 18328 13864
rect 17736 13824 18328 13852
rect 17736 13812 17742 13824
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 20070 13812 20076 13864
rect 20128 13852 20134 13864
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 20128 13824 20545 13852
rect 20128 13812 20134 13824
rect 20533 13821 20545 13824
rect 20579 13852 20591 13855
rect 21100 13852 21128 13883
rect 20579 13824 21128 13852
rect 20579 13821 20591 13824
rect 20533 13815 20591 13821
rect 21266 13812 21272 13864
rect 21324 13812 21330 13864
rect 21726 13812 21732 13864
rect 21784 13852 21790 13864
rect 21913 13855 21971 13861
rect 21913 13852 21925 13855
rect 21784 13824 21925 13852
rect 21784 13812 21790 13824
rect 21913 13821 21925 13824
rect 21959 13852 21971 13855
rect 22066 13852 22094 13892
rect 21959 13824 22094 13852
rect 22204 13852 22232 13892
rect 22278 13880 22284 13932
rect 22336 13880 22342 13932
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 24489 13923 24547 13929
rect 24489 13920 24501 13923
rect 23900 13892 24501 13920
rect 23900 13880 23906 13892
rect 24489 13889 24501 13892
rect 24535 13889 24547 13923
rect 24489 13883 24547 13889
rect 23750 13852 23756 13864
rect 22204 13824 23756 13852
rect 21959 13821 21971 13824
rect 21913 13815 21971 13821
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 25501 13855 25559 13861
rect 25501 13821 25513 13855
rect 25547 13852 25559 13855
rect 25590 13852 25596 13864
rect 25547 13824 25596 13852
rect 25547 13821 25559 13824
rect 25501 13815 25559 13821
rect 25590 13812 25596 13824
rect 25648 13812 25654 13864
rect 3326 13744 3332 13796
rect 3384 13784 3390 13796
rect 4522 13784 4528 13796
rect 3384 13756 4528 13784
rect 3384 13744 3390 13756
rect 4522 13744 4528 13756
rect 4580 13744 4586 13796
rect 4706 13744 4712 13796
rect 4764 13784 4770 13796
rect 7282 13784 7288 13796
rect 4764 13756 7288 13784
rect 4764 13744 4770 13756
rect 7282 13744 7288 13756
rect 7340 13744 7346 13796
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 11514 13784 11520 13796
rect 10836 13756 11520 13784
rect 10836 13744 10842 13756
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 12618 13744 12624 13796
rect 12676 13784 12682 13796
rect 13630 13784 13636 13796
rect 12676 13756 13636 13784
rect 12676 13744 12682 13756
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 15838 13744 15844 13796
rect 15896 13784 15902 13796
rect 18414 13784 18420 13796
rect 15896 13756 18420 13784
rect 15896 13744 15902 13756
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 20898 13744 20904 13796
rect 20956 13784 20962 13796
rect 21174 13784 21180 13796
rect 20956 13756 21180 13784
rect 20956 13744 20962 13756
rect 21174 13744 21180 13756
rect 21232 13744 21238 13796
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 6086 13716 6092 13728
rect 4028 13688 6092 13716
rect 4028 13676 4034 13688
rect 6086 13676 6092 13688
rect 6144 13676 6150 13728
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 11146 13716 11152 13728
rect 9364 13688 11152 13716
rect 9364 13676 9370 13688
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 13896 13719 13954 13725
rect 13896 13685 13908 13719
rect 13942 13716 13954 13719
rect 15102 13716 15108 13728
rect 13942 13688 15108 13716
rect 13942 13685 13954 13688
rect 13896 13679 13954 13685
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 21358 13716 21364 13728
rect 15252 13688 21364 13716
rect 15252 13676 15258 13688
rect 21358 13676 21364 13688
rect 21416 13676 21422 13728
rect 22544 13719 22602 13725
rect 22544 13685 22556 13719
rect 22590 13716 22602 13719
rect 25406 13716 25412 13728
rect 22590 13688 25412 13716
rect 22590 13685 22602 13688
rect 22544 13679 22602 13685
rect 25406 13676 25412 13688
rect 25464 13676 25470 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 2406 13512 2412 13524
rect 2363 13484 2412 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 2958 13512 2964 13524
rect 2556 13484 2964 13512
rect 2556 13472 2562 13484
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 3234 13472 3240 13524
rect 3292 13472 3298 13524
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4706 13512 4712 13524
rect 4212 13484 4712 13512
rect 4212 13472 4218 13484
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 5442 13472 5448 13524
rect 5500 13472 5506 13524
rect 6730 13512 6736 13524
rect 5552 13484 6736 13512
rect 2777 13447 2835 13453
rect 2777 13413 2789 13447
rect 2823 13444 2835 13447
rect 4430 13444 4436 13456
rect 2823 13416 4436 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 4430 13404 4436 13416
rect 4488 13404 4494 13456
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 3973 13379 4031 13385
rect 3973 13376 3985 13379
rect 2188 13348 3985 13376
rect 2188 13336 2194 13348
rect 3973 13345 3985 13348
rect 4019 13345 4031 13379
rect 3973 13339 4031 13345
rect 4246 13336 4252 13388
rect 4304 13336 4310 13388
rect 5552 13376 5580 13484
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 7064 13484 8585 13512
rect 7064 13472 7070 13484
rect 8573 13481 8585 13484
rect 8619 13481 8631 13515
rect 8573 13475 8631 13481
rect 8938 13472 8944 13524
rect 8996 13472 9002 13524
rect 9214 13472 9220 13524
rect 9272 13472 9278 13524
rect 10134 13512 10140 13524
rect 9646 13484 10140 13512
rect 6086 13404 6092 13456
rect 6144 13444 6150 13456
rect 6144 13416 6960 13444
rect 6144 13404 6150 13416
rect 5092 13348 5580 13376
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 1673 13311 1731 13317
rect 1673 13308 1685 13311
rect 1360 13280 1685 13308
rect 1360 13268 1366 13280
rect 1673 13277 1685 13280
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 2866 13268 2872 13320
rect 2924 13308 2930 13320
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 2924 13280 3433 13308
rect 2924 13268 2930 13280
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 2372 13212 2774 13240
rect 2372 13200 2378 13212
rect 2746 13172 2774 13212
rect 2958 13200 2964 13252
rect 3016 13240 3022 13252
rect 3786 13240 3792 13252
rect 3016 13212 3792 13240
rect 3016 13200 3022 13212
rect 3786 13200 3792 13212
rect 3844 13200 3850 13252
rect 5092 13172 5120 13348
rect 5626 13336 5632 13388
rect 5684 13376 5690 13388
rect 6932 13376 6960 13416
rect 9122 13404 9128 13456
rect 9180 13444 9186 13456
rect 9646 13444 9674 13484
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10594 13472 10600 13524
rect 10652 13512 10658 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10652 13484 10793 13512
rect 10652 13472 10658 13484
rect 10781 13481 10793 13484
rect 10827 13481 10839 13515
rect 10781 13475 10839 13481
rect 11514 13472 11520 13524
rect 11572 13512 11578 13524
rect 12618 13512 12624 13524
rect 11572 13484 12624 13512
rect 11572 13472 11578 13484
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 15013 13515 15071 13521
rect 15013 13512 15025 13515
rect 14884 13484 15025 13512
rect 14884 13472 14890 13484
rect 15013 13481 15025 13484
rect 15059 13481 15071 13515
rect 17126 13512 17132 13524
rect 15013 13475 15071 13481
rect 15120 13484 17132 13512
rect 9180 13416 9674 13444
rect 13449 13447 13507 13453
rect 9180 13404 9186 13416
rect 13449 13413 13461 13447
rect 13495 13444 13507 13447
rect 15120 13444 15148 13484
rect 17126 13472 17132 13484
rect 17184 13472 17190 13524
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 17920 13484 23428 13512
rect 17920 13472 17926 13484
rect 13495 13416 15148 13444
rect 17957 13447 18015 13453
rect 13495 13413 13507 13416
rect 13449 13407 13507 13413
rect 17957 13413 17969 13447
rect 18003 13444 18015 13447
rect 18782 13444 18788 13456
rect 18003 13416 18788 13444
rect 18003 13413 18015 13416
rect 17957 13407 18015 13413
rect 9950 13376 9956 13388
rect 5684 13348 6868 13376
rect 6932 13348 9956 13376
rect 5684 13336 5690 13348
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5721 13311 5779 13317
rect 5721 13308 5733 13311
rect 5307 13280 5733 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5721 13277 5733 13280
rect 5767 13308 5779 13311
rect 6454 13308 6460 13320
rect 5767 13280 6460 13308
rect 5767 13277 5779 13280
rect 5721 13271 5779 13277
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 6840 13317 6868 13348
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10042 13336 10048 13388
rect 10100 13376 10106 13388
rect 10594 13376 10600 13388
rect 10100 13348 10600 13376
rect 10100 13336 10106 13348
rect 10594 13336 10600 13348
rect 10652 13376 10658 13388
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 10652 13348 11713 13376
rect 10652 13336 10658 13348
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 7098 13268 7104 13320
rect 7156 13308 7162 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7156 13280 7941 13308
rect 7156 13268 7162 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 9582 13308 9588 13320
rect 9539 13280 9588 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 5166 13200 5172 13252
rect 5224 13240 5230 13252
rect 7190 13240 7196 13252
rect 5224 13212 7196 13240
rect 5224 13200 5230 13212
rect 7190 13200 7196 13212
rect 7248 13200 7254 13252
rect 7469 13243 7527 13249
rect 7469 13209 7481 13243
rect 7515 13240 7527 13243
rect 7515 13212 9536 13240
rect 7515 13209 7527 13212
rect 7469 13203 7527 13209
rect 9508 13184 9536 13212
rect 11146 13200 11152 13252
rect 11204 13240 11210 13252
rect 11977 13243 12035 13249
rect 11977 13240 11989 13243
rect 11204 13212 11989 13240
rect 11204 13200 11210 13212
rect 11977 13209 11989 13212
rect 12023 13209 12035 13243
rect 11977 13203 12035 13209
rect 12250 13200 12256 13252
rect 12308 13240 12314 13252
rect 12308 13212 12466 13240
rect 12308 13200 12314 13212
rect 13464 13184 13492 13407
rect 18782 13404 18788 13416
rect 18840 13404 18846 13456
rect 21174 13404 21180 13456
rect 21232 13444 21238 13456
rect 21358 13444 21364 13456
rect 21232 13416 21364 13444
rect 21232 13404 21238 13416
rect 21358 13404 21364 13416
rect 21416 13404 21422 13456
rect 23400 13444 23428 13484
rect 23474 13472 23480 13524
rect 23532 13512 23538 13524
rect 23661 13515 23719 13521
rect 23661 13512 23673 13515
rect 23532 13484 23673 13512
rect 23532 13472 23538 13484
rect 23661 13481 23673 13484
rect 23707 13512 23719 13515
rect 23934 13512 23940 13524
rect 23707 13484 23940 13512
rect 23707 13481 23719 13484
rect 23661 13475 23719 13481
rect 23934 13472 23940 13484
rect 23992 13472 23998 13524
rect 24029 13515 24087 13521
rect 24029 13481 24041 13515
rect 24075 13512 24087 13515
rect 24670 13512 24676 13524
rect 24075 13484 24676 13512
rect 24075 13481 24087 13484
rect 24029 13475 24087 13481
rect 24670 13472 24676 13484
rect 24728 13472 24734 13524
rect 25225 13515 25283 13521
rect 25225 13481 25237 13515
rect 25271 13512 25283 13515
rect 26878 13512 26884 13524
rect 25271 13484 26884 13512
rect 25271 13481 25283 13484
rect 25225 13475 25283 13481
rect 26878 13472 26884 13484
rect 26936 13472 26942 13524
rect 24688 13444 24716 13472
rect 26234 13444 26240 13456
rect 23400 13416 23704 13444
rect 24688 13416 26240 13444
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 15378 13376 15384 13388
rect 14516 13348 15384 13376
rect 14516 13336 14522 13348
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 16666 13376 16672 13388
rect 15703 13348 16672 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 18509 13379 18567 13385
rect 18509 13376 18521 13379
rect 17420 13348 18521 13376
rect 14366 13268 14372 13320
rect 14424 13268 14430 13320
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 15010 13308 15016 13320
rect 14792 13280 15016 13308
rect 14792 13268 14798 13280
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 17034 13268 17040 13320
rect 17092 13268 17098 13320
rect 15933 13243 15991 13249
rect 15304 13212 15516 13240
rect 2746 13144 5120 13172
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6052 13144 6377 13172
rect 6052 13132 6058 13144
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 6638 13132 6644 13184
rect 6696 13172 6702 13184
rect 7006 13172 7012 13184
rect 6696 13144 7012 13172
rect 6696 13132 6702 13144
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 9490 13132 9496 13184
rect 9548 13132 9554 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 13262 13172 13268 13184
rect 11112 13144 13268 13172
rect 11112 13132 11118 13144
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 13446 13132 13452 13184
rect 13504 13132 13510 13184
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 15304 13172 15332 13212
rect 15488 13184 15516 13212
rect 15933 13209 15945 13243
rect 15979 13240 15991 13243
rect 16206 13240 16212 13252
rect 15979 13212 16212 13240
rect 15979 13209 15991 13212
rect 15933 13203 15991 13209
rect 16206 13200 16212 13212
rect 16264 13200 16270 13252
rect 13964 13144 15332 13172
rect 13964 13132 13970 13144
rect 15378 13132 15384 13184
rect 15436 13132 15442 13184
rect 15470 13132 15476 13184
rect 15528 13132 15534 13184
rect 16666 13132 16672 13184
rect 16724 13172 16730 13184
rect 17420 13181 17448 13348
rect 18509 13345 18521 13348
rect 18555 13345 18567 13379
rect 18509 13339 18567 13345
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19392 13348 19717 13376
rect 19392 13336 19398 13348
rect 19705 13345 19717 13348
rect 19751 13376 19763 13379
rect 21910 13376 21916 13388
rect 19751 13348 21916 13376
rect 19751 13345 19763 13348
rect 19705 13339 19763 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22189 13379 22247 13385
rect 22189 13345 22201 13379
rect 22235 13376 22247 13379
rect 23566 13376 23572 13388
rect 22235 13348 23572 13376
rect 22235 13345 22247 13348
rect 22189 13339 22247 13345
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 23676 13376 23704 13416
rect 26234 13404 26240 13416
rect 26292 13404 26298 13456
rect 25222 13376 25228 13388
rect 23676 13348 25228 13376
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13308 24639 13311
rect 24946 13308 24952 13320
rect 24627 13280 24952 13308
rect 24627 13277 24639 13280
rect 24581 13271 24639 13277
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 18417 13243 18475 13249
rect 18417 13209 18429 13243
rect 18463 13240 18475 13243
rect 18506 13240 18512 13252
rect 18463 13212 18512 13240
rect 18463 13209 18475 13212
rect 18417 13203 18475 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 19518 13240 19524 13252
rect 18984 13212 19524 13240
rect 18984 13184 19012 13212
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 19978 13200 19984 13252
rect 20036 13200 20042 13252
rect 23658 13240 23664 13252
rect 21206 13212 21956 13240
rect 23414 13212 23664 13240
rect 17405 13175 17463 13181
rect 17405 13172 17417 13175
rect 16724 13144 17417 13172
rect 16724 13132 16730 13144
rect 17405 13141 17417 13144
rect 17451 13141 17463 13175
rect 17405 13135 17463 13141
rect 18322 13132 18328 13184
rect 18380 13132 18386 13184
rect 18966 13132 18972 13184
rect 19024 13132 19030 13184
rect 19429 13175 19487 13181
rect 19429 13141 19441 13175
rect 19475 13172 19487 13175
rect 19702 13172 19708 13184
rect 19475 13144 19708 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 19702 13132 19708 13144
rect 19760 13172 19766 13184
rect 19886 13172 19892 13184
rect 19760 13144 19892 13172
rect 19760 13132 19766 13144
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 21284 13172 21312 13212
rect 20772 13144 21312 13172
rect 20772 13132 20778 13144
rect 21450 13132 21456 13184
rect 21508 13132 21514 13184
rect 21928 13172 21956 13212
rect 23492 13172 23520 13212
rect 23658 13200 23664 13212
rect 23716 13200 23722 13252
rect 24213 13243 24271 13249
rect 24213 13209 24225 13243
rect 24259 13240 24271 13243
rect 24762 13240 24768 13252
rect 24259 13212 24768 13240
rect 24259 13209 24271 13212
rect 24213 13203 24271 13209
rect 24762 13200 24768 13212
rect 24820 13240 24826 13252
rect 25590 13240 25596 13252
rect 24820 13212 25596 13240
rect 24820 13200 24826 13212
rect 25590 13200 25596 13212
rect 25648 13200 25654 13252
rect 21928 13144 23520 13172
rect 24578 13132 24584 13184
rect 24636 13172 24642 13184
rect 24946 13172 24952 13184
rect 24636 13144 24952 13172
rect 24636 13132 24642 13144
rect 24946 13132 24952 13144
rect 25004 13132 25010 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 2038 12928 2044 12980
rect 2096 12928 2102 12980
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 4672 12940 4721 12968
rect 4672 12928 4678 12940
rect 4709 12937 4721 12940
rect 4755 12968 4767 12971
rect 4798 12968 4804 12980
rect 4755 12940 4804 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12968 5043 12971
rect 5077 12971 5135 12977
rect 5077 12968 5089 12971
rect 5031 12940 5089 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 5077 12937 5089 12940
rect 5123 12968 5135 12971
rect 5166 12968 5172 12980
rect 5123 12940 5172 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5810 12928 5816 12980
rect 5868 12928 5874 12980
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 6822 12968 6828 12980
rect 6595 12940 6828 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 10045 12971 10103 12977
rect 10045 12968 10057 12971
rect 7852 12940 10057 12968
rect 4433 12903 4491 12909
rect 4433 12869 4445 12903
rect 4479 12900 4491 12903
rect 4890 12900 4896 12912
rect 4479 12872 4896 12900
rect 4479 12869 4491 12872
rect 4433 12863 4491 12869
rect 4890 12860 4896 12872
rect 4948 12860 4954 12912
rect 6178 12860 6184 12912
rect 6236 12900 6242 12912
rect 7852 12900 7880 12940
rect 10045 12937 10057 12940
rect 10091 12937 10103 12971
rect 10045 12931 10103 12937
rect 11146 12928 11152 12980
rect 11204 12928 11210 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 13906 12968 13912 12980
rect 11756 12940 13912 12968
rect 11756 12928 11762 12940
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 14274 12928 14280 12980
rect 14332 12968 14338 12980
rect 14332 12940 14872 12968
rect 14332 12928 14338 12940
rect 6236 12872 7880 12900
rect 6236 12860 6242 12872
rect 7926 12860 7932 12912
rect 7984 12900 7990 12912
rect 7984 12872 10640 12900
rect 7984 12860 7990 12872
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 3602 12832 3608 12844
rect 3559 12804 3608 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 1964 12696 1992 12795
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 4663 12804 6745 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 6733 12801 6745 12804
rect 6779 12832 6791 12835
rect 6822 12832 6828 12844
rect 6779 12804 6828 12832
rect 6779 12801 6791 12804
rect 6733 12795 6791 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 6972 12804 7205 12832
rect 6972 12792 6978 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12832 8723 12835
rect 8938 12832 8944 12844
rect 8711 12804 8944 12832
rect 8711 12801 8723 12804
rect 8665 12795 8723 12801
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 9122 12792 9128 12844
rect 9180 12792 9186 12844
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 10226 12832 10232 12844
rect 9447 12804 10232 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 10502 12792 10508 12844
rect 10560 12792 10566 12844
rect 10612 12832 10640 12872
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 12434 12900 12440 12912
rect 11112 12872 12440 12900
rect 11112 12860 11118 12872
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 12805 12903 12863 12909
rect 12805 12869 12817 12903
rect 12851 12900 12863 12903
rect 13541 12903 13599 12909
rect 13541 12900 13553 12903
rect 12851 12872 13553 12900
rect 12851 12869 12863 12872
rect 12805 12863 12863 12869
rect 13541 12869 13553 12872
rect 13587 12869 13599 12903
rect 14844 12900 14872 12940
rect 15010 12928 15016 12980
rect 15068 12928 15074 12980
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 15930 12968 15936 12980
rect 15436 12940 15936 12968
rect 15436 12928 15442 12940
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 16301 12971 16359 12977
rect 16301 12937 16313 12971
rect 16347 12968 16359 12971
rect 16574 12968 16580 12980
rect 16347 12940 16580 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 18966 12968 18972 12980
rect 16960 12940 18972 12968
rect 16960 12900 16988 12940
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19306 12940 19441 12968
rect 14844 12872 16988 12900
rect 13541 12863 13599 12869
rect 17126 12860 17132 12912
rect 17184 12900 17190 12912
rect 17184 12872 17618 12900
rect 17184 12860 17190 12872
rect 19150 12860 19156 12912
rect 19208 12900 19214 12912
rect 19306 12900 19334 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19429 12931 19487 12937
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 19576 12940 20392 12968
rect 19576 12928 19582 12940
rect 20254 12900 20260 12912
rect 19208 12872 19334 12900
rect 19536 12872 20260 12900
rect 19208 12860 19214 12872
rect 11514 12832 11520 12844
rect 10612 12804 11520 12832
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 12158 12792 12164 12844
rect 12216 12792 12222 12844
rect 12618 12792 12624 12844
rect 12676 12832 12682 12844
rect 13170 12832 13176 12844
rect 12676 12804 13176 12832
rect 12676 12792 12682 12804
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 14642 12792 14648 12844
rect 14700 12792 14706 12844
rect 15657 12835 15715 12841
rect 15657 12801 15669 12835
rect 15703 12832 15715 12835
rect 16298 12832 16304 12844
rect 15703 12804 16304 12832
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 2590 12724 2596 12776
rect 2648 12724 2654 12776
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 3237 12767 3295 12773
rect 3237 12764 3249 12767
rect 2832 12736 3249 12764
rect 2832 12724 2838 12736
rect 3237 12733 3249 12736
rect 3283 12733 3295 12767
rect 3237 12727 3295 12733
rect 7466 12724 7472 12776
rect 7524 12724 7530 12776
rect 10042 12724 10048 12776
rect 10100 12764 10106 12776
rect 13265 12767 13323 12773
rect 13265 12764 13277 12767
rect 10100 12736 13277 12764
rect 10100 12724 10106 12736
rect 13265 12733 13277 12736
rect 13311 12733 13323 12767
rect 14660 12764 14688 12792
rect 15746 12764 15752 12776
rect 13265 12727 13323 12733
rect 13372 12736 14688 12764
rect 14844 12736 15752 12764
rect 7282 12696 7288 12708
rect 1964 12668 7288 12696
rect 7282 12656 7288 12668
rect 7340 12656 7346 12708
rect 8481 12699 8539 12705
rect 8481 12665 8493 12699
rect 8527 12696 8539 12699
rect 11422 12696 11428 12708
rect 8527 12668 11428 12696
rect 8527 12665 8539 12668
rect 8481 12659 8539 12665
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 11514 12656 11520 12708
rect 11572 12696 11578 12708
rect 12250 12696 12256 12708
rect 11572 12668 12256 12696
rect 11572 12656 11578 12668
rect 12250 12656 12256 12668
rect 12308 12696 12314 12708
rect 13372 12696 13400 12736
rect 12308 12668 13400 12696
rect 12308 12656 12314 12668
rect 14642 12656 14648 12708
rect 14700 12696 14706 12708
rect 14844 12696 14872 12736
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 17678 12764 17684 12776
rect 17175 12736 17684 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 19536 12773 19564 12872
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 20364 12832 20392 12940
rect 20622 12928 20628 12980
rect 20680 12968 20686 12980
rect 20717 12971 20775 12977
rect 20717 12968 20729 12971
rect 20680 12940 20729 12968
rect 20680 12928 20686 12940
rect 20717 12937 20729 12940
rect 20763 12937 20775 12971
rect 20717 12931 20775 12937
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 21545 12971 21603 12977
rect 21545 12968 21557 12971
rect 21232 12940 21557 12968
rect 21232 12928 21238 12940
rect 21545 12937 21557 12940
rect 21591 12937 21603 12971
rect 21545 12931 21603 12937
rect 21726 12928 21732 12980
rect 21784 12968 21790 12980
rect 21913 12971 21971 12977
rect 21913 12968 21925 12971
rect 21784 12940 21925 12968
rect 21784 12928 21790 12940
rect 21913 12937 21925 12940
rect 21959 12937 21971 12971
rect 21913 12931 21971 12937
rect 22370 12928 22376 12980
rect 22428 12968 22434 12980
rect 22830 12968 22836 12980
rect 22428 12940 22836 12968
rect 22428 12928 22434 12940
rect 22830 12928 22836 12940
rect 22888 12928 22894 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 24121 12971 24179 12977
rect 24121 12968 24133 12971
rect 23532 12940 24133 12968
rect 23532 12928 23538 12940
rect 24121 12937 24133 12940
rect 24167 12968 24179 12971
rect 24486 12968 24492 12980
rect 24167 12940 24492 12968
rect 24167 12937 24179 12940
rect 24121 12931 24179 12937
rect 24486 12928 24492 12940
rect 24544 12928 24550 12980
rect 20438 12860 20444 12912
rect 20496 12900 20502 12912
rect 20990 12900 20996 12912
rect 20496 12872 20996 12900
rect 20496 12860 20502 12872
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 22922 12900 22928 12912
rect 21100 12872 22928 12900
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20364 12804 20637 12832
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 21100 12832 21128 12872
rect 22922 12860 22928 12872
rect 22980 12860 22986 12912
rect 23658 12860 23664 12912
rect 23716 12860 23722 12912
rect 20625 12795 20683 12801
rect 20732 12804 21128 12832
rect 21453 12835 21511 12841
rect 19521 12767 19579 12773
rect 18656 12736 19196 12764
rect 18656 12724 18662 12736
rect 19061 12699 19119 12705
rect 19061 12696 19073 12699
rect 14700 12668 14872 12696
rect 14936 12668 15424 12696
rect 14700 12656 14706 12668
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6546 12628 6552 12640
rect 6144 12600 6552 12628
rect 6144 12588 6150 12600
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 14936 12628 14964 12668
rect 6880 12600 14964 12628
rect 6880 12588 6886 12600
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15289 12631 15347 12637
rect 15289 12628 15301 12631
rect 15252 12600 15301 12628
rect 15252 12588 15258 12600
rect 15289 12597 15301 12600
rect 15335 12597 15347 12631
rect 15396 12628 15424 12668
rect 18156 12668 19073 12696
rect 18156 12628 18184 12668
rect 19061 12665 19073 12668
rect 19107 12665 19119 12699
rect 19168 12696 19196 12736
rect 19521 12733 19533 12767
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 20732 12764 20760 12804
rect 21453 12801 21465 12835
rect 21499 12832 21511 12835
rect 21726 12832 21732 12844
rect 21499 12804 21732 12832
rect 21499 12801 21511 12804
rect 21453 12795 21511 12801
rect 21726 12792 21732 12804
rect 21784 12792 21790 12844
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 21968 12804 22385 12832
rect 21968 12792 21974 12804
rect 22373 12801 22385 12804
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 24026 12792 24032 12844
rect 24084 12832 24090 12844
rect 24581 12835 24639 12841
rect 24581 12832 24593 12835
rect 24084 12804 24593 12832
rect 24084 12792 24090 12804
rect 24581 12801 24593 12804
rect 24627 12801 24639 12835
rect 24581 12795 24639 12801
rect 19613 12727 19671 12733
rect 19720 12736 20760 12764
rect 20901 12767 20959 12773
rect 19628 12696 19656 12727
rect 19168 12668 19656 12696
rect 19061 12659 19119 12665
rect 15396 12600 18184 12628
rect 15289 12591 15347 12597
rect 18874 12588 18880 12640
rect 18932 12588 18938 12640
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 19720 12628 19748 12736
rect 20901 12733 20913 12767
rect 20947 12764 20959 12767
rect 21174 12764 21180 12776
rect 20947 12736 21180 12764
rect 20947 12733 20959 12736
rect 20901 12727 20959 12733
rect 21174 12724 21180 12736
rect 21232 12724 21238 12776
rect 26142 12764 26148 12776
rect 22480 12736 26148 12764
rect 20530 12656 20536 12708
rect 20588 12696 20594 12708
rect 22480 12696 22508 12736
rect 26142 12724 26148 12736
rect 26200 12724 26206 12776
rect 20588 12668 22508 12696
rect 20588 12656 20594 12668
rect 19208 12600 19748 12628
rect 19208 12588 19214 12600
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21450 12628 21456 12640
rect 20864 12600 21456 12628
rect 20864 12588 20870 12600
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 21818 12588 21824 12640
rect 21876 12628 21882 12640
rect 22002 12628 22008 12640
rect 21876 12600 22008 12628
rect 21876 12588 21882 12600
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22370 12628 22376 12640
rect 22152 12600 22376 12628
rect 22152 12588 22158 12600
rect 22370 12588 22376 12600
rect 22428 12588 22434 12640
rect 22646 12637 22652 12640
rect 22630 12631 22652 12637
rect 22630 12597 22642 12631
rect 22630 12591 22652 12597
rect 22646 12588 22652 12591
rect 22704 12588 22710 12640
rect 25225 12631 25283 12637
rect 25225 12597 25237 12631
rect 25271 12628 25283 12631
rect 25314 12628 25320 12640
rect 25271 12600 25320 12628
rect 25271 12597 25283 12600
rect 25225 12591 25283 12597
rect 25314 12588 25320 12600
rect 25372 12588 25378 12640
rect 25958 12588 25964 12640
rect 26016 12628 26022 12640
rect 26142 12628 26148 12640
rect 26016 12600 26148 12628
rect 26016 12588 26022 12600
rect 26142 12588 26148 12600
rect 26200 12588 26206 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 2593 12427 2651 12433
rect 2593 12393 2605 12427
rect 2639 12424 2651 12427
rect 2774 12424 2780 12436
rect 2639 12396 2780 12424
rect 2639 12393 2651 12396
rect 2593 12387 2651 12393
rect 2774 12384 2780 12396
rect 2832 12384 2838 12436
rect 9125 12427 9183 12433
rect 9125 12393 9137 12427
rect 9171 12424 9183 12427
rect 10318 12424 10324 12436
rect 9171 12396 10324 12424
rect 9171 12393 9183 12396
rect 9125 12387 9183 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 12250 12424 12256 12436
rect 10560 12396 12256 12424
rect 10560 12384 10566 12396
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 12526 12384 12532 12436
rect 12584 12384 12590 12436
rect 12621 12427 12679 12433
rect 12621 12393 12633 12427
rect 12667 12424 12679 12427
rect 13722 12424 13728 12436
rect 12667 12396 13728 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 18509 12427 18567 12433
rect 18509 12424 18521 12427
rect 15160 12396 18521 12424
rect 15160 12384 15166 12396
rect 18509 12393 18521 12396
rect 18555 12393 18567 12427
rect 21174 12424 21180 12436
rect 18509 12387 18567 12393
rect 18984 12396 21180 12424
rect 2222 12316 2228 12368
rect 2280 12356 2286 12368
rect 2280 12328 5028 12356
rect 2280 12316 2286 12328
rect 842 12248 848 12300
rect 900 12288 906 12300
rect 5000 12297 5028 12328
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 9214 12356 9220 12368
rect 8444 12328 9220 12356
rect 8444 12316 8450 12328
rect 9214 12316 9220 12328
rect 9272 12316 9278 12368
rect 12544 12356 12572 12384
rect 18984 12368 19012 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 23753 12427 23811 12433
rect 23753 12424 23765 12427
rect 22152 12396 23765 12424
rect 22152 12384 22158 12396
rect 23753 12393 23765 12396
rect 23799 12393 23811 12427
rect 23753 12387 23811 12393
rect 24118 12384 24124 12436
rect 24176 12424 24182 12436
rect 24486 12424 24492 12436
rect 24176 12396 24492 12424
rect 24176 12384 24182 12396
rect 24486 12384 24492 12396
rect 24544 12384 24550 12436
rect 25314 12384 25320 12436
rect 25372 12424 25378 12436
rect 25372 12396 25544 12424
rect 25372 12384 25378 12396
rect 14921 12359 14979 12365
rect 14921 12356 14933 12359
rect 9508 12328 12480 12356
rect 12544 12328 14933 12356
rect 3237 12291 3295 12297
rect 3237 12288 3249 12291
rect 900 12260 3249 12288
rect 900 12248 906 12260
rect 3237 12257 3249 12260
rect 3283 12257 3295 12291
rect 3237 12251 3295 12257
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12288 6699 12291
rect 6917 12291 6975 12297
rect 6687 12260 6868 12288
rect 6687 12257 6699 12260
rect 6641 12251 6699 12257
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 2498 12220 2504 12232
rect 1903 12192 2504 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12220 2835 12223
rect 4154 12220 4160 12232
rect 2823 12192 4160 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12220 4307 12223
rect 4614 12220 4620 12232
rect 4295 12192 4620 12220
rect 4295 12189 4307 12192
rect 4249 12183 4307 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 5442 12220 5448 12232
rect 4755 12192 5448 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 6178 12180 6184 12232
rect 6236 12180 6242 12232
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 6454 12152 6460 12164
rect 5684 12124 6460 12152
rect 5684 12112 5690 12124
rect 6454 12112 6460 12124
rect 6512 12112 6518 12164
rect 4065 12087 4123 12093
rect 4065 12053 4077 12087
rect 4111 12084 4123 12087
rect 5902 12084 5908 12096
rect 4111 12056 5908 12084
rect 4111 12053 4123 12056
rect 4065 12047 4123 12053
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 5994 12044 6000 12096
rect 6052 12044 6058 12096
rect 6840 12084 6868 12260
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 9398 12288 9404 12300
rect 6963 12260 9404 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7708 12192 7941 12220
rect 7708 12180 7714 12192
rect 7929 12189 7941 12192
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 9180 12192 9321 12220
rect 9180 12180 9186 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 7466 12112 7472 12164
rect 7524 12152 7530 12164
rect 9508 12152 9536 12328
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 9640 12260 11100 12288
rect 9640 12248 9646 12260
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12220 9827 12223
rect 10226 12220 10232 12232
rect 9815 12192 10232 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 10962 12220 10968 12232
rect 10919 12192 10968 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 11072 12220 11100 12260
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 12452 12288 12480 12328
rect 14921 12325 14933 12328
rect 14967 12325 14979 12359
rect 14921 12319 14979 12325
rect 15286 12316 15292 12368
rect 15344 12316 15350 12368
rect 15470 12316 15476 12368
rect 15528 12356 15534 12368
rect 18322 12356 18328 12368
rect 15528 12328 18328 12356
rect 15528 12316 15534 12328
rect 18322 12316 18328 12328
rect 18380 12316 18386 12368
rect 18966 12316 18972 12368
rect 19024 12316 19030 12368
rect 21560 12328 22094 12356
rect 16758 12288 16764 12300
rect 11664 12260 12112 12288
rect 12452 12260 16764 12288
rect 11664 12248 11670 12260
rect 11790 12220 11796 12232
rect 11072 12192 11796 12220
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11974 12180 11980 12232
rect 12032 12180 12038 12232
rect 12084 12220 12112 12260
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 17034 12288 17040 12300
rect 16908 12260 17040 12288
rect 16908 12248 16914 12260
rect 17034 12248 17040 12260
rect 17092 12288 17098 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 17092 12260 19441 12288
rect 17092 12248 17098 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 19705 12291 19763 12297
rect 19705 12257 19717 12291
rect 19751 12288 19763 12291
rect 20162 12288 20168 12300
rect 19751 12260 20168 12288
rect 19751 12257 19763 12260
rect 19705 12251 19763 12257
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 21560 12297 21588 12328
rect 21545 12291 21603 12297
rect 21545 12257 21557 12291
rect 21591 12257 21603 12291
rect 22066 12288 22094 12328
rect 22830 12288 22836 12300
rect 22066 12260 22836 12288
rect 21545 12251 21603 12257
rect 22830 12248 22836 12260
rect 22888 12248 22894 12300
rect 24670 12288 24676 12300
rect 24136 12260 24676 12288
rect 24136 12232 24164 12260
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 25038 12248 25044 12300
rect 25096 12288 25102 12300
rect 25314 12288 25320 12300
rect 25096 12260 25320 12288
rect 25096 12248 25102 12260
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 12986 12220 12992 12232
rect 12084 12192 12992 12220
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13446 12220 13452 12232
rect 13127 12192 13452 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 14550 12220 14556 12232
rect 14323 12192 14556 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 15654 12180 15660 12232
rect 15712 12180 15718 12232
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 17865 12223 17923 12229
rect 17865 12220 17877 12223
rect 16724 12192 17877 12220
rect 16724 12180 16730 12192
rect 17865 12189 17877 12192
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 18506 12180 18512 12232
rect 18564 12220 18570 12232
rect 18785 12223 18843 12229
rect 18785 12220 18797 12223
rect 18564 12192 18797 12220
rect 18564 12180 18570 12192
rect 18785 12189 18797 12192
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 21910 12220 21916 12232
rect 21324 12192 21916 12220
rect 21324 12180 21330 12192
rect 21910 12180 21916 12192
rect 21968 12220 21974 12232
rect 22005 12223 22063 12229
rect 22005 12220 22017 12223
rect 21968 12192 22017 12220
rect 21968 12180 21974 12192
rect 22005 12189 22017 12192
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 24118 12180 24124 12232
rect 24176 12180 24182 12232
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12220 24639 12223
rect 24946 12220 24952 12232
rect 24627 12192 24952 12220
rect 24627 12189 24639 12192
rect 24581 12183 24639 12189
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 7524 12124 9536 12152
rect 10413 12155 10471 12161
rect 7524 12112 7530 12124
rect 10413 12121 10425 12155
rect 10459 12152 10471 12155
rect 19061 12155 19119 12161
rect 10459 12124 17816 12152
rect 10459 12121 10471 12124
rect 10413 12115 10471 12121
rect 8386 12084 8392 12096
rect 6840 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8570 12044 8576 12096
rect 8628 12044 8634 12096
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 11238 12084 11244 12096
rect 8904 12056 11244 12084
rect 8904 12044 8910 12056
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 11517 12087 11575 12093
rect 11517 12053 11529 12087
rect 11563 12084 11575 12087
rect 11606 12084 11612 12096
rect 11563 12056 11612 12084
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 13725 12087 13783 12093
rect 13725 12053 13737 12087
rect 13771 12084 13783 12087
rect 13906 12084 13912 12096
rect 13771 12056 13912 12084
rect 13771 12053 13783 12056
rect 13725 12047 13783 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 16482 12084 16488 12096
rect 16172 12056 16488 12084
rect 16172 12044 16178 12056
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 16942 12044 16948 12096
rect 17000 12044 17006 12096
rect 17788 12084 17816 12124
rect 19061 12121 19073 12155
rect 19107 12152 19119 12155
rect 19610 12152 19616 12164
rect 19107 12124 19616 12152
rect 19107 12121 19119 12124
rect 19061 12115 19119 12121
rect 19610 12112 19616 12124
rect 19668 12112 19674 12164
rect 20714 12112 20720 12164
rect 20772 12112 20778 12164
rect 22281 12155 22339 12161
rect 22281 12152 22293 12155
rect 21008 12124 22293 12152
rect 21008 12084 21036 12124
rect 22281 12121 22293 12124
rect 22327 12121 22339 12155
rect 23658 12152 23664 12164
rect 23506 12124 23664 12152
rect 22281 12115 22339 12121
rect 23658 12112 23664 12124
rect 23716 12112 23722 12164
rect 25516 12152 25544 12396
rect 25590 12316 25596 12368
rect 25648 12356 25654 12368
rect 25648 12328 25912 12356
rect 25648 12316 25654 12328
rect 25590 12152 25596 12164
rect 25516 12124 25596 12152
rect 25590 12112 25596 12124
rect 25648 12112 25654 12164
rect 17788 12056 21036 12084
rect 21542 12044 21548 12096
rect 21600 12084 21606 12096
rect 21637 12087 21695 12093
rect 21637 12084 21649 12087
rect 21600 12056 21649 12084
rect 21600 12044 21606 12056
rect 21637 12053 21649 12056
rect 21683 12053 21695 12087
rect 21637 12047 21695 12053
rect 23934 12044 23940 12096
rect 23992 12084 23998 12096
rect 24118 12084 24124 12096
rect 23992 12056 24124 12084
rect 23992 12044 23998 12056
rect 24118 12044 24124 12056
rect 24176 12044 24182 12096
rect 24578 12044 24584 12096
rect 24636 12084 24642 12096
rect 25225 12087 25283 12093
rect 25225 12084 25237 12087
rect 24636 12056 25237 12084
rect 24636 12044 24642 12056
rect 25225 12053 25237 12056
rect 25271 12053 25283 12087
rect 25225 12047 25283 12053
rect 25884 12016 25912 12328
rect 26326 12016 26332 12028
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 25884 11988 26332 12016
rect 26326 11976 26332 11988
rect 26384 11976 26390 12028
rect 1104 11920 25852 11942
rect 2774 11840 2780 11892
rect 2832 11840 2838 11892
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 2924 11852 3157 11880
rect 2924 11840 2930 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 8846 11880 8852 11892
rect 3145 11843 3203 11849
rect 3988 11852 8852 11880
rect 658 11772 664 11824
rect 716 11812 722 11824
rect 2792 11812 2820 11840
rect 716 11784 2728 11812
rect 2792 11784 2912 11812
rect 716 11772 722 11784
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 2038 11744 2044 11756
rect 1627 11716 2044 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2700 11753 2728 11784
rect 2884 11756 2912 11784
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11744 2743 11747
rect 2774 11744 2780 11756
rect 2731 11716 2780 11744
rect 2731 11713 2743 11716
rect 2685 11707 2743 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 2866 11704 2872 11756
rect 2924 11704 2930 11756
rect 3786 11704 3792 11756
rect 3844 11704 3850 11756
rect 2222 11636 2228 11688
rect 2280 11676 2286 11688
rect 3988 11676 4016 11852
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 9861 11883 9919 11889
rect 9861 11849 9873 11883
rect 9907 11880 9919 11883
rect 10134 11880 10140 11892
rect 9907 11852 10140 11880
rect 9907 11849 9919 11852
rect 9861 11843 9919 11849
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10962 11840 10968 11892
rect 11020 11840 11026 11892
rect 11238 11840 11244 11892
rect 11296 11840 11302 11892
rect 11606 11840 11612 11892
rect 11664 11840 11670 11892
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 12216 11852 13461 11880
rect 12216 11840 12222 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 13449 11843 13507 11849
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 14553 11883 14611 11889
rect 14553 11880 14565 11883
rect 14424 11852 14565 11880
rect 14424 11840 14430 11852
rect 14553 11849 14565 11852
rect 14599 11849 14611 11883
rect 14553 11843 14611 11849
rect 14918 11840 14924 11892
rect 14976 11880 14982 11892
rect 15013 11883 15071 11889
rect 15013 11880 15025 11883
rect 14976 11852 15025 11880
rect 14976 11840 14982 11852
rect 15013 11849 15025 11852
rect 15059 11849 15071 11883
rect 15013 11843 15071 11849
rect 16298 11840 16304 11892
rect 16356 11840 16362 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 17218 11880 17224 11892
rect 16540 11852 17224 11880
rect 16540 11840 16546 11852
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 21450 11880 21456 11892
rect 17696 11852 21456 11880
rect 7650 11812 7656 11824
rect 5184 11784 7656 11812
rect 5184 11753 5212 11784
rect 7650 11772 7656 11784
rect 7708 11772 7714 11824
rect 8570 11772 8576 11824
rect 8628 11812 8634 11824
rect 8628 11784 10180 11812
rect 8628 11772 8634 11784
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 5960 11716 6561 11744
rect 5960 11704 5966 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 2280 11648 4016 11676
rect 4065 11679 4123 11685
rect 2280 11636 2286 11648
rect 4065 11645 4077 11679
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 1854 11568 1860 11620
rect 1912 11568 1918 11620
rect 4080 11608 4108 11639
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 4396 11648 5457 11676
rect 4396 11636 4402 11648
rect 5445 11645 5457 11648
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 5592 11648 6837 11676
rect 5592 11636 5598 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 7944 11676 7972 11707
rect 9214 11704 9220 11756
rect 9272 11704 9278 11756
rect 10152 11744 10180 11784
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 10152 11716 10333 11744
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11624 11744 11652 11840
rect 12342 11772 12348 11824
rect 12400 11772 12406 11824
rect 17696 11812 17724 11852
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 21545 11883 21603 11889
rect 21545 11849 21557 11883
rect 21591 11880 21603 11883
rect 21634 11880 21640 11892
rect 21591 11852 21640 11880
rect 21591 11849 21603 11852
rect 21545 11843 21603 11849
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 25222 11880 25228 11892
rect 22066 11852 25228 11880
rect 12728 11784 17724 11812
rect 11689 11747 11747 11753
rect 11689 11744 11701 11747
rect 10928 11716 11100 11744
rect 11624 11716 11701 11744
rect 10928 11704 10934 11716
rect 9674 11676 9680 11688
rect 7944 11648 9680 11676
rect 6825 11639 6883 11645
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 11072 11676 11100 11716
rect 11689 11713 11701 11716
rect 11735 11713 11747 11747
rect 11689 11707 11747 11713
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 12728 11744 12756 11784
rect 18690 11772 18696 11824
rect 18748 11812 18754 11824
rect 19886 11812 19892 11824
rect 18748 11784 19892 11812
rect 18748 11772 18754 11784
rect 19886 11772 19892 11784
rect 19944 11772 19950 11824
rect 11848 11716 12756 11744
rect 12805 11747 12863 11753
rect 11848 11704 11854 11716
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 12820 11676 12848 11707
rect 13906 11704 13912 11756
rect 13964 11704 13970 11756
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11744 15715 11747
rect 16022 11744 16028 11756
rect 15703 11716 16028 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16298 11704 16304 11756
rect 16356 11744 16362 11756
rect 16356 11716 16988 11744
rect 16356 11704 16362 11716
rect 11072 11648 12848 11676
rect 12986 11636 12992 11688
rect 13044 11676 13050 11688
rect 16761 11679 16819 11685
rect 13044 11648 16712 11676
rect 13044 11636 13050 11648
rect 15286 11608 15292 11620
rect 4080 11580 15292 11608
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 7742 11540 7748 11552
rect 2547 11512 7748 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 8570 11500 8576 11552
rect 8628 11500 8634 11552
rect 8846 11500 8852 11552
rect 8904 11500 8910 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9582 11540 9588 11552
rect 9088 11512 9588 11540
rect 9088 11500 9094 11512
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 16684 11540 16712 11648
rect 16761 11645 16773 11679
rect 16807 11676 16819 11679
rect 16850 11676 16856 11688
rect 16807 11648 16856 11676
rect 16807 11645 16819 11648
rect 16761 11639 16819 11645
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 16960 11676 16988 11716
rect 17034 11704 17040 11756
rect 17092 11704 17098 11756
rect 18414 11704 18420 11756
rect 18472 11704 18478 11756
rect 19334 11704 19340 11756
rect 19392 11704 19398 11756
rect 20714 11704 20720 11756
rect 20772 11704 20778 11756
rect 20898 11704 20904 11756
rect 20956 11744 20962 11756
rect 21358 11744 21364 11756
rect 20956 11716 21364 11744
rect 20956 11704 20962 11716
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 21634 11704 21640 11756
rect 21692 11744 21698 11756
rect 22066 11744 22094 11852
rect 25222 11840 25228 11852
rect 25280 11840 25286 11892
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 21692 11716 22094 11744
rect 22281 11747 22339 11753
rect 21692 11704 21698 11716
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22738 11744 22744 11756
rect 22327 11716 22744 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22738 11704 22744 11716
rect 22796 11704 22802 11756
rect 23934 11704 23940 11756
rect 23992 11704 23998 11756
rect 24670 11704 24676 11756
rect 24728 11744 24734 11756
rect 26694 11744 26700 11756
rect 24728 11716 26700 11744
rect 24728 11704 24734 11716
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 17313 11679 17371 11685
rect 16960 11648 17172 11676
rect 16850 11540 16856 11552
rect 16684 11512 16856 11540
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17144 11540 17172 11648
rect 17313 11645 17325 11679
rect 17359 11676 17371 11679
rect 17678 11676 17684 11688
rect 17359 11648 17684 11676
rect 17359 11645 17371 11648
rect 17313 11639 17371 11645
rect 17678 11636 17684 11648
rect 17736 11636 17742 11688
rect 18966 11676 18972 11688
rect 18432 11648 18972 11676
rect 18432 11540 18460 11648
rect 18966 11636 18972 11648
rect 19024 11636 19030 11688
rect 19613 11679 19671 11685
rect 19613 11645 19625 11679
rect 19659 11676 19671 11679
rect 20346 11676 20352 11688
rect 19659 11648 20352 11676
rect 19659 11645 19671 11648
rect 19613 11639 19671 11645
rect 20346 11636 20352 11648
rect 20404 11636 20410 11688
rect 24946 11676 24952 11688
rect 20640 11648 24952 11676
rect 18506 11568 18512 11620
rect 18564 11608 18570 11620
rect 18564 11580 19472 11608
rect 18564 11568 18570 11580
rect 17144 11512 18460 11540
rect 18782 11500 18788 11552
rect 18840 11540 18846 11552
rect 19242 11540 19248 11552
rect 18840 11512 19248 11540
rect 18840 11500 18846 11512
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 19444 11540 19472 11580
rect 20640 11540 20668 11648
rect 24946 11636 24952 11648
rect 25004 11636 25010 11688
rect 20898 11568 20904 11620
rect 20956 11608 20962 11620
rect 23474 11608 23480 11620
rect 20956 11580 23480 11608
rect 20956 11568 20962 11580
rect 23474 11568 23480 11580
rect 23532 11568 23538 11620
rect 19444 11512 20668 11540
rect 21082 11500 21088 11552
rect 21140 11500 21146 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 1854 11296 1860 11348
rect 1912 11296 1918 11348
rect 2774 11296 2780 11348
rect 2832 11296 2838 11348
rect 3786 11296 3792 11348
rect 3844 11296 3850 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 6788 11308 7849 11336
rect 6788 11296 6794 11308
rect 7837 11305 7849 11308
rect 7883 11305 7895 11339
rect 7837 11299 7895 11305
rect 8386 11296 8392 11348
rect 8444 11296 8450 11348
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 10321 11339 10379 11345
rect 10321 11336 10333 11339
rect 9916 11308 10333 11336
rect 9916 11296 9922 11308
rect 10321 11305 10333 11308
rect 10367 11336 10379 11339
rect 10367 11308 10916 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 5721 11271 5779 11277
rect 5721 11268 5733 11271
rect 4540 11240 5733 11268
rect 4540 11209 4568 11240
rect 5721 11237 5733 11240
rect 5767 11268 5779 11271
rect 7006 11268 7012 11280
rect 5767 11240 7012 11268
rect 5767 11237 5779 11240
rect 5721 11231 5779 11237
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 9582 11268 9588 11280
rect 8628 11240 9588 11268
rect 8628 11228 8634 11240
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 10781 11271 10839 11277
rect 10781 11237 10793 11271
rect 10827 11237 10839 11271
rect 10888 11268 10916 11308
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 12032 11308 13185 11336
rect 12032 11296 12038 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 13173 11299 13231 11305
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 15654 11336 15660 11348
rect 13320 11308 15660 11336
rect 13320 11296 13326 11308
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 19150 11336 19156 11348
rect 15764 11308 19156 11336
rect 15764 11268 15792 11308
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 20530 11336 20536 11348
rect 19260 11308 20536 11336
rect 10888 11240 15792 11268
rect 10781 11231 10839 11237
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 5810 11200 5816 11212
rect 4847 11172 5816 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6641 11203 6699 11209
rect 6641 11169 6653 11203
rect 6687 11200 6699 11203
rect 7098 11200 7104 11212
rect 6687 11172 7104 11200
rect 6687 11169 6699 11172
rect 6641 11163 6699 11169
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11200 9183 11203
rect 9674 11200 9680 11212
rect 9171 11172 9680 11200
rect 9171 11169 9183 11172
rect 9125 11163 9183 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11200 10563 11203
rect 10594 11200 10600 11212
rect 10551 11172 10600 11200
rect 10551 11169 10563 11172
rect 10505 11163 10563 11169
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 10796 11200 10824 11231
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 18785 11271 18843 11277
rect 18785 11268 18797 11271
rect 18564 11240 18797 11268
rect 18564 11228 18570 11240
rect 18785 11237 18797 11240
rect 18831 11237 18843 11271
rect 18785 11231 18843 11237
rect 13538 11200 13544 11212
rect 10796 11172 13544 11200
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 16942 11200 16948 11212
rect 15703 11172 16948 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17126 11200 17132 11212
rect 17052 11172 17132 11200
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 1912 11104 2237 11132
rect 1912 11092 1918 11104
rect 2225 11101 2237 11104
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 3786 11132 3792 11144
rect 3467 11104 3792 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 6362 11092 6368 11144
rect 6420 11092 6426 11144
rect 7742 11092 7748 11144
rect 7800 11092 7806 11144
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 8846 11132 8852 11144
rect 8628 11104 8852 11132
rect 8628 11092 8634 11104
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 10870 11132 10876 11144
rect 9447 11104 10876 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 12529 11135 12587 11141
rect 11471 11104 12434 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 2406 11024 2412 11076
rect 2464 11024 2470 11076
rect 2498 11024 2504 11076
rect 2556 11064 2562 11076
rect 9306 11064 9312 11076
rect 2556 11036 9312 11064
rect 2556 11024 2562 11036
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 10594 11024 10600 11076
rect 10652 11064 10658 11076
rect 10980 11064 11008 11092
rect 10652 11036 11008 11064
rect 10652 11024 10658 11036
rect 12066 11024 12072 11076
rect 12124 11024 12130 11076
rect 12406 11064 12434 11104
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12618 11132 12624 11144
rect 12575 11104 12624 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12618 11092 12624 11104
rect 12676 11132 12682 11144
rect 13354 11132 13360 11144
rect 12676 11104 13360 11132
rect 12676 11092 12682 11104
rect 13354 11092 13360 11104
rect 13412 11132 13418 11144
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 13412 11104 13461 11132
rect 13412 11092 13418 11104
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 15010 11132 15016 11144
rect 14599 11104 15016 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 17052 11118 17080 11172
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 17402 11160 17408 11212
rect 17460 11160 17466 11212
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 19260 11200 19288 11308
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 21174 11296 21180 11348
rect 21232 11296 21238 11348
rect 22554 11336 22560 11348
rect 21284 11308 22560 11336
rect 19702 11228 19708 11280
rect 19760 11268 19766 11280
rect 21284 11268 21312 11308
rect 22554 11296 22560 11308
rect 22612 11296 22618 11348
rect 19760 11240 21312 11268
rect 19760 11228 19766 11240
rect 21450 11228 21456 11280
rect 21508 11268 21514 11280
rect 21508 11240 21956 11268
rect 21508 11228 21514 11240
rect 21928 11200 21956 11240
rect 22189 11203 22247 11209
rect 22189 11200 22201 11203
rect 18012 11172 19288 11200
rect 19444 11172 21864 11200
rect 21928 11172 22201 11200
rect 18012 11160 18018 11172
rect 17862 11092 17868 11144
rect 17920 11092 17926 11144
rect 19444 11141 19472 11172
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 20533 11135 20591 11141
rect 20533 11101 20545 11135
rect 20579 11132 20591 11135
rect 20622 11132 20628 11144
rect 20579 11104 20628 11132
rect 20579 11101 20591 11104
rect 20533 11095 20591 11101
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 21450 11092 21456 11144
rect 21508 11132 21514 11144
rect 21729 11135 21787 11141
rect 21729 11132 21741 11135
rect 21508 11104 21741 11132
rect 21508 11092 21514 11104
rect 21729 11101 21741 11104
rect 21775 11101 21787 11135
rect 21729 11095 21787 11101
rect 14918 11064 14924 11076
rect 12406 11036 14924 11064
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 15102 11024 15108 11076
rect 15160 11064 15166 11076
rect 15197 11067 15255 11073
rect 15197 11064 15209 11067
rect 15160 11036 15209 11064
rect 15160 11024 15166 11036
rect 15197 11033 15209 11036
rect 15243 11033 15255 11067
rect 15197 11027 15255 11033
rect 15933 11067 15991 11073
rect 15933 11033 15945 11067
rect 15979 11033 15991 11067
rect 18414 11064 18420 11076
rect 15933 11027 15991 11033
rect 17236 11036 18420 11064
rect 3234 10956 3240 11008
rect 3292 10956 3298 11008
rect 8754 10956 8760 11008
rect 8812 10996 8818 11008
rect 11146 10996 11152 11008
rect 8812 10968 11152 10996
rect 8812 10956 8818 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 12158 10956 12164 11008
rect 12216 10996 12222 11008
rect 12434 10996 12440 11008
rect 12216 10968 12440 10996
rect 12216 10956 12222 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 15948 10996 15976 11027
rect 16850 10996 16856 11008
rect 15948 10968 16856 10996
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17236 10996 17264 11036
rect 18414 11024 18420 11036
rect 18472 11064 18478 11076
rect 18969 11067 19027 11073
rect 18969 11064 18981 11067
rect 18472 11036 18981 11064
rect 18472 11024 18478 11036
rect 18969 11033 18981 11036
rect 19015 11033 19027 11067
rect 18969 11027 19027 11033
rect 19150 11024 19156 11076
rect 19208 11064 19214 11076
rect 20073 11067 20131 11073
rect 20073 11064 20085 11067
rect 19208 11036 20085 11064
rect 19208 11024 19214 11036
rect 20073 11033 20085 11036
rect 20119 11033 20131 11067
rect 20073 11027 20131 11033
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 20990 11064 20996 11076
rect 20220 11036 20996 11064
rect 20220 11024 20226 11036
rect 20990 11024 20996 11036
rect 21048 11024 21054 11076
rect 21836 11064 21864 11172
rect 22189 11169 22201 11172
rect 22235 11169 22247 11203
rect 22189 11163 22247 11169
rect 23845 11203 23903 11209
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 25038 11200 25044 11212
rect 23891 11172 25044 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 25038 11160 25044 11172
rect 25096 11160 25102 11212
rect 21910 11092 21916 11144
rect 21968 11092 21974 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 24578 11092 24584 11144
rect 24636 11092 24642 11144
rect 25498 11132 25504 11144
rect 24688 11104 25504 11132
rect 24688 11064 24716 11104
rect 25498 11092 25504 11104
rect 25556 11092 25562 11144
rect 21836 11036 24716 11064
rect 25222 11024 25228 11076
rect 25280 11024 25286 11076
rect 17000 10968 17264 10996
rect 17000 10956 17006 10968
rect 17494 10956 17500 11008
rect 17552 10996 17558 11008
rect 18046 10996 18052 11008
rect 17552 10968 18052 10996
rect 17552 10956 17558 10968
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 18506 10956 18512 11008
rect 18564 10956 18570 11008
rect 19242 10956 19248 11008
rect 19300 10996 19306 11008
rect 24210 10996 24216 11008
rect 19300 10968 24216 10996
rect 19300 10956 19306 10968
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 3329 10795 3387 10801
rect 3329 10792 3341 10795
rect 2148 10764 3341 10792
rect 2148 10665 2176 10764
rect 3329 10761 3341 10764
rect 3375 10792 3387 10795
rect 3694 10792 3700 10804
rect 3375 10764 3700 10792
rect 3375 10761 3387 10764
rect 3329 10755 3387 10761
rect 3694 10752 3700 10764
rect 3752 10752 3758 10804
rect 7098 10752 7104 10804
rect 7156 10752 7162 10804
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 7708 10764 7757 10792
rect 7708 10752 7714 10764
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 8389 10795 8447 10801
rect 8389 10761 8401 10795
rect 8435 10792 8447 10795
rect 12158 10792 12164 10804
rect 8435 10764 12164 10792
rect 8435 10761 8447 10764
rect 8389 10755 8447 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 13541 10795 13599 10801
rect 12308 10764 12572 10792
rect 12308 10752 12314 10764
rect 3234 10684 3240 10736
rect 3292 10724 3298 10736
rect 3789 10727 3847 10733
rect 3789 10724 3801 10727
rect 3292 10696 3801 10724
rect 3292 10684 3298 10696
rect 3789 10693 3801 10696
rect 3835 10693 3847 10727
rect 3789 10687 3847 10693
rect 3970 10684 3976 10736
rect 4028 10684 4034 10736
rect 11054 10724 11060 10736
rect 7944 10696 11060 10724
rect 7944 10665 7972 10696
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 11146 10684 11152 10736
rect 11204 10724 11210 10736
rect 12544 10724 12572 10764
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 13814 10792 13820 10804
rect 13587 10764 13820 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 15749 10795 15807 10801
rect 15749 10761 15761 10795
rect 15795 10792 15807 10795
rect 16666 10792 16672 10804
rect 15795 10764 16672 10792
rect 15795 10761 15807 10764
rect 15749 10755 15807 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 17770 10752 17776 10804
rect 17828 10792 17834 10804
rect 18693 10795 18751 10801
rect 18693 10792 18705 10795
rect 17828 10764 18705 10792
rect 17828 10752 17834 10764
rect 18693 10761 18705 10764
rect 18739 10761 18751 10795
rect 18693 10755 18751 10761
rect 18966 10752 18972 10804
rect 19024 10792 19030 10804
rect 20901 10795 20959 10801
rect 19024 10764 20852 10792
rect 19024 10752 19030 10764
rect 15470 10724 15476 10736
rect 11204 10696 12434 10724
rect 12544 10696 15476 10724
rect 11204 10684 11210 10696
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 2133 10619 2191 10625
rect 2332 10628 6745 10656
rect 1026 10548 1032 10600
rect 1084 10588 1090 10600
rect 2332 10588 2360 10628
rect 6733 10625 6745 10628
rect 6779 10656 6791 10659
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 6779 10628 7297 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10656 8631 10659
rect 8938 10656 8944 10668
rect 8619 10628 8944 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9214 10616 9220 10668
rect 9272 10616 9278 10668
rect 9858 10616 9864 10668
rect 9916 10616 9922 10668
rect 10594 10616 10600 10668
rect 10652 10616 10658 10668
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 12406 10656 12434 10696
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 17218 10684 17224 10736
rect 17276 10724 17282 10736
rect 19797 10727 19855 10733
rect 19797 10724 19809 10727
rect 17276 10696 19809 10724
rect 17276 10684 17282 10696
rect 19797 10693 19809 10696
rect 19843 10693 19855 10727
rect 19797 10687 19855 10693
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12406 10628 12909 10656
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 15102 10616 15108 10668
rect 15160 10616 15166 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 17310 10656 17316 10668
rect 16899 10628 17316 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18506 10656 18512 10668
rect 18095 10628 18512 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 19150 10616 19156 10668
rect 19208 10616 19214 10668
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10656 20315 10659
rect 20438 10656 20444 10668
rect 20303 10628 20444 10656
rect 20303 10625 20315 10628
rect 20257 10619 20315 10625
rect 20438 10616 20444 10628
rect 20496 10616 20502 10668
rect 20824 10656 20852 10764
rect 20901 10761 20913 10795
rect 20947 10792 20959 10795
rect 21174 10792 21180 10804
rect 20947 10764 21180 10792
rect 20947 10761 20959 10764
rect 20901 10755 20959 10761
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 21453 10795 21511 10801
rect 21453 10761 21465 10795
rect 21499 10792 21511 10795
rect 21726 10792 21732 10804
rect 21499 10764 21732 10792
rect 21499 10761 21511 10764
rect 21453 10755 21511 10761
rect 21726 10752 21732 10764
rect 21784 10752 21790 10804
rect 26510 10792 26516 10804
rect 21836 10764 26516 10792
rect 21836 10656 21864 10764
rect 26510 10752 26516 10764
rect 26568 10752 26574 10804
rect 25130 10684 25136 10736
rect 25188 10684 25194 10736
rect 20824 10628 21864 10656
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 1084 10560 2360 10588
rect 1084 10548 1090 10560
rect 2406 10548 2412 10600
rect 2464 10548 2470 10600
rect 4430 10548 4436 10600
rect 4488 10548 4494 10600
rect 4709 10591 4767 10597
rect 4709 10557 4721 10591
rect 4755 10588 4767 10591
rect 5166 10588 5172 10600
rect 4755 10560 5172 10588
rect 4755 10557 4767 10560
rect 4709 10551 4767 10557
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 5629 10523 5687 10529
rect 5629 10520 5641 10523
rect 2746 10492 5641 10520
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 2746 10452 2774 10492
rect 5629 10489 5641 10492
rect 5675 10520 5687 10523
rect 5828 10520 5856 10551
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 6512 10560 10333 10588
rect 6512 10548 6518 10560
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 14884 10560 21680 10588
rect 14884 10548 14890 10560
rect 5675 10492 5856 10520
rect 5675 10489 5687 10492
rect 5629 10483 5687 10489
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 8846 10520 8852 10532
rect 7892 10492 8852 10520
rect 7892 10480 7898 10492
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 9677 10523 9735 10529
rect 9677 10489 9689 10523
rect 9723 10520 9735 10523
rect 14458 10520 14464 10532
rect 9723 10492 14464 10520
rect 9723 10489 9735 10492
rect 9677 10483 9735 10489
rect 14458 10480 14464 10492
rect 14516 10480 14522 10532
rect 16114 10480 16120 10532
rect 16172 10520 16178 10532
rect 17770 10520 17776 10532
rect 16172 10492 17776 10520
rect 16172 10480 16178 10492
rect 17770 10480 17776 10492
rect 17828 10480 17834 10532
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 21542 10520 21548 10532
rect 20772 10492 21548 10520
rect 20772 10480 20778 10492
rect 21542 10480 21548 10492
rect 21600 10480 21606 10532
rect 21652 10520 21680 10560
rect 21726 10548 21732 10600
rect 21784 10588 21790 10600
rect 22112 10588 22140 10619
rect 23658 10616 23664 10668
rect 23716 10656 23722 10668
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 23716 10628 23949 10656
rect 23716 10616 23722 10628
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 21784 10560 22140 10588
rect 23293 10591 23351 10597
rect 21784 10548 21790 10560
rect 23293 10557 23305 10591
rect 23339 10588 23351 10591
rect 24854 10588 24860 10600
rect 23339 10560 24860 10588
rect 23339 10557 23351 10560
rect 23293 10551 23351 10557
rect 24854 10548 24860 10560
rect 24912 10548 24918 10600
rect 22094 10520 22100 10532
rect 21652 10492 22100 10520
rect 22094 10480 22100 10492
rect 22152 10480 22158 10532
rect 992 10424 2774 10452
rect 992 10412 998 10424
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 6454 10452 6460 10464
rect 3936 10424 6460 10452
rect 3936 10412 3942 10424
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 9033 10455 9091 10461
rect 9033 10421 9045 10455
rect 9079 10452 9091 10455
rect 11330 10452 11336 10464
rect 9079 10424 11336 10452
rect 9079 10421 9091 10424
rect 9033 10415 9091 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 14645 10455 14703 10461
rect 14645 10421 14657 10455
rect 14691 10452 14703 10455
rect 15654 10452 15660 10464
rect 14691 10424 15660 10452
rect 14691 10421 14703 10424
rect 14645 10415 14703 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 16022 10412 16028 10464
rect 16080 10412 16086 10464
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 17497 10455 17555 10461
rect 17497 10452 17509 10455
rect 17000 10424 17509 10452
rect 17000 10412 17006 10424
rect 17497 10421 17509 10424
rect 17543 10421 17555 10455
rect 17497 10415 17555 10421
rect 18506 10412 18512 10464
rect 18564 10452 18570 10464
rect 20070 10452 20076 10464
rect 18564 10424 20076 10452
rect 18564 10412 18570 10424
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 21174 10412 21180 10464
rect 21232 10452 21238 10464
rect 21269 10455 21327 10461
rect 21269 10452 21281 10455
rect 21232 10424 21281 10452
rect 21232 10412 21238 10424
rect 21269 10421 21281 10424
rect 21315 10452 21327 10455
rect 21818 10452 21824 10464
rect 21315 10424 21824 10452
rect 21315 10421 21327 10424
rect 21269 10415 21327 10421
rect 21818 10412 21824 10424
rect 21876 10412 21882 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 1544 10220 6040 10248
rect 1544 10208 1550 10220
rect 2314 10140 2320 10192
rect 2372 10140 2378 10192
rect 4430 10140 4436 10192
rect 4488 10180 4494 10192
rect 5353 10183 5411 10189
rect 5353 10180 5365 10183
rect 4488 10152 5365 10180
rect 4488 10140 4494 10152
rect 5353 10149 5365 10152
rect 5399 10149 5411 10183
rect 5353 10143 5411 10149
rect 5905 10183 5963 10189
rect 5905 10149 5917 10183
rect 5951 10149 5963 10183
rect 6012 10180 6040 10220
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 6604 10220 6745 10248
rect 6604 10208 6610 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 9125 10251 9183 10257
rect 9125 10217 9137 10251
rect 9171 10248 9183 10251
rect 9214 10248 9220 10260
rect 9171 10220 9220 10248
rect 9171 10217 9183 10220
rect 9125 10211 9183 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11664 10220 11713 10248
rect 11664 10208 11670 10220
rect 11701 10217 11713 10220
rect 11747 10248 11759 10251
rect 12342 10248 12348 10260
rect 11747 10220 12348 10248
rect 11747 10217 11759 10220
rect 11701 10211 11759 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 16485 10251 16543 10257
rect 16485 10248 16497 10251
rect 14056 10220 16497 10248
rect 14056 10208 14062 10220
rect 16485 10217 16497 10220
rect 16531 10217 16543 10251
rect 16485 10211 16543 10217
rect 18966 10208 18972 10260
rect 19024 10208 19030 10260
rect 19334 10208 19340 10260
rect 19392 10208 19398 10260
rect 20349 10251 20407 10257
rect 20349 10217 20361 10251
rect 20395 10248 20407 10251
rect 23842 10248 23848 10260
rect 20395 10220 23848 10248
rect 20395 10217 20407 10220
rect 20349 10211 20407 10217
rect 23842 10208 23848 10220
rect 23900 10208 23906 10260
rect 24210 10208 24216 10260
rect 24268 10208 24274 10260
rect 8297 10183 8355 10189
rect 8297 10180 8309 10183
rect 6012 10152 8309 10180
rect 5905 10143 5963 10149
rect 8297 10149 8309 10152
rect 8343 10149 8355 10183
rect 8297 10143 8355 10149
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 5920 10112 5948 10143
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 12621 10183 12679 10189
rect 10744 10152 12434 10180
rect 10744 10140 10750 10152
rect 4111 10084 5948 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 12406 10112 12434 10152
rect 12621 10149 12633 10183
rect 12667 10180 12679 10183
rect 12667 10152 16160 10180
rect 12667 10149 12679 10152
rect 12621 10143 12679 10149
rect 16022 10112 16028 10124
rect 6512 10084 10824 10112
rect 12406 10084 16028 10112
rect 6512 10072 6518 10084
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10044 2191 10047
rect 2179 10016 4292 10044
rect 2179 10013 2191 10016
rect 2133 10007 2191 10013
rect 2774 9936 2780 9988
rect 2832 9936 2838 9988
rect 4264 9976 4292 10016
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10044 5687 10047
rect 6086 10044 6092 10056
rect 5675 10016 6092 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 5994 9976 6000 9988
rect 4264 9948 6000 9976
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 6641 9979 6699 9985
rect 6641 9945 6653 9979
rect 6687 9976 6699 9979
rect 8386 9976 8392 9988
rect 6687 9948 8392 9976
rect 6687 9945 6699 9948
rect 6641 9939 6699 9945
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 8496 9976 8524 10007
rect 9398 10004 9404 10056
rect 9456 10004 9462 10056
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10044 9735 10047
rect 10410 10044 10416 10056
rect 9723 10016 10416 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 10594 10004 10600 10056
rect 10652 10044 10658 10056
rect 10689 10047 10747 10053
rect 10689 10044 10701 10047
rect 10652 10016 10701 10044
rect 10652 10004 10658 10016
rect 10689 10013 10701 10016
rect 10735 10013 10747 10047
rect 10796 10044 10824 10084
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 10796 10016 11989 10044
rect 10689 10007 10747 10013
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10013 13139 10047
rect 13081 10007 13139 10013
rect 13096 9976 13124 10007
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14752 10053 14780 10084
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 16132 10112 16160 10152
rect 16206 10140 16212 10192
rect 16264 10180 16270 10192
rect 18693 10183 18751 10189
rect 18693 10180 18705 10183
rect 16264 10152 18705 10180
rect 16264 10140 16270 10152
rect 18693 10149 18705 10152
rect 18739 10149 18751 10183
rect 18693 10143 18751 10149
rect 20993 10183 21051 10189
rect 20993 10149 21005 10183
rect 21039 10180 21051 10183
rect 21174 10180 21180 10192
rect 21039 10152 21180 10180
rect 21039 10149 21051 10152
rect 20993 10143 21051 10149
rect 21174 10140 21180 10152
rect 21232 10140 21238 10192
rect 24118 10140 24124 10192
rect 24176 10180 24182 10192
rect 24581 10183 24639 10189
rect 24581 10180 24593 10183
rect 24176 10152 24593 10180
rect 24176 10140 24182 10152
rect 24581 10149 24593 10152
rect 24627 10149 24639 10183
rect 24581 10143 24639 10149
rect 16482 10112 16488 10124
rect 16132 10084 16488 10112
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 17126 10072 17132 10124
rect 17184 10112 17190 10124
rect 20898 10112 20904 10124
rect 17184 10084 20904 10112
rect 17184 10072 17190 10084
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 21266 10072 21272 10124
rect 21324 10072 21330 10124
rect 25038 10072 25044 10124
rect 25096 10072 25102 10124
rect 25133 10115 25191 10121
rect 25133 10081 25145 10115
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 14056 10016 14105 10044
rect 14056 10004 14062 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10044 15899 10047
rect 16574 10044 16580 10056
rect 15887 10016 16580 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 16574 10004 16580 10016
rect 16632 10004 16638 10056
rect 16942 10004 16948 10056
rect 17000 10004 17006 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10044 17647 10047
rect 18049 10047 18107 10053
rect 18049 10044 18061 10047
rect 17635 10016 18061 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 18049 10013 18061 10016
rect 18095 10013 18107 10047
rect 19242 10044 19248 10056
rect 18049 10007 18107 10013
rect 19076 10016 19248 10044
rect 19076 9976 19104 10016
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10044 19763 10047
rect 20438 10044 20444 10056
rect 19751 10016 20444 10044
rect 19751 10013 19763 10016
rect 19705 10007 19763 10013
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 20714 10004 20720 10056
rect 20772 10004 20778 10056
rect 25148 10044 25176 10075
rect 23032 10016 25176 10044
rect 8496 9948 13032 9976
rect 13096 9948 19104 9976
rect 5074 9868 5080 9920
rect 5132 9908 5138 9920
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 5132 9880 7665 9908
rect 5132 9868 5138 9880
rect 7653 9877 7665 9880
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 8938 9908 8944 9920
rect 7800 9880 8944 9908
rect 7800 9868 7806 9880
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 11330 9868 11336 9920
rect 11388 9868 11394 9920
rect 13004 9908 13032 9948
rect 19150 9936 19156 9988
rect 19208 9976 19214 9988
rect 21545 9979 21603 9985
rect 21545 9976 21557 9979
rect 19208 9948 21557 9976
rect 19208 9936 19214 9948
rect 21545 9945 21557 9948
rect 21591 9945 21603 9979
rect 21545 9939 21603 9945
rect 21818 9936 21824 9988
rect 21876 9976 21882 9988
rect 21876 9948 22034 9976
rect 21876 9936 21882 9948
rect 13630 9908 13636 9920
rect 13004 9880 13636 9908
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 13722 9868 13728 9920
rect 13780 9868 13786 9920
rect 15381 9911 15439 9917
rect 15381 9877 15393 9911
rect 15427 9908 15439 9911
rect 17494 9908 17500 9920
rect 15427 9880 17500 9908
rect 15427 9877 15439 9880
rect 15381 9871 15439 9877
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 17862 9868 17868 9920
rect 17920 9908 17926 9920
rect 21726 9908 21732 9920
rect 17920 9880 21732 9908
rect 17920 9868 17926 9880
rect 21726 9868 21732 9880
rect 21784 9868 21790 9920
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 23032 9917 23060 10016
rect 23474 9936 23480 9988
rect 23532 9976 23538 9988
rect 23661 9979 23719 9985
rect 23661 9976 23673 9979
rect 23532 9948 23673 9976
rect 23532 9936 23538 9948
rect 23661 9945 23673 9948
rect 23707 9945 23719 9979
rect 23661 9939 23719 9945
rect 23017 9911 23075 9917
rect 23017 9908 23029 9911
rect 22980 9880 23029 9908
rect 22980 9868 22986 9880
rect 23017 9877 23029 9880
rect 23063 9877 23075 9911
rect 23017 9871 23075 9877
rect 23750 9868 23756 9920
rect 23808 9868 23814 9920
rect 24302 9868 24308 9920
rect 24360 9908 24366 9920
rect 24397 9911 24455 9917
rect 24397 9908 24409 9911
rect 24360 9880 24409 9908
rect 24360 9868 24366 9880
rect 24397 9877 24409 9880
rect 24443 9908 24455 9911
rect 24949 9911 25007 9917
rect 24949 9908 24961 9911
rect 24443 9880 24961 9908
rect 24443 9877 24455 9880
rect 24397 9871 24455 9877
rect 24949 9877 24961 9880
rect 24995 9877 25007 9911
rect 24949 9871 25007 9877
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 1118 9664 1124 9716
rect 1176 9704 1182 9716
rect 7742 9704 7748 9716
rect 1176 9676 7748 9704
rect 1176 9664 1182 9676
rect 7742 9664 7748 9676
rect 7800 9664 7806 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 14826 9704 14832 9716
rect 11848 9676 14832 9704
rect 11848 9664 11854 9676
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 14918 9664 14924 9716
rect 14976 9704 14982 9716
rect 14976 9676 15240 9704
rect 14976 9664 14982 9676
rect 4614 9636 4620 9648
rect 2976 9608 4620 9636
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 2314 9568 2320 9580
rect 1903 9540 2320 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2976 9577 3004 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 4706 9596 4712 9648
rect 4764 9596 4770 9648
rect 5166 9596 5172 9648
rect 5224 9596 5230 9648
rect 8294 9636 8300 9648
rect 5920 9608 8300 9636
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 5184 9568 5212 9596
rect 5920 9577 5948 9608
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 14090 9636 14096 9648
rect 9324 9608 14096 9636
rect 4295 9540 5212 9568
rect 5905 9571 5963 9577
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 5905 9537 5917 9571
rect 5951 9537 5963 9571
rect 5905 9531 5963 9537
rect 3620 9500 3648 9531
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 9324 9577 9352 9608
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 15212 9645 15240 9676
rect 16592 9676 18920 9704
rect 15197 9639 15255 9645
rect 15197 9605 15209 9639
rect 15243 9605 15255 9639
rect 16592 9636 16620 9676
rect 15197 9599 15255 9605
rect 15580 9608 16620 9636
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11848 9540 11897 9568
rect 11848 9528 11854 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 12342 9528 12348 9580
rect 12400 9528 12406 9580
rect 13449 9571 13507 9577
rect 13449 9537 13461 9571
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 14550 9568 14556 9580
rect 14507 9540 14556 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 3620 9472 5396 9500
rect 2130 9392 2136 9444
rect 2188 9392 2194 9444
rect 2777 9435 2835 9441
rect 2777 9401 2789 9435
rect 2823 9432 2835 9435
rect 2866 9432 2872 9444
rect 2823 9404 2872 9432
rect 2823 9401 2835 9404
rect 2777 9395 2835 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3421 9435 3479 9441
rect 3421 9401 3433 9435
rect 3467 9432 3479 9435
rect 3510 9432 3516 9444
rect 3467 9404 3516 9432
rect 3467 9401 3479 9404
rect 3421 9395 3479 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 5368 9376 5396 9472
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7432 9472 8033 9500
rect 7432 9460 7438 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9500 10379 9503
rect 10778 9500 10784 9512
rect 10367 9472 10784 9500
rect 10367 9469 10379 9472
rect 10321 9463 10379 9469
rect 5721 9435 5779 9441
rect 5721 9401 5733 9435
rect 5767 9432 5779 9435
rect 6362 9432 6368 9444
rect 5767 9404 6368 9432
rect 5767 9401 5779 9404
rect 5721 9395 5779 9401
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 9048 9432 9076 9463
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 13464 9500 13492 9531
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 14918 9528 14924 9580
rect 14976 9568 14982 9580
rect 15580 9568 15608 9608
rect 17678 9596 17684 9648
rect 17736 9636 17742 9648
rect 18785 9639 18843 9645
rect 18785 9636 18797 9639
rect 17736 9608 18797 9636
rect 17736 9596 17742 9608
rect 18785 9605 18797 9608
rect 18831 9605 18843 9639
rect 18785 9599 18843 9605
rect 14976 9540 15608 9568
rect 15657 9571 15715 9577
rect 14976 9528 14982 9540
rect 15657 9537 15669 9571
rect 15703 9568 15715 9571
rect 16298 9568 16304 9580
rect 15703 9540 16304 9568
rect 15703 9537 15715 9540
rect 15657 9531 15715 9537
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 16942 9500 16948 9512
rect 13464 9472 16948 9500
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17052 9500 17080 9531
rect 17218 9528 17224 9580
rect 17276 9568 17282 9580
rect 17862 9568 17868 9580
rect 17276 9540 17868 9568
rect 17276 9528 17282 9540
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 18012 9540 18153 9568
rect 18012 9528 18018 9540
rect 18141 9537 18153 9540
rect 18187 9537 18199 9571
rect 18141 9531 18199 9537
rect 18598 9500 18604 9512
rect 17052 9472 18604 9500
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 18892 9500 18920 9676
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 20162 9704 20168 9716
rect 19116 9676 20168 9704
rect 19116 9664 19122 9676
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 20438 9664 20444 9716
rect 20496 9664 20502 9716
rect 21174 9704 21180 9716
rect 20640 9676 21180 9704
rect 20640 9648 20668 9676
rect 21174 9664 21180 9676
rect 21232 9664 21238 9716
rect 20622 9636 20628 9648
rect 19306 9608 20628 9636
rect 19058 9528 19064 9580
rect 19116 9568 19122 9580
rect 19306 9568 19334 9608
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 23293 9639 23351 9645
rect 20916 9608 23060 9636
rect 19116 9540 19334 9568
rect 19797 9571 19855 9577
rect 19116 9528 19122 9540
rect 19797 9537 19809 9571
rect 19843 9568 19855 9571
rect 20806 9568 20812 9580
rect 19843 9540 20812 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 20916 9500 20944 9608
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9537 21051 9571
rect 20993 9531 21051 9537
rect 18892 9472 20944 9500
rect 11606 9432 11612 9444
rect 9048 9404 11612 9432
rect 11606 9392 11612 9404
rect 11664 9392 11670 9444
rect 11701 9435 11759 9441
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 11882 9432 11888 9444
rect 11747 9404 11888 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 14093 9435 14151 9441
rect 14093 9401 14105 9435
rect 14139 9432 14151 9435
rect 14139 9404 18000 9432
rect 14139 9401 14151 9404
rect 14093 9395 14151 9401
rect 566 9324 572 9376
rect 624 9364 630 9376
rect 3602 9364 3608 9376
rect 624 9336 3608 9364
rect 624 9324 630 9336
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 4062 9324 4068 9376
rect 4120 9324 4126 9376
rect 5350 9324 5356 9376
rect 5408 9324 5414 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 5500 9336 7021 9364
rect 5500 9324 5506 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 12158 9364 12164 9376
rect 7616 9336 12164 9364
rect 7616 9324 7622 9336
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 12768 9336 13001 9364
rect 12768 9324 12774 9336
rect 12989 9333 13001 9336
rect 13035 9333 13047 9367
rect 12989 9327 13047 9333
rect 16301 9367 16359 9373
rect 16301 9333 16313 9367
rect 16347 9364 16359 9367
rect 16574 9364 16580 9376
rect 16347 9336 16580 9364
rect 16347 9333 16359 9336
rect 16301 9327 16359 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 17126 9364 17132 9376
rect 16724 9336 17132 9364
rect 16724 9324 16730 9336
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 17368 9336 17693 9364
rect 17368 9324 17374 9336
rect 17681 9333 17693 9336
rect 17727 9333 17739 9367
rect 17972 9364 18000 9404
rect 18046 9392 18052 9444
rect 18104 9432 18110 9444
rect 21008 9432 21036 9531
rect 22186 9528 22192 9580
rect 22244 9528 22250 9580
rect 23032 9568 23060 9608
rect 23293 9605 23305 9639
rect 23339 9636 23351 9639
rect 24854 9636 24860 9648
rect 23339 9608 24860 9636
rect 23339 9605 23351 9608
rect 23293 9599 23351 9605
rect 24854 9596 24860 9608
rect 24912 9596 24918 9648
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23032 9540 23949 9568
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 22646 9460 22652 9512
rect 22704 9500 22710 9512
rect 22922 9500 22928 9512
rect 22704 9472 22928 9500
rect 22704 9460 22710 9472
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 18104 9404 21036 9432
rect 18104 9392 18110 9404
rect 21174 9392 21180 9444
rect 21232 9392 21238 9444
rect 18598 9364 18604 9376
rect 17972 9336 18604 9364
rect 17681 9327 17739 9333
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 19058 9324 19064 9376
rect 19116 9324 19122 9376
rect 20438 9324 20444 9376
rect 20496 9364 20502 9376
rect 20622 9364 20628 9376
rect 20496 9336 20628 9364
rect 20496 9324 20502 9336
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 21545 9367 21603 9373
rect 21545 9364 21557 9367
rect 20864 9336 21557 9364
rect 20864 9324 20870 9336
rect 21545 9333 21557 9336
rect 21591 9364 21603 9367
rect 23382 9364 23388 9376
rect 21591 9336 23388 9364
rect 21591 9333 21603 9336
rect 21545 9327 21603 9333
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 1578 9120 1584 9172
rect 1636 9120 1642 9172
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2498 9160 2504 9172
rect 1995 9132 2504 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3326 9160 3332 9172
rect 3283 9132 3332 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 3660 9132 5304 9160
rect 3660 9120 3666 9132
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 5169 9095 5227 9101
rect 5169 9092 5181 9095
rect 5132 9064 5181 9092
rect 5132 9052 5138 9064
rect 5169 9061 5181 9064
rect 5215 9061 5227 9095
rect 5276 9092 5304 9132
rect 5718 9120 5724 9172
rect 5776 9160 5782 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 5776 9132 5825 9160
rect 5776 9120 5782 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 7282 9120 7288 9172
rect 7340 9120 7346 9172
rect 7834 9120 7840 9172
rect 7892 9120 7898 9172
rect 7926 9120 7932 9172
rect 7984 9160 7990 9172
rect 8662 9160 8668 9172
rect 7984 9132 8668 9160
rect 7984 9120 7990 9132
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 8938 9120 8944 9172
rect 8996 9120 9002 9172
rect 11790 9160 11796 9172
rect 9048 9132 11796 9160
rect 9048 9092 9076 9132
rect 11790 9120 11796 9132
rect 11848 9160 11854 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 11848 9132 12357 9160
rect 11848 9120 11854 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13538 9160 13544 9172
rect 13320 9132 13544 9160
rect 13320 9120 13326 9132
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 16666 9160 16672 9172
rect 15160 9132 16672 9160
rect 15160 9120 15166 9132
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 16850 9120 16856 9172
rect 16908 9120 16914 9172
rect 17954 9120 17960 9172
rect 18012 9120 18018 9172
rect 19058 9160 19064 9172
rect 18524 9132 19064 9160
rect 5276 9064 9076 9092
rect 5169 9055 5227 9061
rect 9490 9052 9496 9104
rect 9548 9092 9554 9104
rect 14550 9092 14556 9104
rect 9548 9064 10180 9092
rect 9548 9052 9554 9064
rect 750 8984 756 9036
rect 808 9024 814 9036
rect 3602 9024 3608 9036
rect 808 8996 2774 9024
rect 808 8984 814 8996
rect 2746 8968 2774 8996
rect 3436 8996 3608 9024
rect 1578 8916 1584 8968
rect 1636 8956 1642 8968
rect 2133 8959 2191 8965
rect 2133 8956 2145 8959
rect 1636 8928 2145 8956
rect 1636 8916 1642 8928
rect 2133 8925 2145 8928
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2590 8916 2596 8968
rect 2648 8916 2654 8968
rect 2746 8928 2780 8968
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3436 8965 3464 8996
rect 3602 8984 3608 8996
rect 3660 9024 3666 9036
rect 4246 9024 4252 9036
rect 3660 8996 4252 9024
rect 3660 8984 3666 8996
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8956 4951 8959
rect 5092 8956 5120 9052
rect 7926 9024 7932 9036
rect 6012 8996 7932 9024
rect 6012 8965 6040 8996
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9309 9027 9367 9033
rect 9309 9024 9321 9027
rect 8536 8996 9321 9024
rect 8536 8984 8542 8996
rect 9309 8993 9321 8996
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 10152 9024 10180 9064
rect 11348 9064 14556 9092
rect 11348 9024 11376 9064
rect 14550 9052 14556 9064
rect 14608 9052 14614 9104
rect 10152 8996 11376 9024
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 9024 12127 9027
rect 12618 9024 12624 9036
rect 12115 8996 12624 9024
rect 12115 8993 12127 8996
rect 12069 8987 12127 8993
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 15378 8984 15384 9036
rect 15436 9024 15442 9036
rect 15436 8996 17448 9024
rect 15436 8984 15442 8996
rect 4939 8928 5120 8956
rect 5997 8959 6055 8965
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6733 8959 6791 8965
rect 6733 8956 6745 8959
rect 6328 8928 6745 8956
rect 6328 8916 6334 8928
rect 6733 8925 6745 8928
rect 6779 8956 6791 8959
rect 6822 8956 6828 8968
rect 6779 8928 6828 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 7834 8956 7840 8968
rect 7515 8928 7840 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 8573 8959 8631 8965
rect 8573 8952 8585 8959
rect 8496 8925 8585 8952
rect 8619 8925 8631 8959
rect 8496 8924 8631 8925
rect 2608 8888 2636 8916
rect 8021 8891 8079 8897
rect 8021 8888 8033 8891
rect 2608 8860 8033 8888
rect 8021 8857 8033 8860
rect 8067 8888 8079 8891
rect 8496 8888 8524 8924
rect 8573 8919 8631 8924
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 8720 8928 10088 8956
rect 8720 8916 8726 8928
rect 8067 8860 8524 8888
rect 8067 8857 8079 8860
rect 8021 8851 8079 8857
rect 2593 8823 2651 8829
rect 2593 8789 2605 8823
rect 2639 8820 2651 8823
rect 3878 8820 3884 8832
rect 2639 8792 3884 8820
rect 2639 8789 2651 8792
rect 2593 8783 2651 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 3970 8780 3976 8832
rect 4028 8780 4034 8832
rect 4706 8780 4712 8832
rect 4764 8780 4770 8832
rect 6546 8780 6552 8832
rect 6604 8780 6610 8832
rect 8389 8823 8447 8829
rect 8389 8789 8401 8823
rect 8435 8820 8447 8823
rect 8846 8820 8852 8832
rect 8435 8792 8852 8820
rect 8435 8789 8447 8792
rect 8389 8783 8447 8789
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 10060 8820 10088 8928
rect 11422 8916 11428 8968
rect 11480 8916 11486 8968
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 12216 8928 13093 8956
rect 12216 8916 12222 8928
rect 13081 8925 13093 8928
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 14366 8916 14372 8968
rect 14424 8916 14430 8968
rect 15102 8916 15108 8968
rect 15160 8916 15166 8968
rect 15654 8916 15660 8968
rect 15712 8956 15718 8968
rect 16209 8959 16267 8965
rect 16209 8956 16221 8959
rect 15712 8928 16221 8956
rect 15712 8916 15718 8928
rect 16209 8925 16221 8928
rect 16255 8925 16267 8959
rect 16209 8919 16267 8925
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 17218 8956 17224 8968
rect 16724 8928 17224 8956
rect 16724 8916 16730 8928
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17310 8916 17316 8968
rect 17368 8916 17374 8968
rect 17420 8956 17448 8996
rect 18417 8959 18475 8965
rect 17420 8928 18184 8956
rect 10318 8848 10324 8900
rect 10376 8848 10382 8900
rect 11606 8848 11612 8900
rect 11664 8888 11670 8900
rect 18046 8888 18052 8900
rect 11664 8860 18052 8888
rect 11664 8848 11670 8860
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 18156 8888 18184 8928
rect 18417 8925 18429 8959
rect 18463 8956 18475 8959
rect 18524 8956 18552 9132
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 19886 9120 19892 9172
rect 19944 9160 19950 9172
rect 21177 9163 21235 9169
rect 21177 9160 21189 9163
rect 19944 9132 21189 9160
rect 19944 9120 19950 9132
rect 21177 9129 21189 9132
rect 21223 9129 21235 9163
rect 22094 9160 22100 9172
rect 21177 9123 21235 9129
rect 22066 9120 22100 9160
rect 22152 9120 22158 9172
rect 25225 9163 25283 9169
rect 25225 9129 25237 9163
rect 25271 9160 25283 9163
rect 25774 9160 25780 9172
rect 25271 9132 25780 9160
rect 25271 9129 25283 9132
rect 25225 9123 25283 9129
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 18598 9052 18604 9104
rect 18656 9092 18662 9104
rect 22066 9092 22094 9120
rect 18656 9064 22094 9092
rect 18656 9052 18662 9064
rect 19058 8984 19064 9036
rect 19116 9024 19122 9036
rect 19116 8996 19564 9024
rect 19116 8984 19122 8996
rect 18463 8928 18552 8956
rect 18463 8925 18475 8928
rect 18417 8919 18475 8925
rect 18598 8916 18604 8968
rect 18656 8956 18662 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 18656 8928 19441 8956
rect 18656 8916 18662 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 18693 8891 18751 8897
rect 18693 8888 18705 8891
rect 18156 8860 18705 8888
rect 18693 8857 18705 8860
rect 18739 8857 18751 8891
rect 19536 8888 19564 8996
rect 19610 8984 19616 9036
rect 19668 9024 19674 9036
rect 19668 8996 22692 9024
rect 19668 8984 19674 8996
rect 22664 8965 22692 8996
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8956 20591 8959
rect 22649 8959 22707 8965
rect 20579 8928 22600 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 21729 8891 21787 8897
rect 21729 8888 21741 8891
rect 19536 8860 21741 8888
rect 18693 8851 18751 8857
rect 21729 8857 21741 8860
rect 21775 8888 21787 8891
rect 22189 8891 22247 8897
rect 22189 8888 22201 8891
rect 21775 8860 22201 8888
rect 21775 8857 21787 8860
rect 21729 8851 21787 8857
rect 22189 8857 22201 8860
rect 22235 8857 22247 8891
rect 22189 8851 22247 8857
rect 11698 8820 11704 8832
rect 10060 8792 11704 8820
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 13630 8780 13636 8832
rect 13688 8820 13694 8832
rect 13725 8823 13783 8829
rect 13725 8820 13737 8823
rect 13688 8792 13737 8820
rect 13688 8780 13694 8792
rect 13725 8789 13737 8792
rect 13771 8789 13783 8823
rect 13725 8783 13783 8789
rect 15746 8780 15752 8832
rect 15804 8780 15810 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 20073 8823 20131 8829
rect 20073 8820 20085 8823
rect 17644 8792 20085 8820
rect 17644 8780 17650 8792
rect 20073 8789 20085 8792
rect 20119 8789 20131 8823
rect 20073 8783 20131 8789
rect 21818 8780 21824 8832
rect 21876 8780 21882 8832
rect 22572 8820 22600 8928
rect 22649 8925 22661 8959
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 25222 8956 25228 8968
rect 24627 8928 25228 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 25222 8916 25228 8928
rect 25280 8916 25286 8968
rect 23845 8891 23903 8897
rect 23845 8857 23857 8891
rect 23891 8888 23903 8891
rect 24946 8888 24952 8900
rect 23891 8860 24952 8888
rect 23891 8857 23903 8860
rect 23845 8851 23903 8857
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 25590 8820 25596 8832
rect 22572 8792 25596 8820
rect 25590 8780 25596 8792
rect 25648 8780 25654 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 1949 8619 2007 8625
rect 1949 8585 1961 8619
rect 1995 8616 2007 8619
rect 2222 8616 2228 8628
rect 1995 8588 2228 8616
rect 1995 8585 2007 8588
rect 1949 8579 2007 8585
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 2590 8576 2596 8628
rect 2648 8576 2654 8628
rect 3234 8576 3240 8628
rect 3292 8576 3298 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4212 8588 4445 8616
rect 4212 8576 4218 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 6822 8576 6828 8628
rect 6880 8576 6886 8628
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 8665 8619 8723 8625
rect 8665 8616 8677 8619
rect 8444 8588 8677 8616
rect 8444 8576 8450 8588
rect 8665 8585 8677 8588
rect 8711 8585 8723 8619
rect 8665 8579 8723 8585
rect 9674 8576 9680 8628
rect 9732 8576 9738 8628
rect 15102 8616 15108 8628
rect 10152 8588 15108 8616
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 9030 8548 9036 8560
rect 4028 8520 9036 8548
rect 4028 8508 4034 8520
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4212 8452 4629 8480
rect 4212 8440 4218 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8812 8452 8861 8480
rect 8812 8440 8818 8452
rect 8849 8449 8861 8452
rect 8895 8480 8907 8483
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 8895 8452 9137 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9125 8449 9137 8452
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9447 8452 9873 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9861 8449 9873 8452
rect 9907 8480 9919 8483
rect 10042 8480 10048 8492
rect 9907 8452 10048 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 10152 8412 10180 8588
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 16758 8616 16764 8628
rect 15243 8588 16764 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 18598 8576 18604 8628
rect 18656 8576 18662 8628
rect 20809 8619 20867 8625
rect 20809 8585 20821 8619
rect 20855 8616 20867 8619
rect 20990 8616 20996 8628
rect 20855 8588 20996 8616
rect 20855 8585 20867 8588
rect 20809 8579 20867 8585
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 19610 8548 19616 8560
rect 12124 8520 15700 8548
rect 12124 8508 12130 8520
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 13262 8480 13268 8492
rect 12023 8452 13268 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 14274 8480 14280 8492
rect 13495 8452 14280 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14550 8440 14556 8492
rect 14608 8440 14614 8492
rect 15672 8489 15700 8520
rect 16776 8520 19616 8548
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 16666 8480 16672 8492
rect 15657 8443 15715 8449
rect 16224 8452 16672 8480
rect 4856 8384 10180 8412
rect 10321 8415 10379 8421
rect 4856 8372 4862 8384
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10502 8412 10508 8424
rect 10367 8384 10508 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 11698 8372 11704 8424
rect 11756 8372 11762 8424
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 16224 8412 16252 8452
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 12676 8384 16252 8412
rect 12676 8372 12682 8384
rect 16298 8372 16304 8424
rect 16356 8372 16362 8424
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 3973 8347 4031 8353
rect 3973 8344 3985 8347
rect 3844 8316 3985 8344
rect 3844 8304 3850 8316
rect 3973 8313 3985 8316
rect 4019 8313 4031 8347
rect 3973 8307 4031 8313
rect 14093 8347 14151 8353
rect 14093 8313 14105 8347
rect 14139 8344 14151 8347
rect 14826 8344 14832 8356
rect 14139 8316 14832 8344
rect 14139 8313 14151 8316
rect 14093 8307 14151 8313
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 13814 8276 13820 8288
rect 11204 8248 13820 8276
rect 11204 8236 11210 8248
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 16776 8276 16804 8520
rect 19610 8508 19616 8520
rect 19668 8508 19674 8560
rect 19794 8508 19800 8560
rect 19852 8548 19858 8560
rect 21269 8551 21327 8557
rect 21269 8548 21281 8551
rect 19852 8520 21281 8548
rect 19852 8508 19858 8520
rect 21269 8517 21281 8520
rect 21315 8517 21327 8551
rect 21269 8511 21327 8517
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 16868 8344 16896 8443
rect 17954 8440 17960 8492
rect 18012 8440 18018 8492
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 19061 8483 19119 8489
rect 19061 8480 19073 8483
rect 18840 8452 19073 8480
rect 18840 8440 18846 8452
rect 19061 8449 19073 8452
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 20070 8440 20076 8492
rect 20128 8480 20134 8492
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 20128 8452 20177 8480
rect 20128 8440 20134 8452
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 22094 8440 22100 8492
rect 22152 8440 22158 8492
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 17310 8372 17316 8424
rect 17368 8412 17374 8424
rect 17497 8415 17555 8421
rect 17497 8412 17509 8415
rect 17368 8384 17509 8412
rect 17368 8372 17374 8384
rect 17497 8381 17509 8384
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 17586 8372 17592 8424
rect 17644 8412 17650 8424
rect 18874 8412 18880 8424
rect 17644 8384 18880 8412
rect 17644 8372 17650 8384
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 22002 8412 22008 8424
rect 19392 8384 22008 8412
rect 19392 8372 19398 8384
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 23382 8412 23388 8424
rect 23339 8384 23388 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 23382 8372 23388 8384
rect 23440 8372 23446 8424
rect 24210 8344 24216 8356
rect 16868 8316 24216 8344
rect 24210 8304 24216 8316
rect 24268 8304 24274 8356
rect 15896 8248 16804 8276
rect 15896 8236 15902 8248
rect 16850 8236 16856 8288
rect 16908 8276 16914 8288
rect 19058 8276 19064 8288
rect 16908 8248 19064 8276
rect 16908 8236 16914 8248
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 19705 8279 19763 8285
rect 19705 8276 19717 8279
rect 19484 8248 19717 8276
rect 19484 8236 19490 8248
rect 19705 8245 19717 8248
rect 19751 8245 19763 8279
rect 19705 8239 19763 8245
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 2004 8044 2145 8072
rect 2004 8032 2010 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2133 8035 2191 8041
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2869 8075 2927 8081
rect 2869 8072 2881 8075
rect 2832 8044 2881 8072
rect 2832 8032 2838 8044
rect 2869 8041 2881 8044
rect 2915 8041 2927 8075
rect 2869 8035 2927 8041
rect 3602 8032 3608 8084
rect 3660 8032 3666 8084
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 10505 8075 10563 8081
rect 10505 8072 10517 8075
rect 10376 8044 10517 8072
rect 10376 8032 10382 8044
rect 10505 8041 10517 8044
rect 10551 8041 10563 8075
rect 10505 8035 10563 8041
rect 12158 8032 12164 8084
rect 12216 8072 12222 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 12216 8044 12357 8072
rect 12216 8032 12222 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12584 8044 12909 8072
rect 12584 8032 12590 8044
rect 12897 8041 12909 8044
rect 12943 8072 12955 8075
rect 13906 8072 13912 8084
rect 12943 8044 13912 8072
rect 12943 8041 12955 8044
rect 12897 8035 12955 8041
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 14185 8075 14243 8081
rect 14185 8041 14197 8075
rect 14231 8072 14243 8075
rect 14274 8072 14280 8084
rect 14231 8044 14280 8072
rect 14231 8041 14243 8044
rect 14185 8035 14243 8041
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 16850 8072 16856 8084
rect 14476 8044 16856 8072
rect 2590 7964 2596 8016
rect 2648 7964 2654 8016
rect 3878 7964 3884 8016
rect 3936 8004 3942 8016
rect 14476 8004 14504 8044
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 17000 8044 17325 8072
rect 17000 8032 17006 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18417 8075 18475 8081
rect 18417 8072 18429 8075
rect 18012 8044 18429 8072
rect 18012 8032 18018 8044
rect 18417 8041 18429 8044
rect 18463 8041 18475 8075
rect 18417 8035 18475 8041
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 19150 8072 19156 8084
rect 18932 8044 19156 8072
rect 18932 8032 18938 8044
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 20070 8032 20076 8084
rect 20128 8032 20134 8084
rect 3936 7976 14504 8004
rect 3936 7964 3942 7976
rect 15102 7964 15108 8016
rect 15160 7964 15166 8016
rect 22186 8004 22192 8016
rect 17236 7976 22192 8004
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 17236 7936 17264 7976
rect 22186 7964 22192 7976
rect 22244 7964 22250 8016
rect 11287 7908 17264 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 20714 7896 20720 7948
rect 20772 7936 20778 7948
rect 20809 7939 20867 7945
rect 20809 7936 20821 7939
rect 20772 7908 20821 7936
rect 20772 7896 20778 7908
rect 20809 7905 20821 7908
rect 20855 7905 20867 7939
rect 23658 7936 23664 7948
rect 20809 7899 20867 7905
rect 20916 7908 23664 7936
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2590 7868 2596 7880
rect 2363 7840 2596 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13495 7840 13737 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 13725 7837 13737 7840
rect 13771 7868 13783 7871
rect 13998 7868 14004 7880
rect 13771 7840 14004 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7868 14519 7871
rect 15194 7868 15200 7880
rect 14507 7840 15200 7868
rect 14507 7837 14519 7840
rect 14461 7831 14519 7837
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7868 15623 7871
rect 16390 7868 16396 7880
rect 15611 7840 16396 7868
rect 15611 7837 15623 7840
rect 15565 7831 15623 7837
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7837 16727 7871
rect 16669 7831 16727 7837
rect 6546 7760 6552 7812
rect 6604 7800 6610 7812
rect 11606 7800 11612 7812
rect 6604 7772 11612 7800
rect 6604 7760 6610 7772
rect 11606 7760 11612 7772
rect 11664 7760 11670 7812
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 16684 7800 16712 7831
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 17460 7840 17785 7868
rect 17460 7828 17466 7840
rect 17773 7837 17785 7840
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 19426 7828 19432 7880
rect 19484 7828 19490 7880
rect 20438 7828 20444 7880
rect 20496 7868 20502 7880
rect 20625 7871 20683 7877
rect 20625 7868 20637 7871
rect 20496 7840 20637 7868
rect 20496 7828 20502 7840
rect 20625 7837 20637 7840
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 13872 7772 16712 7800
rect 13872 7760 13878 7772
rect 16758 7760 16764 7812
rect 16816 7800 16822 7812
rect 20916 7800 20944 7908
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 26234 7936 26240 7948
rect 23768 7908 26240 7936
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 22370 7868 22376 7880
rect 21591 7840 22376 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 22370 7828 22376 7840
rect 22428 7828 22434 7880
rect 22830 7828 22836 7880
rect 22888 7828 22894 7880
rect 23768 7800 23796 7908
rect 26234 7896 26240 7908
rect 26292 7896 26298 7948
rect 24394 7828 24400 7880
rect 24452 7868 24458 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24452 7840 24593 7868
rect 24452 7828 24458 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 16816 7772 20944 7800
rect 22066 7772 23796 7800
rect 23845 7803 23903 7809
rect 16816 7760 16822 7772
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 11330 7732 11336 7744
rect 1728 7704 11336 7732
rect 1728 7692 1734 7704
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 13722 7732 13728 7744
rect 13587 7704 13728 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 16206 7692 16212 7744
rect 16264 7692 16270 7744
rect 16666 7692 16672 7744
rect 16724 7732 16730 7744
rect 22066 7732 22094 7772
rect 23845 7769 23857 7803
rect 23891 7800 23903 7803
rect 24946 7800 24952 7812
rect 23891 7772 24952 7800
rect 23891 7769 23903 7772
rect 23845 7763 23903 7769
rect 24946 7760 24952 7772
rect 25004 7760 25010 7812
rect 16724 7704 22094 7732
rect 16724 7692 16730 7704
rect 22186 7692 22192 7744
rect 22244 7692 22250 7744
rect 25222 7692 25228 7744
rect 25280 7692 25286 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 10965 7531 11023 7537
rect 10965 7528 10977 7531
rect 10560 7500 10977 7528
rect 10560 7488 10566 7500
rect 10965 7497 10977 7500
rect 11011 7497 11023 7531
rect 10965 7491 11023 7497
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 12250 7528 12256 7540
rect 11839 7500 12256 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 15010 7488 15016 7540
rect 15068 7488 15074 7540
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 15930 7528 15936 7540
rect 15252 7500 15936 7528
rect 15252 7488 15258 7500
rect 15930 7488 15936 7500
rect 15988 7528 15994 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 15988 7500 16129 7528
rect 15988 7488 15994 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16117 7491 16175 7497
rect 16390 7488 16396 7540
rect 16448 7488 16454 7540
rect 17402 7488 17408 7540
rect 17460 7528 17466 7540
rect 18506 7528 18512 7540
rect 17460 7500 18512 7528
rect 17460 7488 17466 7500
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 18785 7531 18843 7537
rect 18785 7497 18797 7531
rect 18831 7528 18843 7531
rect 23842 7528 23848 7540
rect 18831 7500 23848 7528
rect 18831 7497 18843 7500
rect 18785 7491 18843 7497
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 6236 7432 12572 7460
rect 6236 7420 6242 7432
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 6788 7364 10517 7392
rect 6788 7352 6794 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7392 10931 7395
rect 11146 7392 11152 7404
rect 10919 7364 11152 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 12544 7392 12572 7432
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 12952 7432 15884 7460
rect 12952 7420 12958 7432
rect 12713 7395 12771 7401
rect 12544 7364 12664 7392
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12526 7324 12532 7336
rect 12483 7296 12532 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 12636 7324 12664 7364
rect 12713 7361 12725 7395
rect 12759 7392 12771 7395
rect 14001 7395 14059 7401
rect 12759 7364 13952 7392
rect 12759 7361 12771 7364
rect 12713 7355 12771 7361
rect 12894 7324 12900 7336
rect 12636 7296 12900 7324
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 13814 7324 13820 7336
rect 13771 7296 13820 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 13924 7324 13952 7364
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14642 7392 14648 7404
rect 14047 7364 14648 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 15194 7352 15200 7404
rect 15252 7352 15258 7404
rect 15856 7401 15884 7432
rect 16574 7420 16580 7472
rect 16632 7460 16638 7472
rect 19889 7463 19947 7469
rect 16632 7432 19380 7460
rect 16632 7420 16638 7432
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 18138 7352 18144 7404
rect 18196 7352 18202 7404
rect 19242 7352 19248 7404
rect 19300 7352 19306 7404
rect 19352 7392 19380 7432
rect 19889 7429 19901 7463
rect 19935 7460 19947 7463
rect 25866 7460 25872 7472
rect 19935 7432 25872 7460
rect 19935 7429 19947 7432
rect 19889 7423 19947 7429
rect 25866 7420 25872 7432
rect 25924 7420 25930 7472
rect 20349 7395 20407 7401
rect 20349 7392 20361 7395
rect 19352 7364 20361 7392
rect 20349 7361 20361 7364
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 20438 7352 20444 7404
rect 20496 7392 20502 7404
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 20496 7364 21281 7392
rect 20496 7352 20502 7364
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 16758 7324 16764 7336
rect 13924 7296 16764 7324
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 16850 7284 16856 7336
rect 16908 7284 16914 7336
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7293 17187 7327
rect 17129 7287 17187 7293
rect 4522 7216 4528 7268
rect 4580 7256 4586 7268
rect 16206 7256 16212 7268
rect 4580 7228 16212 7256
rect 4580 7216 4586 7228
rect 16206 7216 16212 7228
rect 16264 7216 16270 7268
rect 17144 7256 17172 7287
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 22112 7324 22140 7355
rect 23934 7352 23940 7404
rect 23992 7352 23998 7404
rect 24670 7352 24676 7404
rect 24728 7392 24734 7404
rect 24728 7364 24808 7392
rect 24728 7352 24734 7364
rect 18104 7296 22140 7324
rect 18104 7284 18110 7296
rect 23290 7284 23296 7336
rect 23348 7284 23354 7336
rect 24780 7333 24808 7364
rect 24765 7327 24823 7333
rect 24765 7293 24777 7327
rect 24811 7293 24823 7327
rect 24765 7287 24823 7293
rect 22738 7256 22744 7268
rect 17144 7228 22744 7256
rect 22738 7216 22744 7228
rect 22796 7216 22802 7268
rect 10318 7148 10324 7200
rect 10376 7148 10382 7200
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 12308 7160 15669 7188
rect 12308 7148 12314 7160
rect 15657 7157 15669 7160
rect 15703 7157 15715 7191
rect 15657 7151 15715 7157
rect 20714 7148 20720 7200
rect 20772 7188 20778 7200
rect 20993 7191 21051 7197
rect 20993 7188 21005 7191
rect 20772 7160 21005 7188
rect 20772 7148 20778 7160
rect 20993 7157 21005 7160
rect 21039 7157 21051 7191
rect 20993 7151 21051 7157
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 12618 6944 12624 6996
rect 12676 6993 12682 6996
rect 12676 6987 12725 6993
rect 12676 6953 12679 6987
rect 12713 6953 12725 6987
rect 12676 6947 12725 6953
rect 12676 6944 12682 6947
rect 14550 6944 14556 6996
rect 14608 6984 14614 6996
rect 18046 6984 18052 6996
rect 14608 6956 18052 6984
rect 14608 6944 14614 6956
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 18877 6987 18935 6993
rect 18877 6984 18889 6987
rect 18196 6956 18889 6984
rect 18196 6944 18202 6956
rect 18877 6953 18889 6956
rect 18923 6953 18935 6987
rect 26786 6984 26792 6996
rect 18877 6947 18935 6953
rect 18984 6956 26792 6984
rect 15194 6876 15200 6928
rect 15252 6916 15258 6928
rect 16761 6919 16819 6925
rect 16761 6916 16773 6919
rect 15252 6888 16773 6916
rect 15252 6876 15258 6888
rect 16761 6885 16773 6888
rect 16807 6916 16819 6919
rect 18984 6916 19012 6956
rect 26786 6944 26792 6956
rect 26844 6944 26850 6996
rect 16807 6888 19012 6916
rect 16807 6885 16819 6888
rect 16761 6879 16819 6885
rect 19242 6876 19248 6928
rect 19300 6876 19306 6928
rect 22002 6876 22008 6928
rect 22060 6916 22066 6928
rect 22060 6888 22324 6916
rect 22060 6876 22066 6888
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 10134 6848 10140 6860
rect 5408 6820 10140 6848
rect 5408 6808 5414 6820
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 11624 6820 17172 6848
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 11333 6783 11391 6789
rect 11333 6780 11345 6783
rect 1452 6752 11345 6780
rect 1452 6740 1458 6752
rect 11333 6749 11345 6752
rect 11379 6780 11391 6783
rect 11514 6780 11520 6792
rect 11379 6752 11520 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 3418 6672 3424 6724
rect 3476 6712 3482 6724
rect 8294 6712 8300 6724
rect 3476 6684 8300 6712
rect 3476 6672 3482 6684
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 9582 6672 9588 6724
rect 9640 6712 9646 6724
rect 11624 6712 11652 6820
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 12544 6752 12848 6780
rect 12544 6712 12572 6752
rect 9640 6684 11652 6712
rect 11808 6684 12572 6712
rect 12820 6712 12848 6752
rect 13262 6740 13268 6792
rect 13320 6780 13326 6792
rect 14921 6783 14979 6789
rect 13320 6752 14872 6780
rect 13320 6740 13326 6752
rect 13446 6712 13452 6724
rect 12820 6684 13452 6712
rect 9640 6672 9646 6684
rect 11146 6604 11152 6656
rect 11204 6604 11210 6656
rect 11808 6653 11836 6684
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 14844 6712 14872 6752
rect 14921 6749 14933 6783
rect 14967 6780 14979 6783
rect 15102 6780 15108 6792
rect 14967 6752 15108 6780
rect 14967 6749 14979 6752
rect 14921 6743 14979 6749
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 15565 6783 15623 6789
rect 15565 6749 15577 6783
rect 15611 6780 15623 6783
rect 15930 6780 15936 6792
rect 15611 6752 15936 6780
rect 15611 6749 15623 6752
rect 15565 6743 15623 6749
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16206 6740 16212 6792
rect 16264 6740 16270 6792
rect 16574 6740 16580 6792
rect 16632 6740 16638 6792
rect 17144 6789 17172 6820
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 19150 6848 19156 6860
rect 17552 6820 19156 6848
rect 17552 6808 17558 6820
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 20346 6808 20352 6860
rect 20404 6808 20410 6860
rect 22186 6848 22192 6860
rect 20824 6820 22192 6848
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17276 6752 18245 6780
rect 17276 6740 17282 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6780 19763 6783
rect 20714 6780 20720 6792
rect 19751 6752 20720 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 20714 6740 20720 6752
rect 20772 6740 20778 6792
rect 20824 6789 20852 6820
rect 22186 6808 22192 6820
rect 22244 6808 22250 6860
rect 22296 6848 22324 6888
rect 22554 6848 22560 6860
rect 22296 6820 22560 6848
rect 22554 6808 22560 6820
rect 22612 6808 22618 6860
rect 20809 6783 20867 6789
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 22097 6783 22155 6789
rect 22097 6749 22109 6783
rect 22143 6780 22155 6783
rect 22278 6780 22284 6792
rect 22143 6752 22284 6780
rect 22143 6749 22155 6752
rect 22097 6743 22155 6749
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 25222 6780 25228 6792
rect 24627 6752 25228 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 13556 6684 14780 6712
rect 14844 6684 17785 6712
rect 11701 6647 11759 6653
rect 11701 6613 11713 6647
rect 11747 6644 11759 6647
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11747 6616 11805 6644
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 13556 6644 13584 6684
rect 11940 6616 13584 6644
rect 11940 6604 11946 6616
rect 14458 6604 14464 6656
rect 14516 6604 14522 6656
rect 14752 6653 14780 6684
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 22664 6712 22692 6743
rect 25222 6740 25228 6752
rect 25280 6740 25286 6792
rect 17773 6675 17831 6681
rect 17880 6684 22692 6712
rect 23845 6715 23903 6721
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6613 14795 6647
rect 14737 6607 14795 6613
rect 15378 6604 15384 6656
rect 15436 6604 15442 6656
rect 16022 6604 16028 6656
rect 16080 6604 16086 6656
rect 16758 6604 16764 6656
rect 16816 6644 16822 6656
rect 17880 6644 17908 6684
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 25682 6712 25688 6724
rect 23891 6684 25688 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 25682 6672 25688 6684
rect 25740 6672 25746 6724
rect 16816 6616 17908 6644
rect 16816 6604 16822 6616
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 21453 6647 21511 6653
rect 21453 6644 21465 6647
rect 20036 6616 21465 6644
rect 20036 6604 20042 6616
rect 21453 6613 21465 6616
rect 21499 6613 21511 6647
rect 21453 6607 21511 6613
rect 21542 6604 21548 6656
rect 21600 6644 21606 6656
rect 21913 6647 21971 6653
rect 21913 6644 21925 6647
rect 21600 6616 21925 6644
rect 21600 6604 21606 6616
rect 21913 6613 21925 6616
rect 21959 6613 21971 6647
rect 21913 6607 21971 6613
rect 25038 6604 25044 6656
rect 25096 6644 25102 6656
rect 25225 6647 25283 6653
rect 25225 6644 25237 6647
rect 25096 6616 25237 6644
rect 25096 6604 25102 6616
rect 25225 6613 25237 6616
rect 25271 6613 25283 6647
rect 25225 6607 25283 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9858 6440 9864 6452
rect 9355 6412 9864 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 11514 6400 11520 6452
rect 11572 6400 11578 6452
rect 12894 6400 12900 6452
rect 12952 6400 12958 6452
rect 14458 6400 14464 6452
rect 14516 6440 14522 6452
rect 15102 6440 15108 6452
rect 14516 6412 15108 6440
rect 14516 6400 14522 6412
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 15470 6400 15476 6452
rect 15528 6400 15534 6452
rect 16025 6443 16083 6449
rect 16025 6409 16037 6443
rect 16071 6440 16083 6443
rect 16114 6440 16120 6452
rect 16071 6412 16120 6440
rect 16071 6409 16083 6412
rect 16025 6403 16083 6409
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 16945 6443 17003 6449
rect 16945 6409 16957 6443
rect 16991 6440 17003 6443
rect 22002 6440 22008 6452
rect 16991 6412 22008 6440
rect 16991 6409 17003 6412
rect 16945 6403 17003 6409
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 11882 6372 11888 6384
rect 7708 6344 11888 6372
rect 7708 6332 7714 6344
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 12710 6332 12716 6384
rect 12768 6372 12774 6384
rect 12768 6344 15608 6372
rect 12768 6332 12774 6344
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 12268 6276 12940 6304
rect 12268 6245 12296 6276
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 12253 6239 12311 6245
rect 12253 6236 12265 6239
rect 12207 6208 12265 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12253 6205 12265 6208
rect 12299 6205 12311 6239
rect 12912 6236 12940 6276
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13412 6276 13737 6304
rect 13412 6264 13418 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 14182 6264 14188 6316
rect 14240 6264 14246 6316
rect 15286 6304 15292 6316
rect 14292 6276 15292 6304
rect 14292 6236 14320 6276
rect 15286 6264 15292 6276
rect 15344 6264 15350 6316
rect 12253 6199 12311 6205
rect 12406 6208 12848 6236
rect 12912 6208 14320 6236
rect 14461 6239 14519 6245
rect 11974 6128 11980 6180
rect 12032 6168 12038 6180
rect 12406 6168 12434 6208
rect 12032 6140 12434 6168
rect 12820 6168 12848 6208
rect 14461 6205 14473 6239
rect 14507 6236 14519 6239
rect 14918 6236 14924 6248
rect 14507 6208 14924 6236
rect 14507 6205 14519 6208
rect 14461 6199 14519 6205
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 15580 6236 15608 6344
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6304 15715 6307
rect 16960 6304 16988 6403
rect 22002 6400 22008 6412
rect 22060 6400 22066 6452
rect 22370 6400 22376 6452
rect 22428 6440 22434 6452
rect 22649 6443 22707 6449
rect 22649 6440 22661 6443
rect 22428 6412 22661 6440
rect 22428 6400 22434 6412
rect 22649 6409 22661 6412
rect 22695 6409 22707 6443
rect 22649 6403 22707 6409
rect 17034 6332 17040 6384
rect 17092 6372 17098 6384
rect 18690 6372 18696 6384
rect 17092 6344 18696 6372
rect 17092 6332 17098 6344
rect 18690 6332 18696 6344
rect 18748 6332 18754 6384
rect 18874 6332 18880 6384
rect 18932 6372 18938 6384
rect 19153 6375 19211 6381
rect 19153 6372 19165 6375
rect 18932 6344 19165 6372
rect 18932 6332 18938 6344
rect 19153 6341 19165 6344
rect 19199 6341 19211 6375
rect 19153 6335 19211 6341
rect 19889 6375 19947 6381
rect 19889 6341 19901 6375
rect 19935 6372 19947 6375
rect 23474 6372 23480 6384
rect 19935 6344 23480 6372
rect 19935 6341 19947 6344
rect 19889 6335 19947 6341
rect 23474 6332 23480 6344
rect 23532 6332 23538 6384
rect 24026 6372 24032 6384
rect 23584 6344 24032 6372
rect 15703 6276 16988 6304
rect 17405 6307 17463 6313
rect 15703 6273 15715 6276
rect 15657 6267 15715 6273
rect 17405 6273 17417 6307
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17218 6236 17224 6248
rect 15580 6208 17224 6236
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 17420 6236 17448 6267
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 17828 6276 18061 6304
rect 17828 6264 17834 6276
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6304 18567 6307
rect 19610 6304 19616 6316
rect 18555 6276 19616 6304
rect 18555 6273 18567 6276
rect 18509 6267 18567 6273
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 19702 6264 19708 6316
rect 19760 6264 19766 6316
rect 20806 6264 20812 6316
rect 20864 6264 20870 6316
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6304 22063 6307
rect 23584 6304 23612 6344
rect 24026 6332 24032 6344
rect 24084 6332 24090 6384
rect 22051 6276 23612 6304
rect 22051 6273 22063 6276
rect 22005 6267 22063 6273
rect 23934 6264 23940 6316
rect 23992 6264 23998 6316
rect 19886 6236 19892 6248
rect 17420 6208 19892 6236
rect 19886 6196 19892 6208
rect 19944 6196 19950 6248
rect 19978 6196 19984 6248
rect 20036 6236 20042 6248
rect 20165 6239 20223 6245
rect 20165 6236 20177 6239
rect 20036 6208 20177 6236
rect 20036 6196 20042 6208
rect 20165 6205 20177 6208
rect 20211 6236 20223 6239
rect 20533 6239 20591 6245
rect 20533 6236 20545 6239
rect 20211 6208 20545 6236
rect 20211 6205 20223 6208
rect 20165 6199 20223 6205
rect 20533 6205 20545 6208
rect 20579 6205 20591 6239
rect 20533 6199 20591 6205
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 23569 6171 23627 6177
rect 23569 6168 23581 6171
rect 12820 6140 23581 6168
rect 12032 6128 12038 6140
rect 23569 6137 23581 6140
rect 23615 6168 23627 6171
rect 23934 6168 23940 6180
rect 23615 6140 23940 6168
rect 23615 6137 23627 6140
rect 23569 6131 23627 6137
rect 23934 6128 23940 6140
rect 23992 6128 23998 6180
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 13262 6100 13268 6112
rect 9364 6072 13268 6100
rect 9364 6060 9370 6072
rect 13262 6060 13268 6072
rect 13320 6060 13326 6112
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 16761 6103 16819 6109
rect 16761 6100 16773 6103
rect 15988 6072 16773 6100
rect 15988 6060 15994 6072
rect 16761 6069 16773 6072
rect 16807 6100 16819 6103
rect 17586 6100 17592 6112
rect 16807 6072 17592 6100
rect 16807 6069 16819 6072
rect 16761 6063 16819 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 18230 6060 18236 6112
rect 18288 6100 18294 6112
rect 18598 6100 18604 6112
rect 18288 6072 18604 6100
rect 18288 6060 18294 6072
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 19978 6060 19984 6112
rect 20036 6100 20042 6112
rect 21634 6100 21640 6112
rect 20036 6072 21640 6100
rect 20036 6060 20042 6072
rect 21634 6060 21640 6072
rect 21692 6060 21698 6112
rect 22830 6060 22836 6112
rect 22888 6100 22894 6112
rect 22925 6103 22983 6109
rect 22925 6100 22937 6103
rect 22888 6072 22937 6100
rect 22888 6060 22894 6072
rect 22925 6069 22937 6072
rect 22971 6069 22983 6103
rect 22925 6063 22983 6069
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 10594 5856 10600 5908
rect 10652 5896 10658 5908
rect 16758 5896 16764 5908
rect 10652 5868 16764 5896
rect 10652 5856 10658 5868
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 16853 5899 16911 5905
rect 16853 5865 16865 5899
rect 16899 5896 16911 5899
rect 16942 5896 16948 5908
rect 16899 5868 16948 5896
rect 16899 5865 16911 5868
rect 16853 5859 16911 5865
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 18414 5856 18420 5908
rect 18472 5896 18478 5908
rect 18472 5868 21680 5896
rect 18472 5856 18478 5868
rect 5626 5788 5632 5840
rect 5684 5828 5690 5840
rect 21542 5828 21548 5840
rect 5684 5800 21548 5828
rect 5684 5788 5690 5800
rect 21542 5788 21548 5800
rect 21600 5788 21606 5840
rect 10226 5720 10232 5772
rect 10284 5760 10290 5772
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 10284 5732 20269 5760
rect 10284 5720 10290 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 21358 5720 21364 5772
rect 21416 5720 21422 5772
rect 21652 5769 21680 5868
rect 21637 5763 21695 5769
rect 21637 5729 21649 5763
rect 21683 5729 21695 5763
rect 21637 5723 21695 5729
rect 21744 5732 24624 5760
rect 13722 5652 13728 5704
rect 13780 5652 13786 5704
rect 14274 5652 14280 5704
rect 14332 5652 14338 5704
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 13740 5624 13768 5652
rect 15580 5624 15608 5655
rect 15838 5652 15844 5704
rect 15896 5652 15902 5704
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5692 17095 5695
rect 17126 5692 17132 5704
rect 17083 5664 17132 5692
rect 17083 5661 17095 5664
rect 17037 5655 17095 5661
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 19613 5695 19671 5701
rect 19613 5692 19625 5695
rect 18432 5664 19625 5692
rect 13740 5596 15608 5624
rect 17586 5584 17592 5636
rect 17644 5584 17650 5636
rect 17770 5584 17776 5636
rect 17828 5584 17834 5636
rect 12897 5559 12955 5565
rect 12897 5525 12909 5559
rect 12943 5556 12955 5559
rect 13354 5556 13360 5568
rect 12943 5528 13360 5556
rect 12943 5525 12955 5528
rect 12897 5519 12955 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13722 5556 13728 5568
rect 13587 5528 13728 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 15746 5516 15752 5568
rect 15804 5556 15810 5568
rect 18432 5556 18460 5664
rect 19613 5661 19625 5664
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 20898 5652 20904 5704
rect 20956 5652 20962 5704
rect 18874 5584 18880 5636
rect 18932 5584 18938 5636
rect 19150 5584 19156 5636
rect 19208 5624 19214 5636
rect 21744 5624 21772 5732
rect 24596 5701 24624 5732
rect 22649 5695 22707 5701
rect 22649 5692 22661 5695
rect 19208 5596 21772 5624
rect 22066 5664 22661 5692
rect 19208 5584 19214 5596
rect 15804 5528 18460 5556
rect 15804 5516 15810 5528
rect 18598 5516 18604 5568
rect 18656 5556 18662 5568
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 18656 5528 19257 5556
rect 18656 5516 18662 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 19245 5519 19303 5525
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 22066 5556 22094 5664
rect 22649 5661 22661 5664
rect 22695 5661 22707 5695
rect 22649 5655 22707 5661
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 23845 5627 23903 5633
rect 23845 5593 23857 5627
rect 23891 5624 23903 5627
rect 24946 5624 24952 5636
rect 23891 5596 24952 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 24946 5584 24952 5596
rect 25004 5584 25010 5636
rect 20763 5528 22094 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 25222 5516 25228 5568
rect 25280 5516 25286 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 13538 5312 13544 5364
rect 13596 5312 13602 5364
rect 14001 5355 14059 5361
rect 14001 5352 14013 5355
rect 13740 5324 14013 5352
rect 2406 5244 2412 5296
rect 2464 5284 2470 5296
rect 2464 5256 2774 5284
rect 2464 5244 2470 5256
rect 2746 5012 2774 5256
rect 12802 5176 12808 5228
rect 12860 5216 12866 5228
rect 13740 5225 13768 5324
rect 14001 5321 14013 5324
rect 14047 5321 14059 5355
rect 14001 5315 14059 5321
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14734 5352 14740 5364
rect 14148 5324 14740 5352
rect 14148 5312 14154 5324
rect 14734 5312 14740 5324
rect 14792 5312 14798 5364
rect 15562 5312 15568 5364
rect 15620 5312 15626 5364
rect 16853 5355 16911 5361
rect 16853 5321 16865 5355
rect 16899 5352 16911 5355
rect 17586 5352 17592 5364
rect 16899 5324 17592 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18233 5355 18291 5361
rect 18233 5352 18245 5355
rect 18012 5324 18245 5352
rect 18012 5312 18018 5324
rect 18233 5321 18245 5324
rect 18279 5352 18291 5355
rect 18966 5352 18972 5364
rect 18279 5324 18972 5352
rect 18279 5321 18291 5324
rect 18233 5315 18291 5321
rect 18966 5312 18972 5324
rect 19024 5312 19030 5364
rect 20898 5352 20904 5364
rect 19628 5324 20904 5352
rect 18506 5244 18512 5296
rect 18564 5284 18570 5296
rect 19628 5284 19656 5324
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 25314 5352 25320 5364
rect 23216 5324 25320 5352
rect 22830 5284 22836 5296
rect 18564 5256 19656 5284
rect 19720 5256 22836 5284
rect 18564 5244 18570 5256
rect 13725 5219 13783 5225
rect 13725 5216 13737 5219
rect 12860 5188 13737 5216
rect 12860 5176 12866 5188
rect 13725 5185 13737 5188
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5216 15807 5219
rect 15795 5188 16160 5216
rect 15795 5185 15807 5188
rect 15749 5179 15807 5185
rect 16132 5157 16160 5188
rect 17034 5176 17040 5228
rect 17092 5176 17098 5228
rect 17586 5176 17592 5228
rect 17644 5220 17650 5228
rect 17681 5220 17739 5225
rect 17644 5219 17739 5220
rect 17644 5192 17693 5219
rect 17644 5176 17650 5192
rect 17681 5185 17693 5192
rect 17727 5185 17739 5219
rect 17681 5179 17739 5185
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 19720 5225 19748 5256
rect 22830 5244 22836 5256
rect 22888 5244 22894 5296
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 18012 5188 18613 5216
rect 18012 5176 18018 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 19705 5219 19763 5225
rect 19705 5185 19717 5219
rect 19751 5185 19763 5219
rect 19705 5179 19763 5185
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 20349 5219 20407 5225
rect 20349 5216 20361 5219
rect 19944 5188 20361 5216
rect 19944 5176 19950 5188
rect 20349 5185 20361 5188
rect 20395 5185 20407 5219
rect 20349 5179 20407 5185
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 21082 5216 21088 5228
rect 20855 5188 21088 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 21082 5176 21088 5188
rect 21140 5176 21146 5228
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 23216 5216 23244 5324
rect 25314 5312 25320 5324
rect 25372 5312 25378 5364
rect 23293 5287 23351 5293
rect 23293 5253 23305 5287
rect 23339 5284 23351 5287
rect 24854 5284 24860 5296
rect 23339 5256 24860 5284
rect 23339 5253 23351 5256
rect 23293 5247 23351 5253
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 22327 5188 23244 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 23934 5176 23940 5228
rect 23992 5176 23998 5228
rect 14921 5151 14979 5157
rect 14921 5117 14933 5151
rect 14967 5117 14979 5151
rect 14921 5111 14979 5117
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5148 16175 5151
rect 16163 5120 18000 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 8478 5040 8484 5092
rect 8536 5080 8542 5092
rect 12250 5080 12256 5092
rect 8536 5052 12256 5080
rect 8536 5040 8542 5052
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 14936 5080 14964 5111
rect 16390 5080 16396 5092
rect 14936 5052 16396 5080
rect 16390 5040 16396 5052
rect 16448 5040 16454 5092
rect 16482 5040 16488 5092
rect 16540 5040 16546 5092
rect 17494 5040 17500 5092
rect 17552 5040 17558 5092
rect 17586 5040 17592 5092
rect 17644 5080 17650 5092
rect 17862 5080 17868 5092
rect 17644 5052 17868 5080
rect 17644 5040 17650 5052
rect 17862 5040 17868 5052
rect 17920 5040 17926 5092
rect 17972 5080 18000 5120
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 23382 5148 23388 5160
rect 18104 5120 23388 5148
rect 18104 5108 18110 5120
rect 23382 5108 23388 5120
rect 23440 5108 23446 5160
rect 24670 5108 24676 5160
rect 24728 5108 24734 5160
rect 26050 5080 26056 5092
rect 17972 5052 26056 5080
rect 26050 5040 26056 5052
rect 26108 5040 26114 5092
rect 13998 5012 14004 5024
rect 2746 4984 14004 5012
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 17957 5015 18015 5021
rect 17957 5012 17969 5015
rect 17184 4984 17969 5012
rect 17184 4972 17190 4984
rect 17957 4981 17969 4984
rect 18003 4981 18015 5015
rect 17957 4975 18015 4981
rect 19242 4972 19248 5024
rect 19300 4972 19306 5024
rect 20438 4972 20444 5024
rect 20496 5012 20502 5024
rect 21453 5015 21511 5021
rect 21453 5012 21465 5015
rect 20496 4984 21465 5012
rect 20496 4972 20502 4984
rect 21453 4981 21465 4984
rect 21499 4981 21511 5015
rect 21453 4975 21511 4981
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 8662 4808 8668 4820
rect 8619 4780 8668 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 16025 4811 16083 4817
rect 16025 4808 16037 4811
rect 10836 4780 16037 4808
rect 10836 4768 10842 4780
rect 16025 4777 16037 4780
rect 16071 4777 16083 4811
rect 16025 4771 16083 4777
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 16850 4808 16856 4820
rect 16715 4780 16856 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 17126 4768 17132 4820
rect 17184 4768 17190 4820
rect 19610 4768 19616 4820
rect 19668 4808 19674 4820
rect 20349 4811 20407 4817
rect 20349 4808 20361 4811
rect 19668 4780 20361 4808
rect 19668 4768 19674 4780
rect 20349 4777 20361 4780
rect 20395 4777 20407 4811
rect 20349 4771 20407 4777
rect 25225 4811 25283 4817
rect 25225 4777 25237 4811
rect 25271 4808 25283 4811
rect 25406 4808 25412 4820
rect 25271 4780 25412 4808
rect 25271 4777 25283 4780
rect 25225 4771 25283 4777
rect 25406 4768 25412 4780
rect 25464 4768 25470 4820
rect 16206 4700 16212 4752
rect 16264 4740 16270 4752
rect 19242 4740 19248 4752
rect 16264 4712 19248 4740
rect 16264 4700 16270 4712
rect 19242 4700 19248 4712
rect 19300 4700 19306 4752
rect 19337 4743 19395 4749
rect 19337 4709 19349 4743
rect 19383 4740 19395 4743
rect 26142 4740 26148 4752
rect 19383 4712 26148 4740
rect 19383 4709 19395 4712
rect 19337 4703 19395 4709
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 17402 4672 17408 4684
rect 14783 4644 17408 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7892 4576 7941 4604
rect 7892 4564 7898 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 15010 4564 15016 4616
rect 15068 4564 15074 4616
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4604 16267 4607
rect 16298 4604 16304 4616
rect 16255 4576 16304 4604
rect 16255 4573 16267 4576
rect 16209 4567 16267 4573
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 16482 4564 16488 4616
rect 16540 4604 16546 4616
rect 16853 4607 16911 4613
rect 16853 4604 16865 4607
rect 16540 4576 16865 4604
rect 16540 4564 16546 4576
rect 16853 4573 16865 4576
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 17126 4564 17132 4616
rect 17184 4604 17190 4616
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 17184 4576 17325 4604
rect 17184 4564 17190 4576
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4604 18199 4607
rect 19352 4604 19380 4703
rect 26142 4700 26148 4712
rect 26200 4700 26206 4752
rect 23750 4672 23756 4684
rect 21008 4644 23756 4672
rect 18187 4576 19380 4604
rect 19705 4607 19763 4613
rect 18187 4573 18199 4576
rect 18141 4567 18199 4573
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 20438 4604 20444 4616
rect 19751 4576 20444 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 20438 4564 20444 4576
rect 20496 4564 20502 4616
rect 21008 4613 21036 4644
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 22462 4564 22468 4616
rect 22520 4604 22526 4616
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22520 4576 22661 4604
rect 22520 4564 22526 4576
rect 22649 4573 22661 4576
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 25038 4604 25044 4616
rect 24627 4576 25044 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 25038 4564 25044 4576
rect 25096 4564 25102 4616
rect 10042 4496 10048 4548
rect 10100 4536 10106 4548
rect 18046 4536 18052 4548
rect 10100 4508 18052 4536
rect 10100 4496 10106 4508
rect 18046 4496 18052 4508
rect 18104 4496 18110 4548
rect 18690 4496 18696 4548
rect 18748 4496 18754 4548
rect 18877 4539 18935 4545
rect 18877 4505 18889 4539
rect 18923 4536 18935 4539
rect 22005 4539 22063 4545
rect 18923 4508 20484 4536
rect 18923 4505 18935 4508
rect 18877 4499 18935 4505
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 17862 4468 17868 4480
rect 14884 4440 17868 4468
rect 14884 4428 14890 4440
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 17954 4428 17960 4480
rect 18012 4428 18018 4480
rect 20456 4468 20484 4508
rect 22005 4505 22017 4539
rect 22051 4536 22063 4539
rect 23382 4536 23388 4548
rect 22051 4508 23388 4536
rect 22051 4505 22063 4508
rect 22005 4499 22063 4505
rect 23382 4496 23388 4508
rect 23440 4496 23446 4548
rect 23845 4539 23903 4545
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 24946 4536 24952 4548
rect 23891 4508 24952 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 22646 4468 22652 4480
rect 20456 4440 22652 4468
rect 22646 4428 22652 4440
rect 22704 4428 22710 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 16298 4224 16304 4276
rect 16356 4224 16362 4276
rect 16390 4224 16396 4276
rect 16448 4264 16454 4276
rect 26326 4264 26332 4276
rect 16448 4236 26332 4264
rect 16448 4224 16454 4236
rect 26326 4224 26332 4236
rect 26384 4224 26390 4276
rect 10318 4156 10324 4208
rect 10376 4196 10382 4208
rect 18690 4196 18696 4208
rect 10376 4168 18696 4196
rect 10376 4156 10382 4168
rect 18690 4156 18696 4168
rect 18748 4156 18754 4208
rect 19150 4156 19156 4208
rect 19208 4196 19214 4208
rect 26418 4196 26424 4208
rect 19208 4168 26424 4196
rect 19208 4156 19214 4168
rect 26418 4156 26424 4168
rect 26476 4156 26482 4208
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4128 6883 4131
rect 9122 4128 9128 4140
rect 6871 4100 9128 4128
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 16942 4128 16948 4140
rect 10928 4100 16948 4128
rect 10928 4088 10934 4100
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17034 4088 17040 4140
rect 17092 4088 17098 4140
rect 18230 4128 18236 4140
rect 17144 4100 18236 4128
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 13538 4060 13544 4072
rect 12492 4032 13544 4060
rect 12492 4020 12498 4032
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 17144 4060 17172 4100
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4128 18383 4131
rect 18598 4128 18604 4140
rect 18371 4100 18604 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4128 19027 4131
rect 19334 4128 19340 4140
rect 19015 4100 19340 4128
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19613 4131 19671 4137
rect 19613 4097 19625 4131
rect 19659 4128 19671 4131
rect 19978 4128 19984 4140
rect 19659 4100 19984 4128
rect 19659 4097 19671 4100
rect 19613 4091 19671 4097
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 22097 4131 22155 4137
rect 22097 4128 22109 4131
rect 20732 4100 22109 4128
rect 14332 4032 17172 4060
rect 17405 4063 17463 4069
rect 14332 4020 14338 4032
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 17494 4060 17500 4072
rect 17451 4032 17500 4060
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 17494 4020 17500 4032
rect 17552 4020 17558 4072
rect 17770 4020 17776 4072
rect 17828 4060 17834 4072
rect 20732 4060 20760 4100
rect 22097 4097 22109 4100
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23937 4131 23995 4137
rect 23937 4128 23949 4131
rect 23532 4100 23949 4128
rect 23532 4088 23538 4100
rect 23937 4097 23949 4100
rect 23983 4097 23995 4131
rect 23937 4091 23995 4097
rect 17828 4032 20760 4060
rect 21269 4063 21327 4069
rect 17828 4020 17834 4032
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 22278 4060 22284 4072
rect 21315 4032 22284 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 22278 4020 22284 4032
rect 22336 4020 22342 4072
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4029 23351 4063
rect 23293 4023 23351 4029
rect 11698 3952 11704 4004
rect 11756 3992 11762 4004
rect 16853 3995 16911 4001
rect 16853 3992 16865 3995
rect 11756 3964 16865 3992
rect 11756 3952 11762 3964
rect 16853 3961 16865 3964
rect 16899 3961 16911 3995
rect 16853 3955 16911 3961
rect 16942 3952 16948 4004
rect 17000 3992 17006 4004
rect 19150 3992 19156 4004
rect 17000 3964 19156 3992
rect 17000 3952 17006 3964
rect 19150 3952 19156 3964
rect 19208 3952 19214 4004
rect 23308 3992 23336 4023
rect 24762 4020 24768 4072
rect 24820 4020 24826 4072
rect 24946 3992 24952 4004
rect 23308 3964 24952 3992
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 7374 3884 7380 3936
rect 7432 3924 7438 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 7432 3896 7481 3924
rect 7432 3884 7438 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 18141 3927 18199 3933
rect 18141 3924 18153 3927
rect 13596 3896 18153 3924
rect 13596 3884 13602 3896
rect 18141 3893 18153 3896
rect 18187 3893 18199 3927
rect 18141 3887 18199 3893
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 18785 3927 18843 3933
rect 18785 3924 18797 3927
rect 18288 3896 18797 3924
rect 18288 3884 18294 3896
rect 18785 3893 18797 3896
rect 18831 3893 18843 3927
rect 18785 3887 18843 3893
rect 19426 3884 19432 3936
rect 19484 3884 19490 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 8205 3723 8263 3729
rect 8205 3720 8217 3723
rect 7892 3692 8217 3720
rect 7892 3680 7898 3692
rect 8205 3689 8217 3692
rect 8251 3689 8263 3723
rect 8205 3683 8263 3689
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 16393 3723 16451 3729
rect 16393 3720 16405 3723
rect 10744 3692 16405 3720
rect 10744 3680 10750 3692
rect 16393 3689 16405 3692
rect 16439 3689 16451 3723
rect 16393 3683 16451 3689
rect 17405 3723 17463 3729
rect 17405 3689 17417 3723
rect 17451 3720 17463 3723
rect 18322 3720 18328 3732
rect 17451 3692 18328 3720
rect 17451 3689 17463 3692
rect 17405 3683 17463 3689
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 6472 3448 6500 3479
rect 7558 3476 7564 3528
rect 7616 3476 7622 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 16408 3516 16436 3683
rect 18322 3680 18328 3692
rect 18380 3680 18386 3732
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 19702 3720 19708 3732
rect 18739 3692 19708 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 19702 3680 19708 3692
rect 19760 3680 19766 3732
rect 20349 3723 20407 3729
rect 20349 3689 20361 3723
rect 20395 3720 20407 3723
rect 20530 3720 20536 3732
rect 20395 3692 20536 3720
rect 20395 3689 20407 3692
rect 20349 3683 20407 3689
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 25225 3723 25283 3729
rect 25225 3689 25237 3723
rect 25271 3720 25283 3723
rect 25590 3720 25596 3732
rect 25271 3692 25596 3720
rect 25271 3689 25283 3692
rect 25225 3683 25283 3689
rect 25590 3680 25596 3692
rect 25648 3680 25654 3732
rect 17678 3612 17684 3664
rect 17736 3652 17742 3664
rect 20070 3652 20076 3664
rect 17736 3624 20076 3652
rect 17736 3612 17742 3624
rect 20070 3612 20076 3624
rect 20128 3612 20134 3664
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3584 16819 3587
rect 19518 3584 19524 3596
rect 16807 3556 19524 3584
rect 16807 3553 16819 3556
rect 16761 3547 16819 3553
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 25130 3584 25136 3596
rect 19720 3556 25136 3584
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 9456 3488 12434 3516
rect 16408 3488 17601 3516
rect 9456 3476 9462 3488
rect 9766 3448 9772 3460
rect 6472 3420 9772 3448
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 12406 3448 12434 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 18230 3476 18236 3528
rect 18288 3476 18294 3528
rect 18874 3476 18880 3528
rect 18932 3476 18938 3528
rect 19720 3525 19748 3556
rect 25130 3544 25136 3556
rect 25188 3544 25194 3596
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 20993 3519 21051 3525
rect 20993 3485 21005 3519
rect 21039 3516 21051 3519
rect 21910 3516 21916 3528
rect 21039 3488 21916 3516
rect 21039 3485 21051 3488
rect 20993 3479 21051 3485
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 22646 3476 22652 3528
rect 22704 3476 22710 3528
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3516 24639 3519
rect 25222 3516 25228 3528
rect 24627 3488 25228 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 19429 3451 19487 3457
rect 12406 3420 18092 3448
rect 7101 3383 7159 3389
rect 7101 3349 7113 3383
rect 7147 3380 7159 3383
rect 8478 3380 8484 3392
rect 7147 3352 8484 3380
rect 7147 3349 7159 3352
rect 7101 3343 7159 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 18064 3389 18092 3420
rect 19429 3417 19441 3451
rect 19475 3448 19487 3451
rect 19978 3448 19984 3460
rect 19475 3420 19984 3448
rect 19475 3417 19487 3420
rect 19429 3411 19487 3417
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 22005 3451 22063 3457
rect 22005 3417 22017 3451
rect 22051 3448 22063 3451
rect 23382 3448 23388 3460
rect 22051 3420 23388 3448
rect 22051 3417 22063 3420
rect 22005 3411 22063 3417
rect 23382 3408 23388 3420
rect 23440 3408 23446 3460
rect 23845 3451 23903 3457
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 25682 3448 25688 3460
rect 23891 3420 25688 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 25682 3408 25688 3420
rect 25740 3408 25746 3460
rect 18049 3383 18107 3389
rect 18049 3349 18061 3383
rect 18095 3349 18107 3383
rect 18049 3343 18107 3349
rect 20438 3340 20444 3392
rect 20496 3380 20502 3392
rect 24486 3380 24492 3392
rect 20496 3352 24492 3380
rect 20496 3340 20502 3352
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 9122 3136 9128 3188
rect 9180 3136 9186 3188
rect 16853 3179 16911 3185
rect 16853 3145 16865 3179
rect 16899 3176 16911 3179
rect 16945 3179 17003 3185
rect 16945 3176 16957 3179
rect 16899 3148 16957 3176
rect 16899 3145 16911 3148
rect 16853 3139 16911 3145
rect 16945 3145 16957 3148
rect 16991 3176 17003 3179
rect 17586 3176 17592 3188
rect 16991 3148 17592 3176
rect 16991 3145 17003 3148
rect 16945 3139 17003 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 20438 3176 20444 3188
rect 17788 3148 20444 3176
rect 16485 3111 16543 3117
rect 16485 3077 16497 3111
rect 16531 3108 16543 3111
rect 17788 3108 17816 3148
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 16531 3080 17816 3108
rect 16531 3077 16543 3080
rect 16485 3071 16543 3077
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 8478 3000 8484 3052
rect 8536 3000 8542 3052
rect 17788 3049 17816 3080
rect 19429 3111 19487 3117
rect 19429 3077 19441 3111
rect 19475 3108 19487 3111
rect 22186 3108 22192 3120
rect 19475 3080 22192 3108
rect 19475 3077 19487 3080
rect 19429 3071 19487 3077
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 23293 3111 23351 3117
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24854 3108 24860 3120
rect 23339 3080 24860 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3009 17831 3043
rect 17773 3003 17831 3009
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 20257 3043 20315 3049
rect 20257 3009 20269 3043
rect 20303 3040 20315 3043
rect 21818 3040 21824 3052
rect 20303 3012 21824 3040
rect 20303 3009 20315 3012
rect 20257 3003 20315 3009
rect 18432 2972 18460 3003
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 22094 3000 22100 3052
rect 22152 3000 22158 3052
rect 24121 3043 24179 3049
rect 24121 3009 24133 3043
rect 24167 3040 24179 3043
rect 26602 3040 26608 3052
rect 24167 3012 26608 3040
rect 24167 3009 24179 3012
rect 24121 3003 24179 3009
rect 26602 3000 26608 3012
rect 26660 3000 26666 3052
rect 21174 2972 21180 2984
rect 18432 2944 21180 2972
rect 21174 2932 21180 2944
rect 21232 2932 21238 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 21315 2944 22094 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 8662 2904 8668 2916
rect 6788 2876 8668 2904
rect 6788 2864 6794 2876
rect 8662 2864 8668 2876
rect 8720 2864 8726 2916
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 17589 2907 17647 2913
rect 17589 2904 17601 2907
rect 11020 2876 17601 2904
rect 11020 2864 11026 2876
rect 17589 2873 17601 2876
rect 17635 2873 17647 2907
rect 22066 2904 22094 2944
rect 24578 2932 24584 2984
rect 24636 2932 24642 2984
rect 25038 2904 25044 2916
rect 22066 2876 25044 2904
rect 17589 2867 17647 2873
rect 25038 2864 25044 2876
rect 25096 2864 25102 2916
rect 7190 2796 7196 2848
rect 7248 2836 7254 2848
rect 8021 2839 8079 2845
rect 8021 2836 8033 2839
rect 7248 2808 8033 2836
rect 7248 2796 7254 2808
rect 8021 2805 8033 2808
rect 8067 2805 8079 2839
rect 8021 2799 8079 2805
rect 20714 2796 20720 2848
rect 20772 2836 20778 2848
rect 22554 2836 22560 2848
rect 20772 2808 22560 2836
rect 20772 2796 20778 2808
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 7558 2632 7564 2644
rect 6779 2604 7564 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8662 2592 8668 2644
rect 8720 2592 8726 2644
rect 9766 2592 9772 2644
rect 9824 2592 9830 2644
rect 17402 2592 17408 2644
rect 17460 2632 17466 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17460 2604 17601 2632
rect 17460 2592 17466 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 17589 2595 17647 2601
rect 18877 2635 18935 2641
rect 18877 2601 18889 2635
rect 18923 2632 18935 2635
rect 22005 2635 22063 2641
rect 18923 2604 20760 2632
rect 18923 2601 18935 2604
rect 18877 2595 18935 2601
rect 7190 2564 7196 2576
rect 5368 2536 7196 2564
rect 5368 2437 5396 2536
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 16945 2567 17003 2573
rect 16945 2533 16957 2567
rect 16991 2564 17003 2567
rect 20732 2564 20760 2604
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 22094 2632 22100 2644
rect 22051 2604 22100 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 22094 2592 22100 2604
rect 22152 2592 22158 2644
rect 25130 2592 25136 2644
rect 25188 2632 25194 2644
rect 25225 2635 25283 2641
rect 25225 2632 25237 2635
rect 25188 2604 25237 2632
rect 25188 2592 25194 2604
rect 25225 2601 25237 2604
rect 25271 2601 25283 2635
rect 25225 2595 25283 2601
rect 23474 2564 23480 2576
rect 16991 2536 20208 2564
rect 20732 2536 23480 2564
rect 16991 2533 17003 2536
rect 16945 2527 17003 2533
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 6932 2468 8033 2496
rect 6932 2437 6960 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8021 2459 8079 2465
rect 13630 2456 13636 2508
rect 13688 2496 13694 2508
rect 18233 2499 18291 2505
rect 18233 2496 18245 2499
rect 13688 2468 18245 2496
rect 13688 2456 13694 2468
rect 18233 2465 18245 2468
rect 18279 2465 18291 2499
rect 18233 2459 18291 2465
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19392 2468 19656 2496
rect 19392 2456 19398 2468
rect 19628 2440 19656 2468
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 5997 2363 6055 2369
rect 5997 2329 6009 2363
rect 6043 2360 6055 2363
rect 7392 2360 7420 2391
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8720 2400 9137 2428
rect 8720 2388 8726 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2397 17187 2431
rect 17129 2391 17187 2397
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2428 17831 2431
rect 19518 2428 19524 2440
rect 17819 2400 19524 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 6043 2332 7420 2360
rect 17144 2360 17172 2391
rect 19518 2388 19524 2400
rect 19576 2388 19582 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2397 20131 2431
rect 20180 2428 20208 2536
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2496 21327 2499
rect 24854 2496 24860 2508
rect 21315 2468 24860 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 20180 2400 22201 2428
rect 20073 2391 20131 2397
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 20088 2360 20116 2391
rect 22646 2388 22652 2440
rect 22704 2388 22710 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 20714 2360 20720 2372
rect 17144 2332 20024 2360
rect 20088 2332 20720 2360
rect 6043 2329 6055 2332
rect 5997 2323 6055 2329
rect 16485 2295 16543 2301
rect 16485 2261 16497 2295
rect 16531 2292 16543 2295
rect 19334 2292 19340 2304
rect 16531 2264 19340 2292
rect 16531 2261 16543 2264
rect 16485 2255 16543 2261
rect 19334 2252 19340 2264
rect 19392 2252 19398 2304
rect 19426 2252 19432 2304
rect 19484 2252 19490 2304
rect 19996 2292 20024 2332
rect 20714 2320 20720 2332
rect 20772 2320 20778 2372
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24946 2360 24952 2372
rect 23891 2332 24952 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 20254 2292 20260 2304
rect 19996 2264 20260 2292
rect 20254 2252 20260 2264
rect 20312 2252 20318 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 15010 2048 15016 2100
rect 15068 2088 15074 2100
rect 22646 2088 22652 2100
rect 15068 2060 22652 2088
rect 15068 2048 15074 2060
rect 22646 2048 22652 2060
rect 22704 2048 22710 2100
rect 12526 1980 12532 2032
rect 12584 2020 12590 2032
rect 19426 2020 19432 2032
rect 12584 1992 19432 2020
rect 12584 1980 12590 1992
rect 19426 1980 19432 1992
rect 19484 1980 19490 2032
rect 19518 1980 19524 2032
rect 19576 2020 19582 2032
rect 24118 2020 24124 2032
rect 19576 1992 24124 2020
rect 19576 1980 19582 1992
rect 24118 1980 24124 1992
rect 24176 1980 24182 2032
rect 17310 1912 17316 1964
rect 17368 1952 17374 1964
rect 24578 1952 24584 1964
rect 17368 1924 24584 1952
rect 17368 1912 17374 1924
rect 24578 1912 24584 1924
rect 24636 1912 24642 1964
rect 13722 1844 13728 1896
rect 13780 1884 13786 1896
rect 19886 1884 19892 1896
rect 13780 1856 19892 1884
rect 13780 1844 13786 1856
rect 19886 1844 19892 1856
rect 19944 1844 19950 1896
rect 11606 1776 11612 1828
rect 11664 1816 11670 1828
rect 20530 1816 20536 1828
rect 11664 1788 20536 1816
rect 11664 1776 11670 1788
rect 20530 1776 20536 1788
rect 20588 1776 20594 1828
<< via1 >>
rect 1032 26324 1084 26376
rect 22560 26324 22612 26376
rect 2136 26256 2188 26308
rect 22192 26256 22244 26308
rect 5448 26188 5500 26240
rect 21272 26188 21324 26240
rect 1584 26120 1636 26172
rect 16672 26120 16724 26172
rect 17316 26120 17368 26172
rect 10968 25916 11020 25968
rect 14188 25916 14240 25968
rect 1860 25848 1912 25900
rect 13728 25848 13780 25900
rect 3424 25780 3476 25832
rect 21732 25780 21784 25832
rect 572 25712 624 25764
rect 20904 25712 20956 25764
rect 2412 25644 2464 25696
rect 15844 25644 15896 25696
rect 2596 25576 2648 25628
rect 20536 25576 20588 25628
rect 7288 25508 7340 25560
rect 22008 25508 22060 25560
rect 4528 25440 4580 25492
rect 24216 25440 24268 25492
rect 5264 25372 5316 25424
rect 24768 25372 24820 25424
rect 4804 25304 4856 25356
rect 19524 25304 19576 25356
rect 4160 25236 4212 25288
rect 17960 25236 18012 25288
rect 3240 25168 3292 25220
rect 9496 25168 9548 25220
rect 12624 25168 12676 25220
rect 24032 25168 24084 25220
rect 6736 25100 6788 25152
rect 13912 25100 13964 25152
rect 1124 24964 1176 25016
rect 14280 25032 14332 25084
rect 756 24896 808 24948
rect 13084 24964 13136 25016
rect 17684 24964 17736 25016
rect 11612 24896 11664 24948
rect 14740 24896 14792 24948
rect 16028 24896 16080 24948
rect 19616 24896 19668 24948
rect 23572 24896 23624 24948
rect 8576 24828 8628 24880
rect 19984 24828 20036 24880
rect 13636 24760 13688 24812
rect 3700 24624 3752 24676
rect 14464 24692 14516 24744
rect 12532 24624 12584 24676
rect 13820 24624 13872 24676
rect 15844 24760 15896 24812
rect 19340 24760 19392 24812
rect 17592 24692 17644 24744
rect 17500 24624 17552 24676
rect 19064 24624 19116 24676
rect 21180 24624 21232 24676
rect 23940 24624 23992 24676
rect 2780 24556 2832 24608
rect 16580 24556 16632 24608
rect 16672 24556 16724 24608
rect 22192 24556 22244 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 6552 24395 6604 24404
rect 6552 24361 6561 24395
rect 6561 24361 6595 24395
rect 6595 24361 6604 24395
rect 6552 24352 6604 24361
rect 8484 24352 8536 24404
rect 15292 24352 15344 24404
rect 3976 24327 4028 24336
rect 3976 24293 3985 24327
rect 3985 24293 4019 24327
rect 4019 24293 4028 24327
rect 3976 24284 4028 24293
rect 6276 24284 6328 24336
rect 6460 24216 6512 24268
rect 6644 24284 6696 24336
rect 16488 24284 16540 24336
rect 2320 24148 2372 24200
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 4436 24148 4488 24200
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 5908 24148 5960 24200
rect 7196 24191 7248 24200
rect 7196 24157 7205 24191
rect 7205 24157 7239 24191
rect 7239 24157 7248 24191
rect 7196 24148 7248 24157
rect 9680 24216 9732 24268
rect 11244 24216 11296 24268
rect 12440 24216 12492 24268
rect 14740 24259 14792 24268
rect 14740 24225 14749 24259
rect 14749 24225 14783 24259
rect 14783 24225 14792 24259
rect 14740 24216 14792 24225
rect 17408 24259 17460 24268
rect 17408 24225 17417 24259
rect 17417 24225 17451 24259
rect 17451 24225 17460 24259
rect 17408 24216 17460 24225
rect 17592 24259 17644 24268
rect 17592 24225 17601 24259
rect 17601 24225 17635 24259
rect 17635 24225 17644 24259
rect 17592 24216 17644 24225
rect 8668 24080 8720 24132
rect 12348 24191 12400 24200
rect 12348 24157 12357 24191
rect 12357 24157 12391 24191
rect 12391 24157 12400 24191
rect 12348 24148 12400 24157
rect 13452 24148 13504 24200
rect 16580 24148 16632 24200
rect 7012 24012 7064 24064
rect 7748 24012 7800 24064
rect 11244 24012 11296 24064
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 16212 24080 16264 24132
rect 16764 24080 16816 24132
rect 18144 24395 18196 24404
rect 18144 24361 18153 24395
rect 18153 24361 18187 24395
rect 18187 24361 18196 24395
rect 18144 24352 18196 24361
rect 18328 24352 18380 24404
rect 19432 24352 19484 24404
rect 19616 24395 19668 24404
rect 19616 24361 19625 24395
rect 19625 24361 19659 24395
rect 19659 24361 19668 24395
rect 19616 24352 19668 24361
rect 19984 24395 20036 24404
rect 19984 24361 19993 24395
rect 19993 24361 20027 24395
rect 20027 24361 20036 24395
rect 19984 24352 20036 24361
rect 21732 24352 21784 24404
rect 23940 24395 23992 24404
rect 23940 24361 23949 24395
rect 23949 24361 23983 24395
rect 23983 24361 23992 24395
rect 23940 24352 23992 24361
rect 25504 24352 25556 24404
rect 18972 24284 19024 24336
rect 20260 24284 20312 24336
rect 19708 24216 19760 24268
rect 19800 24216 19852 24268
rect 21180 24327 21232 24336
rect 21180 24293 21189 24327
rect 21189 24293 21223 24327
rect 21223 24293 21232 24327
rect 21180 24284 21232 24293
rect 25044 24284 25096 24336
rect 22560 24216 22612 24268
rect 25320 24216 25372 24268
rect 23756 24148 23808 24200
rect 25136 24148 25188 24200
rect 15936 24012 15988 24064
rect 16120 24055 16172 24064
rect 16120 24021 16129 24055
rect 16129 24021 16163 24055
rect 16163 24021 16172 24055
rect 16120 24012 16172 24021
rect 17224 24012 17276 24064
rect 18604 24055 18656 24064
rect 18604 24021 18613 24055
rect 18613 24021 18647 24055
rect 18647 24021 18656 24055
rect 18604 24012 18656 24021
rect 19340 24055 19392 24064
rect 19340 24021 19349 24055
rect 19349 24021 19383 24055
rect 19383 24021 19392 24055
rect 19984 24080 20036 24132
rect 21272 24080 21324 24132
rect 19340 24012 19392 24021
rect 20536 24055 20588 24064
rect 20536 24021 20545 24055
rect 20545 24021 20579 24055
rect 20579 24021 20588 24055
rect 20536 24012 20588 24021
rect 22376 24012 22428 24064
rect 23848 24012 23900 24064
rect 25596 24012 25648 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 7380 23808 7432 23860
rect 12164 23740 12216 23792
rect 2596 23672 2648 23724
rect 2964 23715 3016 23724
rect 2964 23681 2973 23715
rect 2973 23681 3007 23715
rect 3007 23681 3016 23715
rect 2964 23672 3016 23681
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 5356 23604 5408 23656
rect 1768 23468 1820 23520
rect 6644 23672 6696 23724
rect 6828 23715 6880 23724
rect 6828 23681 6837 23715
rect 6837 23681 6871 23715
rect 6871 23681 6880 23715
rect 6828 23672 6880 23681
rect 7840 23672 7892 23724
rect 9588 23672 9640 23724
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 10876 23715 10928 23724
rect 10876 23681 10885 23715
rect 10885 23681 10919 23715
rect 10919 23681 10928 23715
rect 10876 23672 10928 23681
rect 7564 23604 7616 23656
rect 9220 23604 9272 23656
rect 12440 23808 12492 23860
rect 13636 23808 13688 23860
rect 13912 23808 13964 23860
rect 15568 23808 15620 23860
rect 13360 23740 13412 23792
rect 18512 23808 18564 23860
rect 18604 23808 18656 23860
rect 18328 23740 18380 23792
rect 20168 23740 20220 23792
rect 22376 23808 22428 23860
rect 20720 23783 20772 23792
rect 20720 23749 20729 23783
rect 20729 23749 20763 23783
rect 20763 23749 20772 23783
rect 20720 23740 20772 23749
rect 22468 23740 22520 23792
rect 23388 23740 23440 23792
rect 11980 23604 12032 23656
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15335 23715
rect 15335 23681 15344 23715
rect 15292 23672 15344 23681
rect 17316 23715 17368 23724
rect 17316 23681 17325 23715
rect 17325 23681 17359 23715
rect 17359 23681 17368 23715
rect 17316 23672 17368 23681
rect 21364 23672 21416 23724
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 25412 23672 25464 23724
rect 7196 23536 7248 23588
rect 9680 23536 9732 23588
rect 5816 23468 5868 23520
rect 6644 23468 6696 23520
rect 11612 23511 11664 23520
rect 11612 23477 11621 23511
rect 11621 23477 11655 23511
rect 11655 23477 11664 23511
rect 11612 23468 11664 23477
rect 11704 23511 11756 23520
rect 11704 23477 11713 23511
rect 11713 23477 11747 23511
rect 11747 23477 11756 23511
rect 11704 23468 11756 23477
rect 13728 23468 13780 23520
rect 14096 23579 14148 23588
rect 14096 23545 14105 23579
rect 14105 23545 14139 23579
rect 14139 23545 14148 23579
rect 14096 23536 14148 23545
rect 14648 23647 14700 23656
rect 14648 23613 14657 23647
rect 14657 23613 14691 23647
rect 14691 23613 14700 23647
rect 14648 23604 14700 23613
rect 16948 23604 17000 23656
rect 14832 23468 14884 23520
rect 16488 23511 16540 23520
rect 16488 23477 16497 23511
rect 16497 23477 16531 23511
rect 16531 23477 16540 23511
rect 16488 23468 16540 23477
rect 17040 23536 17092 23588
rect 17776 23468 17828 23520
rect 18788 23604 18840 23656
rect 19708 23604 19760 23656
rect 20720 23604 20772 23656
rect 20904 23647 20956 23656
rect 20904 23613 20913 23647
rect 20913 23613 20947 23647
rect 20947 23613 20956 23647
rect 20904 23604 20956 23613
rect 20996 23604 21048 23656
rect 22468 23604 22520 23656
rect 22652 23647 22704 23656
rect 22652 23613 22661 23647
rect 22661 23613 22695 23647
rect 22695 23613 22704 23647
rect 22652 23604 22704 23613
rect 21088 23536 21140 23588
rect 25228 23579 25280 23588
rect 25228 23545 25237 23579
rect 25237 23545 25271 23579
rect 25271 23545 25280 23579
rect 25228 23536 25280 23545
rect 18328 23468 18380 23520
rect 19800 23511 19852 23520
rect 19800 23477 19809 23511
rect 19809 23477 19843 23511
rect 19843 23477 19852 23511
rect 19800 23468 19852 23477
rect 20076 23468 20128 23520
rect 21548 23511 21600 23520
rect 21548 23477 21557 23511
rect 21557 23477 21591 23511
rect 21591 23477 21600 23511
rect 21548 23468 21600 23477
rect 24400 23511 24452 23520
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 3700 23264 3752 23316
rect 9680 23264 9732 23316
rect 11888 23264 11940 23316
rect 12532 23264 12584 23316
rect 12624 23264 12676 23316
rect 13452 23264 13504 23316
rect 13544 23264 13596 23316
rect 15844 23264 15896 23316
rect 16580 23264 16632 23316
rect 17868 23264 17920 23316
rect 3148 23196 3200 23248
rect 4620 23128 4672 23180
rect 7656 23128 7708 23180
rect 9312 23128 9364 23180
rect 9404 23128 9456 23180
rect 12992 23196 13044 23248
rect 14648 23128 14700 23180
rect 16304 23196 16356 23248
rect 17408 23128 17460 23180
rect 17500 23128 17552 23180
rect 18696 23239 18748 23248
rect 18696 23205 18705 23239
rect 18705 23205 18739 23239
rect 18739 23205 18748 23239
rect 18696 23196 18748 23205
rect 18880 23196 18932 23248
rect 20260 23264 20312 23316
rect 20720 23264 20772 23316
rect 24308 23264 24360 23316
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 4252 23103 4304 23112
rect 4252 23069 4261 23103
rect 4261 23069 4295 23103
rect 4295 23069 4304 23103
rect 4252 23060 4304 23069
rect 6552 23060 6604 23112
rect 3700 22924 3752 22976
rect 4620 22924 4672 22976
rect 6184 22924 6236 22976
rect 7288 23060 7340 23112
rect 9220 23103 9272 23112
rect 9220 23069 9229 23103
rect 9229 23069 9263 23103
rect 9263 23069 9272 23103
rect 9220 23060 9272 23069
rect 9496 23103 9548 23112
rect 9496 23069 9505 23103
rect 9505 23069 9539 23103
rect 9539 23069 9548 23103
rect 9496 23060 9548 23069
rect 13360 23060 13412 23112
rect 13636 23060 13688 23112
rect 16672 23060 16724 23112
rect 17040 23060 17092 23112
rect 18972 23060 19024 23112
rect 10600 22992 10652 23044
rect 10784 22924 10836 22976
rect 11612 22924 11664 22976
rect 12256 22992 12308 23044
rect 13176 22992 13228 23044
rect 12348 22967 12400 22976
rect 12348 22933 12357 22967
rect 12357 22933 12391 22967
rect 12391 22933 12400 22967
rect 12348 22924 12400 22933
rect 12624 22924 12676 22976
rect 12808 22924 12860 22976
rect 14372 23035 14424 23044
rect 14372 23001 14381 23035
rect 14381 23001 14415 23035
rect 14415 23001 14424 23035
rect 14372 22992 14424 23001
rect 14556 23035 14608 23044
rect 14556 23001 14565 23035
rect 14565 23001 14599 23035
rect 14599 23001 14608 23035
rect 14556 22992 14608 23001
rect 14740 22992 14792 23044
rect 16948 22992 17000 23044
rect 18880 22992 18932 23044
rect 17132 22924 17184 22976
rect 17224 22967 17276 22976
rect 17224 22933 17233 22967
rect 17233 22933 17267 22967
rect 17267 22933 17276 22967
rect 17224 22924 17276 22933
rect 17684 22967 17736 22976
rect 17684 22933 17693 22967
rect 17693 22933 17727 22967
rect 17727 22933 17736 22967
rect 17684 22924 17736 22933
rect 22652 23128 22704 23180
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 23388 23060 23440 23112
rect 24952 23103 25004 23112
rect 24952 23069 24961 23103
rect 24961 23069 24995 23103
rect 24995 23069 25004 23103
rect 24952 23060 25004 23069
rect 25228 23060 25280 23112
rect 19708 23035 19760 23044
rect 19708 23001 19717 23035
rect 19717 23001 19751 23035
rect 19751 23001 19760 23035
rect 19708 22992 19760 23001
rect 20168 22992 20220 23044
rect 21916 23035 21968 23044
rect 21916 23001 21925 23035
rect 21925 23001 21959 23035
rect 21959 23001 21968 23035
rect 21916 22992 21968 23001
rect 20536 22924 20588 22976
rect 22284 22924 22336 22976
rect 26884 22992 26936 23044
rect 23388 22967 23440 22976
rect 23388 22933 23397 22967
rect 23397 22933 23431 22967
rect 23431 22933 23440 22967
rect 23388 22924 23440 22933
rect 23848 22967 23900 22976
rect 23848 22933 23857 22967
rect 23857 22933 23891 22967
rect 23891 22933 23900 22967
rect 23848 22924 23900 22933
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 2504 22720 2556 22772
rect 3424 22720 3476 22772
rect 6000 22720 6052 22772
rect 6736 22720 6788 22772
rect 7012 22763 7064 22772
rect 7012 22729 7021 22763
rect 7021 22729 7055 22763
rect 7055 22729 7064 22763
rect 7012 22720 7064 22729
rect 11796 22720 11848 22772
rect 14740 22720 14792 22772
rect 3148 22652 3200 22704
rect 4160 22652 4212 22704
rect 5724 22695 5776 22704
rect 5724 22661 5733 22695
rect 5733 22661 5767 22695
rect 5767 22661 5776 22695
rect 5724 22652 5776 22661
rect 8760 22695 8812 22704
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 11612 22652 11664 22704
rect 12532 22652 12584 22704
rect 13544 22652 13596 22704
rect 15292 22720 15344 22772
rect 16948 22720 17000 22772
rect 17132 22720 17184 22772
rect 15476 22652 15528 22704
rect 17868 22652 17920 22704
rect 18420 22720 18472 22772
rect 20536 22720 20588 22772
rect 22560 22720 22612 22772
rect 23112 22720 23164 22772
rect 24952 22720 25004 22772
rect 3608 22584 3660 22636
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 7104 22584 7156 22636
rect 6368 22516 6420 22568
rect 8944 22584 8996 22636
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 11152 22584 11204 22636
rect 12164 22584 12216 22636
rect 9772 22516 9824 22568
rect 11704 22559 11756 22568
rect 11704 22525 11713 22559
rect 11713 22525 11747 22559
rect 11747 22525 11756 22559
rect 11704 22516 11756 22525
rect 12072 22516 12124 22568
rect 12440 22516 12492 22568
rect 12716 22584 12768 22636
rect 13452 22584 13504 22636
rect 13636 22627 13688 22636
rect 13636 22593 13645 22627
rect 13645 22593 13679 22627
rect 13679 22593 13688 22627
rect 13636 22584 13688 22593
rect 15936 22627 15988 22636
rect 15936 22593 15945 22627
rect 15945 22593 15979 22627
rect 15979 22593 15988 22627
rect 15936 22584 15988 22593
rect 16028 22584 16080 22636
rect 14004 22516 14056 22568
rect 5540 22448 5592 22500
rect 9404 22448 9456 22500
rect 1676 22380 1728 22432
rect 3424 22380 3476 22432
rect 11336 22380 11388 22432
rect 12992 22423 13044 22432
rect 12992 22389 13001 22423
rect 13001 22389 13035 22423
rect 13035 22389 13044 22423
rect 12992 22380 13044 22389
rect 15752 22448 15804 22500
rect 16948 22516 17000 22568
rect 18604 22584 18656 22636
rect 19616 22627 19668 22636
rect 19616 22593 19625 22627
rect 19625 22593 19659 22627
rect 19659 22593 19668 22627
rect 19616 22584 19668 22593
rect 17592 22516 17644 22568
rect 13912 22380 13964 22432
rect 14648 22380 14700 22432
rect 15844 22380 15896 22432
rect 17776 22448 17828 22500
rect 18236 22448 18288 22500
rect 18420 22448 18472 22500
rect 18972 22516 19024 22568
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 19156 22448 19208 22500
rect 21456 22627 21508 22636
rect 21456 22593 21465 22627
rect 21465 22593 21499 22627
rect 21499 22593 21508 22627
rect 21456 22584 21508 22593
rect 20720 22448 20772 22500
rect 21548 22516 21600 22568
rect 22652 22652 22704 22704
rect 22284 22584 22336 22636
rect 23296 22652 23348 22704
rect 23940 22652 23992 22704
rect 21732 22516 21784 22568
rect 22560 22516 22612 22568
rect 24860 22516 24912 22568
rect 23112 22380 23164 22432
rect 26056 22380 26108 22432
rect 26700 22380 26752 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 1860 22176 1912 22228
rect 5632 22176 5684 22228
rect 13360 22176 13412 22228
rect 13452 22219 13504 22228
rect 13452 22185 13461 22219
rect 13461 22185 13495 22219
rect 13495 22185 13504 22219
rect 13452 22176 13504 22185
rect 14188 22176 14240 22228
rect 15200 22176 15252 22228
rect 15752 22176 15804 22228
rect 16212 22176 16264 22228
rect 9404 22108 9456 22160
rect 12348 22108 12400 22160
rect 17408 22108 17460 22160
rect 17776 22108 17828 22160
rect 19984 22176 20036 22228
rect 20996 22176 21048 22228
rect 24492 22176 24544 22228
rect 2504 22040 2556 22092
rect 3332 22040 3384 22092
rect 3792 22040 3844 22092
rect 7840 22040 7892 22092
rect 8208 22054 8260 22106
rect 8852 22040 8904 22092
rect 9220 22040 9272 22092
rect 1860 21972 1912 22024
rect 3976 21904 4028 21956
rect 5448 22015 5500 22024
rect 5448 21981 5457 22015
rect 5457 21981 5491 22015
rect 5491 21981 5500 22015
rect 5448 21972 5500 21981
rect 7288 21972 7340 22024
rect 7380 22015 7432 22024
rect 7380 21981 7389 22015
rect 7389 21981 7423 22015
rect 7423 21981 7432 22015
rect 7380 21972 7432 21981
rect 12624 22040 12676 22092
rect 12992 22083 13044 22092
rect 12992 22049 13001 22083
rect 13001 22049 13035 22083
rect 13035 22049 13044 22083
rect 12992 22040 13044 22049
rect 14832 22083 14884 22092
rect 14832 22049 14841 22083
rect 14841 22049 14875 22083
rect 14875 22049 14884 22083
rect 14832 22040 14884 22049
rect 17040 22040 17092 22092
rect 18052 22040 18104 22092
rect 19064 22108 19116 22160
rect 20352 22108 20404 22160
rect 10048 21972 10100 22024
rect 12440 21972 12492 22024
rect 6092 21904 6144 21956
rect 6736 21904 6788 21956
rect 11060 21904 11112 21956
rect 12624 21904 12676 21956
rect 14464 21972 14516 22024
rect 15660 21972 15712 22024
rect 17132 21972 17184 22024
rect 17868 21972 17920 22024
rect 14372 21904 14424 21956
rect 18236 21972 18288 22024
rect 18420 21972 18472 22024
rect 19432 22040 19484 22092
rect 19524 22040 19576 22092
rect 19064 21972 19116 22024
rect 4620 21836 4672 21888
rect 4988 21836 5040 21888
rect 5356 21836 5408 21888
rect 8852 21836 8904 21888
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 9220 21836 9272 21888
rect 9680 21836 9732 21888
rect 9864 21836 9916 21888
rect 11152 21836 11204 21888
rect 12440 21879 12492 21888
rect 12440 21845 12449 21879
rect 12449 21845 12483 21879
rect 12483 21845 12492 21879
rect 12440 21836 12492 21845
rect 14004 21836 14056 21888
rect 14280 21879 14332 21888
rect 14280 21845 14289 21879
rect 14289 21845 14323 21879
rect 14323 21845 14332 21879
rect 14280 21836 14332 21845
rect 15292 21879 15344 21888
rect 15292 21845 15301 21879
rect 15301 21845 15335 21879
rect 15335 21845 15344 21879
rect 15292 21836 15344 21845
rect 17500 21879 17552 21888
rect 17500 21845 17509 21879
rect 17509 21845 17543 21879
rect 17543 21845 17552 21879
rect 17500 21836 17552 21845
rect 18144 21836 18196 21888
rect 18880 21904 18932 21956
rect 19432 21836 19484 21888
rect 20076 21836 20128 21888
rect 20720 21836 20772 21888
rect 22192 21972 22244 22024
rect 23480 22040 23532 22092
rect 25504 22108 25556 22160
rect 23020 21972 23072 22024
rect 25688 21972 25740 22024
rect 22008 21904 22060 21956
rect 23112 21947 23164 21956
rect 23112 21913 23121 21947
rect 23121 21913 23155 21947
rect 23155 21913 23164 21947
rect 23112 21904 23164 21913
rect 22284 21836 22336 21888
rect 24584 21879 24636 21888
rect 24584 21845 24593 21879
rect 24593 21845 24627 21879
rect 24627 21845 24636 21879
rect 24584 21836 24636 21845
rect 24860 21836 24912 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 4252 21632 4304 21684
rect 4804 21632 4856 21684
rect 5356 21632 5408 21684
rect 5724 21632 5776 21684
rect 5908 21632 5960 21684
rect 6092 21632 6144 21684
rect 9220 21632 9272 21684
rect 848 21564 900 21616
rect 13912 21632 13964 21684
rect 16488 21632 16540 21684
rect 17684 21632 17736 21684
rect 11336 21564 11388 21616
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 2136 21496 2188 21548
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 5172 21496 5224 21548
rect 8944 21539 8996 21548
rect 8944 21505 8953 21539
rect 8953 21505 8987 21539
rect 8987 21505 8996 21539
rect 8944 21496 8996 21505
rect 11060 21539 11112 21548
rect 11060 21505 11069 21539
rect 11069 21505 11103 21539
rect 11103 21505 11112 21539
rect 11060 21496 11112 21505
rect 11980 21496 12032 21548
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 5908 21428 5960 21480
rect 6276 21428 6328 21480
rect 6920 21428 6972 21480
rect 7288 21428 7340 21480
rect 7472 21428 7524 21480
rect 10968 21428 11020 21480
rect 11612 21428 11664 21480
rect 12072 21428 12124 21480
rect 12256 21564 12308 21616
rect 12992 21564 13044 21616
rect 13636 21564 13688 21616
rect 13728 21607 13780 21616
rect 13728 21573 13737 21607
rect 13737 21573 13771 21607
rect 13771 21573 13780 21607
rect 13728 21564 13780 21573
rect 14004 21564 14056 21616
rect 15108 21564 15160 21616
rect 16396 21564 16448 21616
rect 17316 21564 17368 21616
rect 20444 21632 20496 21684
rect 18604 21607 18656 21616
rect 18604 21573 18613 21607
rect 18613 21573 18647 21607
rect 18647 21573 18656 21607
rect 18604 21564 18656 21573
rect 20168 21564 20220 21616
rect 22008 21632 22060 21684
rect 22376 21632 22428 21684
rect 23756 21632 23808 21684
rect 23940 21632 23992 21684
rect 24216 21632 24268 21684
rect 12624 21428 12676 21480
rect 12716 21471 12768 21480
rect 12716 21437 12725 21471
rect 12725 21437 12759 21471
rect 12759 21437 12768 21471
rect 12716 21428 12768 21437
rect 14372 21428 14424 21480
rect 16028 21428 16080 21480
rect 1308 21292 1360 21344
rect 6092 21292 6144 21344
rect 6460 21335 6512 21344
rect 6460 21301 6469 21335
rect 6469 21301 6503 21335
rect 6503 21301 6512 21335
rect 6460 21292 6512 21301
rect 6644 21335 6696 21344
rect 6644 21301 6653 21335
rect 6653 21301 6687 21335
rect 6687 21301 6696 21335
rect 6644 21292 6696 21301
rect 7564 21292 7616 21344
rect 9588 21292 9640 21344
rect 10692 21335 10744 21344
rect 10692 21301 10701 21335
rect 10701 21301 10735 21335
rect 10735 21301 10744 21335
rect 10692 21292 10744 21301
rect 11612 21335 11664 21344
rect 11612 21301 11621 21335
rect 11621 21301 11655 21335
rect 11655 21301 11664 21335
rect 11612 21292 11664 21301
rect 11704 21335 11756 21344
rect 11704 21301 11713 21335
rect 11713 21301 11747 21335
rect 11747 21301 11756 21335
rect 11704 21292 11756 21301
rect 12072 21292 12124 21344
rect 13452 21360 13504 21412
rect 16212 21360 16264 21412
rect 15292 21292 15344 21344
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 18236 21496 18288 21548
rect 18328 21539 18380 21548
rect 18328 21505 18337 21539
rect 18337 21505 18371 21539
rect 18371 21505 18380 21539
rect 18328 21496 18380 21505
rect 16488 21428 16540 21480
rect 16948 21428 17000 21480
rect 17408 21471 17460 21480
rect 17408 21437 17417 21471
rect 17417 21437 17451 21471
rect 17451 21437 17460 21471
rect 17408 21428 17460 21437
rect 17040 21360 17092 21412
rect 18328 21360 18380 21412
rect 19708 21360 19760 21412
rect 17868 21292 17920 21344
rect 18972 21292 19024 21344
rect 21640 21564 21692 21616
rect 23572 21607 23624 21616
rect 23572 21573 23581 21607
rect 23581 21573 23615 21607
rect 23615 21573 23624 21607
rect 23572 21564 23624 21573
rect 20076 21471 20128 21480
rect 20076 21437 20085 21471
rect 20085 21437 20119 21471
rect 20119 21437 20128 21471
rect 20076 21428 20128 21437
rect 21180 21471 21232 21480
rect 21180 21437 21189 21471
rect 21189 21437 21223 21471
rect 21223 21437 21232 21471
rect 21180 21428 21232 21437
rect 21456 21496 21508 21548
rect 22100 21496 22152 21548
rect 21364 21428 21416 21480
rect 22284 21428 22336 21480
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 23296 21539 23348 21548
rect 23296 21505 23305 21539
rect 23305 21505 23339 21539
rect 23339 21505 23348 21539
rect 23296 21496 23348 21505
rect 23020 21428 23072 21480
rect 23572 21428 23624 21480
rect 19892 21360 19944 21412
rect 21732 21360 21784 21412
rect 21824 21360 21876 21412
rect 23112 21360 23164 21412
rect 25596 21360 25648 21412
rect 26056 21360 26108 21412
rect 20168 21292 20220 21344
rect 21548 21292 21600 21344
rect 23388 21292 23440 21344
rect 25320 21292 25372 21344
rect 25504 21292 25556 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 3976 21088 4028 21140
rect 6828 21088 6880 21140
rect 7380 21088 7432 21140
rect 3332 21020 3384 21072
rect 5724 21020 5776 21072
rect 2780 20995 2832 21004
rect 2780 20961 2789 20995
rect 2789 20961 2823 20995
rect 2823 20961 2832 20995
rect 2780 20952 2832 20961
rect 4160 20952 4212 21004
rect 4620 20952 4672 21004
rect 6828 20952 6880 21004
rect 2228 20927 2280 20936
rect 2228 20893 2237 20927
rect 2237 20893 2271 20927
rect 2271 20893 2280 20927
rect 2228 20884 2280 20893
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 2504 20816 2556 20868
rect 4712 20816 4764 20868
rect 6460 20884 6512 20936
rect 10048 21020 10100 21072
rect 15660 21088 15712 21140
rect 18604 21088 18656 21140
rect 18696 21088 18748 21140
rect 21364 21088 21416 21140
rect 7288 20952 7340 21004
rect 7748 20884 7800 20936
rect 9588 20952 9640 21004
rect 9680 20952 9732 21004
rect 12716 21020 12768 21072
rect 8760 20927 8812 20936
rect 8760 20893 8769 20927
rect 8769 20893 8803 20927
rect 8803 20893 8812 20927
rect 10600 20995 10652 21004
rect 10600 20961 10609 20995
rect 10609 20961 10643 20995
rect 10643 20961 10652 20995
rect 10600 20952 10652 20961
rect 11520 20952 11572 21004
rect 12624 20952 12676 21004
rect 8760 20884 8812 20893
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 13728 20927 13780 20936
rect 13728 20893 13737 20927
rect 13737 20893 13771 20927
rect 13771 20893 13780 20927
rect 13728 20884 13780 20893
rect 2044 20748 2096 20800
rect 2780 20748 2832 20800
rect 3516 20748 3568 20800
rect 5540 20748 5592 20800
rect 6000 20748 6052 20800
rect 12716 20816 12768 20868
rect 13176 20816 13228 20868
rect 13268 20816 13320 20868
rect 14372 20884 14424 20936
rect 14464 20884 14516 20936
rect 14004 20816 14056 20868
rect 15384 20884 15436 20936
rect 16028 20884 16080 20936
rect 16488 20884 16540 20936
rect 17224 21020 17276 21072
rect 17776 20952 17828 21004
rect 19248 21020 19300 21072
rect 21272 21020 21324 21072
rect 18328 20952 18380 21004
rect 19064 20952 19116 21004
rect 20260 20952 20312 21004
rect 20444 20952 20496 21004
rect 21640 21020 21692 21072
rect 22284 21088 22336 21140
rect 25228 21088 25280 21140
rect 22468 20952 22520 21004
rect 22928 20952 22980 21004
rect 23572 20952 23624 21004
rect 16948 20927 17000 20936
rect 16948 20893 16957 20927
rect 16957 20893 16991 20927
rect 16991 20893 17000 20927
rect 16948 20884 17000 20893
rect 21364 20884 21416 20936
rect 16764 20816 16816 20868
rect 9956 20791 10008 20800
rect 9956 20757 9965 20791
rect 9965 20757 9999 20791
rect 9999 20757 10008 20791
rect 9956 20748 10008 20757
rect 11152 20748 11204 20800
rect 15844 20748 15896 20800
rect 16856 20791 16908 20800
rect 16856 20757 16865 20791
rect 16865 20757 16899 20791
rect 16899 20757 16908 20791
rect 16856 20748 16908 20757
rect 17684 20791 17736 20800
rect 17684 20757 17693 20791
rect 17693 20757 17727 20791
rect 17727 20757 17736 20791
rect 17684 20748 17736 20757
rect 18236 20816 18288 20868
rect 19064 20791 19116 20800
rect 19064 20757 19073 20791
rect 19073 20757 19107 20791
rect 19107 20757 19116 20791
rect 19064 20748 19116 20757
rect 19708 20859 19760 20868
rect 19708 20825 19717 20859
rect 19717 20825 19751 20859
rect 19751 20825 19760 20859
rect 19708 20816 19760 20825
rect 20720 20816 20772 20868
rect 24676 21020 24728 21072
rect 24952 21020 25004 21072
rect 24584 20884 24636 20936
rect 21640 20748 21692 20800
rect 21732 20791 21784 20800
rect 21732 20757 21741 20791
rect 21741 20757 21775 20791
rect 21775 20757 21784 20791
rect 21732 20748 21784 20757
rect 22284 20748 22336 20800
rect 22560 20791 22612 20800
rect 22560 20757 22569 20791
rect 22569 20757 22603 20791
rect 22603 20757 22612 20791
rect 22560 20748 22612 20757
rect 22652 20748 22704 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 25412 20748 25464 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 4436 20544 4488 20596
rect 4712 20587 4764 20596
rect 4712 20553 4721 20587
rect 4721 20553 4755 20587
rect 4755 20553 4764 20587
rect 4712 20544 4764 20553
rect 6000 20587 6052 20596
rect 6000 20553 6009 20587
rect 6009 20553 6043 20587
rect 6043 20553 6052 20587
rect 6000 20544 6052 20553
rect 8484 20587 8536 20596
rect 8484 20553 8493 20587
rect 8493 20553 8527 20587
rect 8527 20553 8536 20587
rect 8484 20544 8536 20553
rect 7288 20476 7340 20528
rect 11060 20519 11112 20528
rect 11060 20485 11069 20519
rect 11069 20485 11103 20519
rect 11103 20485 11112 20519
rect 11060 20476 11112 20485
rect 11244 20476 11296 20528
rect 13268 20519 13320 20528
rect 13268 20485 13277 20519
rect 13277 20485 13311 20519
rect 13311 20485 13320 20519
rect 13268 20476 13320 20485
rect 2964 20340 3016 20392
rect 5080 20408 5132 20460
rect 6000 20408 6052 20460
rect 6552 20408 6604 20460
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 8944 20451 8996 20460
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 10968 20408 11020 20460
rect 5632 20340 5684 20392
rect 8300 20340 8352 20392
rect 9680 20340 9732 20392
rect 2320 20272 2372 20324
rect 3700 20272 3752 20324
rect 3976 20272 4028 20324
rect 8852 20272 8904 20324
rect 4252 20204 4304 20256
rect 5080 20204 5132 20256
rect 6552 20204 6604 20256
rect 7840 20204 7892 20256
rect 11980 20272 12032 20324
rect 10508 20204 10560 20256
rect 11244 20204 11296 20256
rect 11704 20247 11756 20256
rect 11704 20213 11713 20247
rect 11713 20213 11747 20247
rect 11747 20213 11756 20247
rect 11704 20204 11756 20213
rect 12072 20247 12124 20256
rect 12072 20213 12081 20247
rect 12081 20213 12115 20247
rect 12115 20213 12124 20247
rect 12072 20204 12124 20213
rect 12624 20383 12676 20392
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 12624 20340 12676 20349
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13544 20476 13596 20528
rect 15384 20587 15436 20596
rect 15384 20553 15393 20587
rect 15393 20553 15427 20587
rect 15427 20553 15436 20587
rect 15384 20544 15436 20553
rect 14004 20476 14056 20528
rect 16488 20519 16540 20528
rect 16488 20485 16497 20519
rect 16497 20485 16531 20519
rect 16531 20485 16540 20519
rect 16488 20476 16540 20485
rect 16948 20476 17000 20528
rect 13636 20451 13688 20460
rect 13176 20408 13228 20417
rect 13636 20417 13652 20451
rect 13652 20417 13686 20451
rect 13686 20417 13688 20451
rect 13636 20408 13688 20417
rect 17040 20408 17092 20460
rect 17408 20383 17460 20392
rect 17408 20349 17417 20383
rect 17417 20349 17451 20383
rect 17451 20349 17460 20383
rect 17408 20340 17460 20349
rect 18420 20340 18472 20392
rect 20168 20476 20220 20528
rect 20628 20544 20680 20596
rect 22376 20587 22428 20596
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 23112 20587 23164 20596
rect 23112 20553 23121 20587
rect 23121 20553 23155 20587
rect 23155 20553 23164 20587
rect 23112 20544 23164 20553
rect 21732 20476 21784 20528
rect 24216 20476 24268 20528
rect 25320 20476 25372 20528
rect 25596 20476 25648 20528
rect 19340 20408 19392 20460
rect 19432 20340 19484 20392
rect 20904 20408 20956 20460
rect 21180 20408 21232 20460
rect 22008 20408 22060 20460
rect 23296 20408 23348 20460
rect 21088 20340 21140 20392
rect 21272 20383 21324 20392
rect 21272 20349 21281 20383
rect 21281 20349 21315 20383
rect 21315 20349 21324 20383
rect 21272 20340 21324 20349
rect 21916 20340 21968 20392
rect 13544 20204 13596 20256
rect 17132 20272 17184 20324
rect 20168 20272 20220 20324
rect 22652 20383 22704 20392
rect 22652 20349 22661 20383
rect 22661 20349 22695 20383
rect 22695 20349 22704 20383
rect 22652 20340 22704 20349
rect 23756 20383 23808 20392
rect 23756 20349 23765 20383
rect 23765 20349 23799 20383
rect 23799 20349 23808 20383
rect 23756 20340 23808 20349
rect 18512 20204 18564 20256
rect 18972 20204 19024 20256
rect 19340 20247 19392 20256
rect 19340 20213 19349 20247
rect 19349 20213 19383 20247
rect 19383 20213 19392 20247
rect 19340 20204 19392 20213
rect 19616 20204 19668 20256
rect 20076 20204 20128 20256
rect 21272 20204 21324 20256
rect 23572 20204 23624 20256
rect 25136 20204 25188 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 3884 20000 3936 20052
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 7472 20000 7524 20052
rect 7656 20000 7708 20052
rect 9404 20000 9456 20052
rect 4160 19932 4212 19984
rect 4344 19932 4396 19984
rect 9956 20000 10008 20052
rect 17132 20000 17184 20052
rect 21824 20000 21876 20052
rect 4528 19796 4580 19848
rect 5632 19864 5684 19916
rect 8668 19864 8720 19916
rect 6736 19796 6788 19848
rect 6828 19839 6880 19848
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 10876 19907 10928 19916
rect 10876 19873 10885 19907
rect 10885 19873 10919 19907
rect 10919 19873 10928 19907
rect 10876 19864 10928 19873
rect 13452 19932 13504 19984
rect 13728 19975 13780 19984
rect 13728 19941 13737 19975
rect 13737 19941 13771 19975
rect 13771 19941 13780 19975
rect 13728 19932 13780 19941
rect 13912 19975 13964 19984
rect 13912 19941 13921 19975
rect 13921 19941 13955 19975
rect 13955 19941 13964 19975
rect 13912 19932 13964 19941
rect 15108 19932 15160 19984
rect 3976 19728 4028 19780
rect 10692 19796 10744 19848
rect 11520 19839 11572 19848
rect 11520 19805 11529 19839
rect 11529 19805 11563 19839
rect 11563 19805 11572 19839
rect 11520 19796 11572 19805
rect 13360 19796 13412 19848
rect 15016 19864 15068 19916
rect 13820 19728 13872 19780
rect 14740 19796 14792 19848
rect 22284 20000 22336 20052
rect 23204 20000 23256 20052
rect 22376 19932 22428 19984
rect 23112 19932 23164 19984
rect 23480 19932 23532 19984
rect 15568 19864 15620 19916
rect 16764 19864 16816 19916
rect 17132 19864 17184 19916
rect 18328 19907 18380 19916
rect 18328 19873 18337 19907
rect 18337 19873 18371 19907
rect 18371 19873 18380 19907
rect 18328 19864 18380 19873
rect 19064 19864 19116 19916
rect 23296 19864 23348 19916
rect 24400 19864 24452 19916
rect 16028 19796 16080 19848
rect 16488 19796 16540 19848
rect 17224 19796 17276 19848
rect 17592 19796 17644 19848
rect 18880 19796 18932 19848
rect 20536 19796 20588 19848
rect 22468 19796 22520 19848
rect 22928 19796 22980 19848
rect 4528 19660 4580 19712
rect 5356 19660 5408 19712
rect 5724 19660 5776 19712
rect 8392 19660 8444 19712
rect 9220 19660 9272 19712
rect 9956 19660 10008 19712
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 10416 19660 10468 19712
rect 14372 19728 14424 19780
rect 14004 19660 14056 19712
rect 14924 19703 14976 19712
rect 14924 19669 14933 19703
rect 14933 19669 14967 19703
rect 14967 19669 14976 19703
rect 14924 19660 14976 19669
rect 15016 19660 15068 19712
rect 18512 19728 18564 19780
rect 16488 19703 16540 19712
rect 16488 19669 16497 19703
rect 16497 19669 16531 19703
rect 16531 19669 16540 19703
rect 16488 19660 16540 19669
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 18696 19660 18748 19712
rect 21180 19771 21232 19780
rect 21180 19737 21189 19771
rect 21189 19737 21223 19771
rect 21223 19737 21232 19771
rect 21180 19728 21232 19737
rect 18972 19703 19024 19712
rect 18972 19669 18981 19703
rect 18981 19669 19015 19703
rect 19015 19669 19024 19703
rect 18972 19660 19024 19669
rect 19524 19660 19576 19712
rect 20444 19703 20496 19712
rect 20444 19669 20453 19703
rect 20453 19669 20487 19703
rect 20487 19669 20496 19703
rect 20444 19660 20496 19669
rect 20720 19660 20772 19712
rect 21456 19660 21508 19712
rect 23020 19660 23072 19712
rect 23204 19660 23256 19712
rect 23756 19660 23808 19712
rect 24584 19703 24636 19712
rect 24584 19669 24593 19703
rect 24593 19669 24627 19703
rect 24627 19669 24636 19703
rect 24584 19660 24636 19669
rect 25320 19660 25372 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 4068 19456 4120 19508
rect 1492 19388 1544 19440
rect 5632 19456 5684 19508
rect 6000 19499 6052 19508
rect 6000 19465 6009 19499
rect 6009 19465 6043 19499
rect 6043 19465 6052 19499
rect 6000 19456 6052 19465
rect 6736 19456 6788 19508
rect 7472 19456 7524 19508
rect 1952 19363 2004 19372
rect 1952 19329 1961 19363
rect 1961 19329 1995 19363
rect 1995 19329 2004 19363
rect 1952 19320 2004 19329
rect 4160 19320 4212 19372
rect 6276 19388 6328 19440
rect 6920 19388 6972 19440
rect 10692 19499 10744 19508
rect 10692 19465 10701 19499
rect 10701 19465 10735 19499
rect 10735 19465 10744 19499
rect 10692 19456 10744 19465
rect 11520 19456 11572 19508
rect 5356 19363 5408 19372
rect 5356 19329 5365 19363
rect 5365 19329 5399 19363
rect 5399 19329 5408 19363
rect 5356 19320 5408 19329
rect 6644 19320 6696 19372
rect 7472 19320 7524 19372
rect 7656 19320 7708 19372
rect 7840 19363 7892 19372
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 8944 19363 8996 19372
rect 8944 19329 8953 19363
rect 8953 19329 8987 19363
rect 8987 19329 8996 19363
rect 8944 19320 8996 19329
rect 10324 19320 10376 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 14280 19456 14332 19508
rect 14740 19499 14792 19508
rect 14740 19465 14749 19499
rect 14749 19465 14783 19499
rect 14783 19465 14792 19499
rect 14740 19456 14792 19465
rect 14832 19456 14884 19508
rect 15108 19456 15160 19508
rect 17684 19456 17736 19508
rect 12808 19431 12860 19440
rect 12808 19397 12817 19431
rect 12817 19397 12851 19431
rect 12851 19397 12860 19431
rect 12808 19388 12860 19397
rect 13912 19320 13964 19372
rect 16948 19388 17000 19440
rect 19616 19499 19668 19508
rect 19616 19465 19625 19499
rect 19625 19465 19659 19499
rect 19659 19465 19668 19499
rect 19616 19456 19668 19465
rect 20996 19456 21048 19508
rect 21364 19456 21416 19508
rect 22560 19456 22612 19508
rect 25228 19456 25280 19508
rect 26516 19456 26568 19508
rect 21456 19388 21508 19440
rect 1584 19252 1636 19304
rect 2596 19252 2648 19304
rect 4528 19252 4580 19304
rect 11060 19252 11112 19304
rect 12256 19252 12308 19304
rect 4160 19184 4212 19236
rect 5264 19184 5316 19236
rect 7012 19184 7064 19236
rect 8760 19184 8812 19236
rect 7288 19116 7340 19168
rect 13360 19252 13412 19304
rect 13452 19252 13504 19304
rect 15108 19363 15160 19372
rect 15108 19329 15117 19363
rect 15117 19329 15151 19363
rect 15151 19329 15160 19363
rect 15108 19320 15160 19329
rect 15384 19320 15436 19372
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 20720 19320 20772 19372
rect 21088 19320 21140 19372
rect 21640 19320 21692 19372
rect 22284 19320 22336 19372
rect 14096 19252 14148 19304
rect 13360 19116 13412 19168
rect 14464 19116 14516 19168
rect 15016 19116 15068 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 16396 19116 16448 19168
rect 16672 19116 16724 19168
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 20904 19252 20956 19304
rect 19984 19184 20036 19236
rect 23112 19320 23164 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 22560 19252 22612 19304
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 23940 19252 23992 19304
rect 24768 19252 24820 19304
rect 25228 19252 25280 19304
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 20812 19116 20864 19168
rect 21640 19116 21692 19168
rect 22928 19184 22980 19236
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 4804 18912 4856 18964
rect 9496 18912 9548 18964
rect 12348 18912 12400 18964
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 3976 18708 4028 18760
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 6368 18708 6420 18760
rect 6644 18708 6696 18760
rect 6828 18751 6880 18760
rect 6828 18717 6837 18751
rect 6837 18717 6871 18751
rect 6871 18717 6880 18751
rect 6828 18708 6880 18717
rect 12072 18844 12124 18896
rect 12256 18844 12308 18896
rect 12992 18887 13044 18896
rect 12992 18853 13001 18887
rect 13001 18853 13035 18887
rect 13035 18853 13044 18887
rect 12992 18844 13044 18853
rect 13176 18844 13228 18896
rect 13728 18844 13780 18896
rect 14372 18912 14424 18964
rect 15568 18844 15620 18896
rect 9312 18776 9364 18828
rect 10968 18776 11020 18828
rect 12624 18776 12676 18828
rect 10140 18708 10192 18760
rect 12256 18708 12308 18760
rect 13084 18708 13136 18760
rect 2228 18572 2280 18624
rect 3424 18615 3476 18624
rect 3424 18581 3433 18615
rect 3433 18581 3467 18615
rect 3467 18581 3476 18615
rect 3424 18572 3476 18581
rect 5632 18640 5684 18692
rect 6000 18640 6052 18692
rect 9496 18640 9548 18692
rect 13452 18819 13504 18828
rect 13452 18785 13461 18819
rect 13461 18785 13495 18819
rect 13495 18785 13504 18819
rect 13452 18776 13504 18785
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 13820 18776 13872 18828
rect 19064 18912 19116 18964
rect 19892 18912 19944 18964
rect 23664 18912 23716 18964
rect 17592 18844 17644 18896
rect 19340 18844 19392 18896
rect 21640 18844 21692 18896
rect 21916 18844 21968 18896
rect 22652 18844 22704 18896
rect 23388 18844 23440 18896
rect 26608 18844 26660 18896
rect 16304 18776 16356 18828
rect 16856 18776 16908 18828
rect 14004 18708 14056 18760
rect 14280 18708 14332 18760
rect 17500 18776 17552 18828
rect 20260 18819 20312 18828
rect 20260 18785 20269 18819
rect 20269 18785 20303 18819
rect 20303 18785 20312 18819
rect 20260 18776 20312 18785
rect 20536 18819 20588 18828
rect 20536 18785 20545 18819
rect 20545 18785 20579 18819
rect 20579 18785 20588 18819
rect 20536 18776 20588 18785
rect 20628 18776 20680 18828
rect 18788 18708 18840 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 13360 18683 13412 18692
rect 13360 18649 13369 18683
rect 13369 18649 13403 18683
rect 13403 18649 13412 18683
rect 13360 18640 13412 18649
rect 14832 18640 14884 18692
rect 16580 18640 16632 18692
rect 5264 18615 5316 18624
rect 5264 18581 5273 18615
rect 5273 18581 5307 18615
rect 5307 18581 5316 18615
rect 5264 18572 5316 18581
rect 5816 18572 5868 18624
rect 6184 18572 6236 18624
rect 6368 18615 6420 18624
rect 6368 18581 6377 18615
rect 6377 18581 6411 18615
rect 6411 18581 6420 18615
rect 6368 18572 6420 18581
rect 7012 18572 7064 18624
rect 7840 18572 7892 18624
rect 11336 18572 11388 18624
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 12348 18572 12400 18624
rect 16672 18572 16724 18624
rect 16856 18572 16908 18624
rect 19156 18640 19208 18692
rect 17592 18615 17644 18624
rect 17592 18581 17601 18615
rect 17601 18581 17635 18615
rect 17635 18581 17644 18615
rect 17592 18572 17644 18581
rect 17776 18572 17828 18624
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 18420 18572 18472 18581
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 18788 18572 18840 18624
rect 20812 18640 20864 18692
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 21456 18572 21508 18624
rect 22744 18708 22796 18760
rect 22836 18708 22888 18760
rect 25044 18819 25096 18828
rect 25044 18785 25053 18819
rect 25053 18785 25087 18819
rect 25087 18785 25096 18819
rect 25044 18776 25096 18785
rect 25136 18819 25188 18828
rect 25136 18785 25145 18819
rect 25145 18785 25179 18819
rect 25179 18785 25188 18819
rect 25136 18776 25188 18785
rect 25320 18708 25372 18760
rect 22192 18640 22244 18692
rect 21916 18572 21968 18624
rect 22652 18572 22704 18624
rect 24676 18640 24728 18692
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 1676 18368 1728 18420
rect 6000 18411 6052 18420
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 6184 18368 6236 18420
rect 6828 18368 6880 18420
rect 14096 18368 14148 18420
rect 14280 18411 14332 18420
rect 14280 18377 14289 18411
rect 14289 18377 14323 18411
rect 14323 18377 14332 18411
rect 14280 18368 14332 18377
rect 14832 18368 14884 18420
rect 16120 18368 16172 18420
rect 16672 18411 16724 18420
rect 16672 18377 16681 18411
rect 16681 18377 16715 18411
rect 16715 18377 16724 18411
rect 16672 18368 16724 18377
rect 5264 18300 5316 18352
rect 12256 18300 12308 18352
rect 18328 18300 18380 18352
rect 18420 18300 18472 18352
rect 18880 18300 18932 18352
rect 20260 18300 20312 18352
rect 20536 18368 20588 18420
rect 22468 18368 22520 18420
rect 23296 18411 23348 18420
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 25872 18368 25924 18420
rect 3884 18232 3936 18284
rect 4252 18275 4304 18284
rect 4252 18241 4261 18275
rect 4261 18241 4295 18275
rect 4295 18241 4304 18275
rect 4252 18232 4304 18241
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 5356 18232 5408 18241
rect 6920 18232 6972 18284
rect 7380 18164 7432 18216
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 10324 18232 10376 18284
rect 10508 18232 10560 18284
rect 11152 18232 11204 18284
rect 13084 18232 13136 18284
rect 13820 18232 13872 18284
rect 14188 18232 14240 18284
rect 6920 18096 6972 18148
rect 11060 18164 11112 18216
rect 11796 18164 11848 18216
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 12624 18164 12676 18216
rect 13268 18164 13320 18216
rect 13452 18164 13504 18216
rect 15660 18164 15712 18216
rect 15752 18164 15804 18216
rect 17132 18232 17184 18284
rect 19432 18232 19484 18284
rect 20536 18232 20588 18284
rect 20812 18275 20864 18284
rect 20812 18241 20821 18275
rect 20821 18241 20855 18275
rect 20855 18241 20864 18275
rect 20812 18232 20864 18241
rect 21088 18232 21140 18284
rect 25320 18343 25372 18352
rect 25320 18309 25329 18343
rect 25329 18309 25363 18343
rect 25363 18309 25372 18343
rect 25320 18300 25372 18309
rect 25596 18232 25648 18284
rect 25872 18232 25924 18284
rect 16120 18207 16172 18216
rect 16120 18173 16129 18207
rect 16129 18173 16163 18207
rect 16163 18173 16172 18207
rect 16120 18164 16172 18173
rect 16488 18164 16540 18216
rect 17592 18164 17644 18216
rect 17776 18164 17828 18216
rect 17868 18164 17920 18216
rect 20720 18164 20772 18216
rect 16396 18096 16448 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 7380 18071 7432 18080
rect 7380 18037 7389 18071
rect 7389 18037 7423 18071
rect 7423 18037 7432 18071
rect 7380 18028 7432 18037
rect 8484 18071 8536 18080
rect 8484 18037 8493 18071
rect 8493 18037 8527 18071
rect 8527 18037 8536 18071
rect 8484 18028 8536 18037
rect 8668 18028 8720 18080
rect 9312 18028 9364 18080
rect 11520 18028 11572 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 12256 18028 12308 18080
rect 13176 18028 13228 18080
rect 13912 18028 13964 18080
rect 14648 18028 14700 18080
rect 15660 18028 15712 18080
rect 16488 18028 16540 18080
rect 18420 18028 18472 18080
rect 19156 18096 19208 18148
rect 24768 18096 24820 18148
rect 19524 18028 19576 18080
rect 20628 18028 20680 18080
rect 22928 18028 22980 18080
rect 24400 18028 24452 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 3976 17799 4028 17808
rect 3976 17765 3985 17799
rect 3985 17765 4019 17799
rect 4019 17765 4028 17799
rect 3976 17756 4028 17765
rect 4620 17824 4672 17876
rect 5356 17824 5408 17876
rect 6920 17824 6972 17876
rect 7380 17824 7432 17876
rect 6736 17756 6788 17808
rect 3424 17688 3476 17740
rect 8208 17756 8260 17808
rect 9128 17756 9180 17808
rect 11244 17867 11296 17876
rect 11244 17833 11253 17867
rect 11253 17833 11287 17867
rect 11287 17833 11296 17867
rect 11244 17824 11296 17833
rect 12072 17824 12124 17876
rect 12348 17824 12400 17876
rect 12440 17824 12492 17876
rect 13544 17824 13596 17876
rect 15752 17824 15804 17876
rect 15844 17824 15896 17876
rect 16580 17824 16632 17876
rect 16948 17824 17000 17876
rect 17224 17824 17276 17876
rect 17408 17824 17460 17876
rect 17592 17824 17644 17876
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 3792 17620 3844 17672
rect 8300 17688 8352 17740
rect 8852 17688 8904 17740
rect 8944 17688 8996 17740
rect 3424 17595 3476 17604
rect 3424 17561 3433 17595
rect 3433 17561 3467 17595
rect 3467 17561 3476 17595
rect 3424 17552 3476 17561
rect 5724 17663 5776 17672
rect 5724 17629 5733 17663
rect 5733 17629 5767 17663
rect 5767 17629 5776 17663
rect 5724 17620 5776 17629
rect 6184 17620 6236 17672
rect 7656 17620 7708 17672
rect 8668 17620 8720 17672
rect 9036 17596 9088 17648
rect 11704 17731 11756 17740
rect 11704 17697 11713 17731
rect 11713 17697 11747 17731
rect 11747 17697 11756 17731
rect 11704 17688 11756 17697
rect 19432 17756 19484 17808
rect 22100 17756 22152 17808
rect 22192 17756 22244 17808
rect 22836 17799 22888 17808
rect 22836 17765 22845 17799
rect 22845 17765 22879 17799
rect 22879 17765 22888 17799
rect 22836 17756 22888 17765
rect 12072 17688 12124 17740
rect 12440 17688 12492 17740
rect 12624 17688 12676 17740
rect 14188 17688 14240 17740
rect 14280 17688 14332 17740
rect 15292 17688 15344 17740
rect 16764 17688 16816 17740
rect 18604 17688 18656 17740
rect 18880 17731 18932 17740
rect 18880 17697 18889 17731
rect 18889 17697 18923 17731
rect 18923 17697 18932 17731
rect 18880 17688 18932 17697
rect 13636 17620 13688 17672
rect 14740 17620 14792 17672
rect 10324 17552 10376 17604
rect 2044 17484 2096 17536
rect 5908 17484 5960 17536
rect 7472 17527 7524 17536
rect 7472 17493 7481 17527
rect 7481 17493 7515 17527
rect 7515 17493 7524 17527
rect 7472 17484 7524 17493
rect 8576 17484 8628 17536
rect 9220 17484 9272 17536
rect 9588 17484 9640 17536
rect 10508 17484 10560 17536
rect 12072 17552 12124 17604
rect 13268 17552 13320 17604
rect 13360 17552 13412 17604
rect 15844 17552 15896 17604
rect 11244 17484 11296 17536
rect 16672 17552 16724 17604
rect 16948 17484 17000 17536
rect 19064 17620 19116 17672
rect 21640 17688 21692 17740
rect 24032 17688 24084 17740
rect 19984 17663 20036 17672
rect 19984 17629 19993 17663
rect 19993 17629 20027 17663
rect 20027 17629 20036 17663
rect 19984 17620 20036 17629
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 24492 17620 24544 17672
rect 18420 17552 18472 17604
rect 20996 17595 21048 17604
rect 20996 17561 21005 17595
rect 21005 17561 21039 17595
rect 21039 17561 21048 17595
rect 20996 17552 21048 17561
rect 21456 17552 21508 17604
rect 23848 17552 23900 17604
rect 22284 17484 22336 17536
rect 23296 17527 23348 17536
rect 23296 17493 23305 17527
rect 23305 17493 23339 17527
rect 23339 17493 23348 17527
rect 23296 17484 23348 17493
rect 24952 17484 25004 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 2688 17323 2740 17332
rect 2688 17289 2697 17323
rect 2697 17289 2731 17323
rect 2731 17289 2740 17323
rect 2688 17280 2740 17289
rect 3792 17323 3844 17332
rect 3792 17289 3801 17323
rect 3801 17289 3835 17323
rect 3835 17289 3844 17323
rect 3792 17280 3844 17289
rect 6460 17323 6512 17332
rect 6460 17289 6469 17323
rect 6469 17289 6503 17323
rect 6503 17289 6512 17323
rect 6460 17280 6512 17289
rect 7288 17280 7340 17332
rect 7380 17280 7432 17332
rect 7656 17323 7708 17332
rect 7656 17289 7665 17323
rect 7665 17289 7699 17323
rect 7699 17289 7708 17323
rect 7656 17280 7708 17289
rect 6736 17212 6788 17264
rect 3424 17144 3476 17196
rect 4252 17187 4304 17196
rect 4252 17153 4261 17187
rect 4261 17153 4295 17187
rect 4295 17153 4304 17187
rect 4252 17144 4304 17153
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 7012 17187 7064 17196
rect 7012 17153 7021 17187
rect 7021 17153 7055 17187
rect 7055 17153 7064 17187
rect 7012 17144 7064 17153
rect 7472 17212 7524 17264
rect 10508 17212 10560 17264
rect 11336 17280 11388 17332
rect 14648 17280 14700 17332
rect 14188 17212 14240 17264
rect 15476 17280 15528 17332
rect 15568 17280 15620 17332
rect 8484 17144 8536 17196
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 14096 17144 14148 17196
rect 5908 17076 5960 17128
rect 7196 17076 7248 17128
rect 5632 17008 5684 17060
rect 7840 17008 7892 17060
rect 8116 17008 8168 17060
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 6000 16940 6052 16949
rect 6736 16983 6788 16992
rect 6736 16949 6745 16983
rect 6745 16949 6779 16983
rect 6779 16949 6788 16983
rect 6736 16940 6788 16949
rect 9220 16940 9272 16992
rect 9496 17076 9548 17128
rect 10692 17008 10744 17060
rect 11244 17051 11296 17060
rect 11244 17017 11253 17051
rect 11253 17017 11287 17051
rect 11287 17017 11296 17051
rect 11244 17008 11296 17017
rect 10600 16940 10652 16992
rect 10968 16983 11020 16992
rect 10968 16949 10977 16983
rect 10977 16949 11011 16983
rect 11011 16949 11020 16983
rect 10968 16940 11020 16949
rect 11704 17076 11756 17128
rect 12072 17051 12124 17060
rect 12072 17017 12081 17051
rect 12081 17017 12115 17051
rect 12115 17017 12124 17051
rect 12072 17008 12124 17017
rect 12440 17008 12492 17060
rect 13360 17076 13412 17128
rect 13452 17076 13504 17128
rect 16672 17212 16724 17264
rect 18604 17212 18656 17264
rect 18696 17255 18748 17264
rect 18696 17221 18705 17255
rect 18705 17221 18739 17255
rect 18739 17221 18748 17255
rect 18696 17212 18748 17221
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 20812 17280 20864 17332
rect 15476 17144 15528 17196
rect 16028 17144 16080 17196
rect 17592 17144 17644 17196
rect 18420 17187 18472 17196
rect 18420 17153 18429 17187
rect 18429 17153 18463 17187
rect 18463 17153 18472 17187
rect 18420 17144 18472 17153
rect 19800 17144 19852 17196
rect 21456 17212 21508 17264
rect 26240 17212 26292 17264
rect 26792 17212 26844 17264
rect 20720 17144 20772 17196
rect 22468 17187 22520 17196
rect 22468 17153 22477 17187
rect 22477 17153 22511 17187
rect 22511 17153 22520 17187
rect 22468 17144 22520 17153
rect 23848 17144 23900 17196
rect 24768 17144 24820 17196
rect 15844 17076 15896 17128
rect 16212 17076 16264 17128
rect 16856 17076 16908 17128
rect 14004 16940 14056 16992
rect 14648 16940 14700 16992
rect 16672 16940 16724 16992
rect 17132 17008 17184 17060
rect 17960 17076 18012 17128
rect 19064 17076 19116 17128
rect 21456 17076 21508 17128
rect 22100 17076 22152 17128
rect 22836 17076 22888 17128
rect 24032 17076 24084 17128
rect 20536 17008 20588 17060
rect 17408 16940 17460 16992
rect 21456 16940 21508 16992
rect 22008 16983 22060 16992
rect 22008 16949 22017 16983
rect 22017 16949 22051 16983
rect 22051 16949 22060 16983
rect 22008 16940 22060 16949
rect 22100 16983 22152 16992
rect 22100 16949 22109 16983
rect 22109 16949 22143 16983
rect 22143 16949 22152 16983
rect 22100 16940 22152 16949
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 4528 16736 4580 16788
rect 9036 16736 9088 16788
rect 4068 16600 4120 16652
rect 2688 16532 2740 16584
rect 3516 16532 3568 16584
rect 4436 16532 4488 16584
rect 5264 16575 5316 16584
rect 5264 16541 5273 16575
rect 5273 16541 5307 16575
rect 5307 16541 5316 16575
rect 5264 16532 5316 16541
rect 6184 16532 6236 16584
rect 6276 16532 6328 16584
rect 8852 16668 8904 16720
rect 9496 16736 9548 16788
rect 23204 16736 23256 16788
rect 9680 16668 9732 16720
rect 8668 16600 8720 16652
rect 8760 16600 8812 16652
rect 2320 16439 2372 16448
rect 2320 16405 2329 16439
rect 2329 16405 2363 16439
rect 2363 16405 2372 16439
rect 2320 16396 2372 16405
rect 2412 16396 2464 16448
rect 4068 16464 4120 16516
rect 5172 16464 5224 16516
rect 7104 16464 7156 16516
rect 8116 16464 8168 16516
rect 8208 16464 8260 16516
rect 8484 16464 8536 16516
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 14004 16668 14056 16720
rect 13728 16600 13780 16652
rect 9220 16464 9272 16516
rect 11704 16532 11756 16584
rect 13360 16532 13412 16584
rect 14096 16600 14148 16652
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 16028 16711 16080 16720
rect 16028 16677 16037 16711
rect 16037 16677 16071 16711
rect 16071 16677 16080 16711
rect 16028 16668 16080 16677
rect 16120 16668 16172 16720
rect 16304 16668 16356 16720
rect 21548 16668 21600 16720
rect 22192 16668 22244 16720
rect 16856 16600 16908 16652
rect 17868 16600 17920 16652
rect 18420 16600 18472 16652
rect 18788 16600 18840 16652
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 23664 16668 23716 16720
rect 24768 16600 24820 16652
rect 25688 16600 25740 16652
rect 16948 16532 17000 16584
rect 22008 16532 22060 16584
rect 23940 16532 23992 16584
rect 4896 16396 4948 16448
rect 4988 16396 5040 16448
rect 8300 16396 8352 16448
rect 8576 16439 8628 16448
rect 8576 16405 8585 16439
rect 8585 16405 8619 16439
rect 8619 16405 8628 16439
rect 8576 16396 8628 16405
rect 11888 16464 11940 16516
rect 12256 16507 12308 16516
rect 12256 16473 12265 16507
rect 12265 16473 12299 16507
rect 12299 16473 12308 16507
rect 12256 16464 12308 16473
rect 15844 16464 15896 16516
rect 9496 16396 9548 16448
rect 10508 16396 10560 16448
rect 10600 16396 10652 16448
rect 11152 16439 11204 16448
rect 11152 16405 11161 16439
rect 11161 16405 11195 16439
rect 11195 16405 11204 16439
rect 11152 16396 11204 16405
rect 12164 16396 12216 16448
rect 14648 16396 14700 16448
rect 17684 16464 17736 16516
rect 18788 16396 18840 16448
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 19708 16507 19760 16516
rect 19708 16473 19717 16507
rect 19717 16473 19751 16507
rect 19751 16473 19760 16507
rect 19708 16464 19760 16473
rect 19800 16396 19852 16448
rect 23848 16464 23900 16516
rect 20996 16396 21048 16448
rect 21732 16396 21784 16448
rect 22192 16396 22244 16448
rect 22744 16396 22796 16448
rect 24032 16439 24084 16448
rect 24032 16405 24041 16439
rect 24041 16405 24075 16439
rect 24075 16405 24084 16439
rect 24032 16396 24084 16405
rect 24216 16396 24268 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 4252 16192 4304 16244
rect 5264 16192 5316 16244
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 2688 16124 2740 16176
rect 5172 16124 5224 16176
rect 5724 16124 5776 16176
rect 7932 16192 7984 16244
rect 8668 16192 8720 16244
rect 8944 16192 8996 16244
rect 10600 16192 10652 16244
rect 12256 16192 12308 16244
rect 13452 16235 13504 16244
rect 13452 16201 13461 16235
rect 13461 16201 13495 16235
rect 13495 16201 13504 16235
rect 13452 16192 13504 16201
rect 13728 16192 13780 16244
rect 18328 16235 18380 16244
rect 18328 16201 18337 16235
rect 18337 16201 18371 16235
rect 18371 16201 18380 16235
rect 18328 16192 18380 16201
rect 18788 16192 18840 16244
rect 20260 16192 20312 16244
rect 20812 16235 20864 16244
rect 20812 16201 20821 16235
rect 20821 16201 20855 16235
rect 20855 16201 20864 16235
rect 20812 16192 20864 16201
rect 21180 16192 21232 16244
rect 21456 16192 21508 16244
rect 21732 16192 21784 16244
rect 3332 16056 3384 16108
rect 6460 16056 6512 16108
rect 6736 16099 6788 16108
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 6736 16056 6788 16065
rect 6828 16056 6880 16108
rect 10968 16124 11020 16176
rect 11888 16124 11940 16176
rect 13360 16124 13412 16176
rect 13912 16124 13964 16176
rect 14832 16124 14884 16176
rect 7012 15988 7064 16040
rect 8300 16099 8352 16108
rect 8300 16065 8309 16099
rect 8309 16065 8343 16099
rect 8343 16065 8352 16099
rect 8300 16056 8352 16065
rect 9680 16056 9732 16108
rect 10140 16056 10192 16108
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 13544 16056 13596 16108
rect 13820 16056 13872 16108
rect 14924 16056 14976 16108
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 16304 16124 16356 16176
rect 18420 16124 18472 16176
rect 19524 16124 19576 16176
rect 19708 16124 19760 16176
rect 22560 16124 22612 16176
rect 23480 16192 23532 16244
rect 25688 16124 25740 16176
rect 9496 15988 9548 16040
rect 11152 15988 11204 16040
rect 12348 15988 12400 16040
rect 14096 15988 14148 16040
rect 5632 15920 5684 15972
rect 6736 15920 6788 15972
rect 7196 15920 7248 15972
rect 8760 15920 8812 15972
rect 15108 15988 15160 16040
rect 19064 16056 19116 16108
rect 15936 16031 15988 16040
rect 15936 15997 15945 16031
rect 15945 15997 15979 16031
rect 15979 15997 15988 16031
rect 15936 15988 15988 15997
rect 16396 15988 16448 16040
rect 19616 15988 19668 16040
rect 20812 16056 20864 16108
rect 22744 16056 22796 16108
rect 24124 16056 24176 16108
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 3884 15852 3936 15904
rect 4896 15852 4948 15904
rect 7472 15852 7524 15904
rect 7932 15852 7984 15904
rect 9956 15852 10008 15904
rect 10416 15852 10468 15904
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 16304 15920 16356 15972
rect 16488 15852 16540 15904
rect 16948 15852 17000 15904
rect 17040 15852 17092 15904
rect 21088 16031 21140 16040
rect 21088 15997 21097 16031
rect 21097 15997 21131 16031
rect 21131 15997 21140 16031
rect 21088 15988 21140 15997
rect 21180 15988 21232 16040
rect 21916 15988 21968 16040
rect 24032 16031 24084 16040
rect 24032 15997 24041 16031
rect 24041 15997 24075 16031
rect 24075 15997 24084 16031
rect 24032 15988 24084 15997
rect 24308 15988 24360 16040
rect 22008 15895 22060 15904
rect 22008 15861 22017 15895
rect 22017 15861 22051 15895
rect 22051 15861 22060 15895
rect 22008 15852 22060 15861
rect 23664 15920 23716 15972
rect 23388 15895 23440 15904
rect 23388 15861 23397 15895
rect 23397 15861 23431 15895
rect 23431 15861 23440 15895
rect 23388 15852 23440 15861
rect 25228 15895 25280 15904
rect 25228 15861 25237 15895
rect 25237 15861 25271 15895
rect 25271 15861 25280 15895
rect 25228 15852 25280 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 4160 15648 4212 15700
rect 7564 15648 7616 15700
rect 10416 15648 10468 15700
rect 2136 15623 2188 15632
rect 2136 15589 2145 15623
rect 2145 15589 2179 15623
rect 2179 15589 2188 15623
rect 2136 15580 2188 15589
rect 2596 15580 2648 15632
rect 7196 15580 7248 15632
rect 9680 15580 9732 15632
rect 11704 15580 11756 15632
rect 12256 15580 12308 15632
rect 12716 15580 12768 15632
rect 13728 15648 13780 15700
rect 13820 15691 13872 15700
rect 13820 15657 13829 15691
rect 13829 15657 13863 15691
rect 13863 15657 13872 15691
rect 13820 15648 13872 15657
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 4252 15512 4304 15564
rect 7748 15512 7800 15564
rect 1492 15376 1544 15428
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 6000 15444 6052 15496
rect 9128 15512 9180 15564
rect 8576 15444 8628 15496
rect 4712 15376 4764 15428
rect 8668 15376 8720 15428
rect 10600 15512 10652 15564
rect 12164 15444 12216 15496
rect 13636 15580 13688 15632
rect 14556 15648 14608 15700
rect 14740 15648 14792 15700
rect 16580 15691 16632 15700
rect 16580 15657 16589 15691
rect 16589 15657 16623 15691
rect 16623 15657 16632 15691
rect 16580 15648 16632 15657
rect 16488 15580 16540 15632
rect 17592 15648 17644 15700
rect 20904 15648 20956 15700
rect 21456 15648 21508 15700
rect 22376 15648 22428 15700
rect 23020 15648 23072 15700
rect 24584 15648 24636 15700
rect 18880 15580 18932 15632
rect 13820 15512 13872 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 19616 15512 19668 15564
rect 19984 15512 20036 15564
rect 20076 15555 20128 15564
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 23940 15580 23992 15632
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 4436 15308 4488 15360
rect 4896 15308 4948 15360
rect 5264 15351 5316 15360
rect 5264 15317 5273 15351
rect 5273 15317 5307 15351
rect 5307 15317 5316 15351
rect 5264 15308 5316 15317
rect 7564 15308 7616 15360
rect 7932 15308 7984 15360
rect 8300 15308 8352 15360
rect 10508 15308 10560 15360
rect 11888 15376 11940 15428
rect 11980 15376 12032 15428
rect 14096 15444 14148 15496
rect 16304 15444 16356 15496
rect 12440 15308 12492 15360
rect 12716 15308 12768 15360
rect 13728 15308 13780 15360
rect 14372 15308 14424 15360
rect 14556 15419 14608 15428
rect 14556 15385 14565 15419
rect 14565 15385 14599 15419
rect 14599 15385 14608 15419
rect 14556 15376 14608 15385
rect 16672 15376 16724 15428
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 16120 15308 16172 15360
rect 17684 15376 17736 15428
rect 20812 15444 20864 15496
rect 21456 15512 21508 15564
rect 19432 15419 19484 15428
rect 19432 15385 19441 15419
rect 19441 15385 19475 15419
rect 19475 15385 19484 15419
rect 19432 15376 19484 15385
rect 20168 15376 20220 15428
rect 19064 15351 19116 15360
rect 19064 15317 19073 15351
rect 19073 15317 19107 15351
rect 19107 15317 19116 15351
rect 19064 15308 19116 15317
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 19800 15308 19852 15360
rect 20996 15376 21048 15428
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 22192 15444 22244 15496
rect 22468 15444 22520 15496
rect 24216 15444 24268 15496
rect 25780 15376 25832 15428
rect 26424 15376 26476 15428
rect 24124 15351 24176 15360
rect 24124 15317 24133 15351
rect 24133 15317 24167 15351
rect 24167 15317 24176 15351
rect 24124 15308 24176 15317
rect 25504 15308 25556 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 2596 15104 2648 15156
rect 5908 15104 5960 15156
rect 6276 15104 6328 15156
rect 7288 15104 7340 15156
rect 7656 15104 7708 15156
rect 1860 15036 1912 15088
rect 2136 15036 2188 15088
rect 2228 15036 2280 15088
rect 4160 14968 4212 15020
rect 1952 14900 2004 14952
rect 3792 14900 3844 14952
rect 1676 14832 1728 14884
rect 4528 14968 4580 15020
rect 5448 14968 5500 15020
rect 8576 14968 8628 15020
rect 13820 15104 13872 15156
rect 15568 15147 15620 15156
rect 15568 15113 15577 15147
rect 15577 15113 15611 15147
rect 15611 15113 15620 15147
rect 15568 15104 15620 15113
rect 9956 15036 10008 15088
rect 10876 15036 10928 15088
rect 11152 15079 11204 15088
rect 11152 15045 11161 15079
rect 11161 15045 11195 15079
rect 11195 15045 11204 15079
rect 11152 15036 11204 15045
rect 12164 15079 12216 15088
rect 12164 15045 12173 15079
rect 12173 15045 12207 15079
rect 12207 15045 12216 15079
rect 12164 15036 12216 15045
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 12532 14968 12584 15020
rect 13268 15036 13320 15088
rect 13452 15036 13504 15088
rect 14740 14968 14792 15020
rect 9036 14900 9088 14952
rect 9496 14900 9548 14952
rect 11244 14900 11296 14952
rect 1860 14764 1912 14816
rect 3516 14764 3568 14816
rect 7748 14832 7800 14884
rect 9220 14832 9272 14884
rect 12164 14832 12216 14884
rect 7564 14764 7616 14816
rect 9680 14764 9732 14816
rect 10876 14764 10928 14816
rect 14832 14900 14884 14952
rect 14096 14832 14148 14884
rect 17960 15104 18012 15156
rect 16120 15079 16172 15088
rect 16120 15045 16129 15079
rect 16129 15045 16163 15079
rect 16163 15045 16172 15079
rect 16120 15036 16172 15045
rect 14280 14764 14332 14816
rect 14740 14764 14792 14816
rect 17040 15036 17092 15088
rect 17684 15036 17736 15088
rect 25136 15104 25188 15156
rect 20076 15036 20128 15088
rect 21456 15079 21508 15088
rect 21456 15045 21465 15079
rect 21465 15045 21499 15079
rect 21499 15045 21508 15079
rect 21456 15036 21508 15045
rect 22376 15036 22428 15088
rect 23572 15036 23624 15088
rect 21548 14968 21600 15020
rect 22284 14968 22336 15020
rect 25596 14968 25648 15020
rect 16488 14832 16540 14884
rect 17224 14900 17276 14952
rect 19340 14943 19392 14952
rect 16580 14764 16632 14816
rect 16856 14764 16908 14816
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 18880 14832 18932 14884
rect 22652 14900 22704 14952
rect 23388 14900 23440 14952
rect 24400 14900 24452 14952
rect 20720 14764 20772 14816
rect 21548 14807 21600 14816
rect 21548 14773 21557 14807
rect 21557 14773 21591 14807
rect 21591 14773 21600 14807
rect 21548 14764 21600 14773
rect 22468 14832 22520 14884
rect 22744 14832 22796 14884
rect 23020 14764 23072 14816
rect 24584 14764 24636 14816
rect 25044 14764 25096 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 1584 14356 1636 14408
rect 3976 14560 4028 14612
rect 5724 14560 5776 14612
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 9220 14603 9272 14612
rect 9220 14569 9229 14603
rect 9229 14569 9263 14603
rect 9263 14569 9272 14603
rect 9220 14560 9272 14569
rect 5264 14492 5316 14544
rect 2320 14424 2372 14476
rect 2688 14356 2740 14408
rect 4068 14356 4120 14408
rect 4436 14356 4488 14408
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 5172 14356 5224 14408
rect 6368 14467 6420 14476
rect 6368 14433 6377 14467
rect 6377 14433 6411 14467
rect 6411 14433 6420 14467
rect 6368 14424 6420 14433
rect 7288 14424 7340 14476
rect 8944 14424 8996 14476
rect 8300 14356 8352 14408
rect 9680 14492 9732 14544
rect 12164 14560 12216 14612
rect 12348 14535 12400 14544
rect 10600 14467 10652 14476
rect 10600 14433 10609 14467
rect 10609 14433 10643 14467
rect 10643 14433 10652 14467
rect 10600 14424 10652 14433
rect 12348 14501 12357 14535
rect 12357 14501 12391 14535
rect 12391 14501 12400 14535
rect 12348 14492 12400 14501
rect 12532 14560 12584 14612
rect 13544 14560 13596 14612
rect 15752 14560 15804 14612
rect 16028 14603 16080 14612
rect 16028 14569 16037 14603
rect 16037 14569 16071 14603
rect 16071 14569 16080 14603
rect 16028 14560 16080 14569
rect 16764 14560 16816 14612
rect 17408 14560 17460 14612
rect 17776 14560 17828 14612
rect 18604 14560 18656 14612
rect 21916 14560 21968 14612
rect 22100 14560 22152 14612
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 10968 14424 11020 14476
rect 14096 14424 14148 14476
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 15200 14424 15252 14476
rect 11888 14356 11940 14408
rect 12256 14356 12308 14408
rect 2320 14288 2372 14340
rect 3516 14288 3568 14340
rect 5816 14288 5868 14340
rect 6552 14288 6604 14340
rect 1584 14220 1636 14272
rect 3976 14263 4028 14272
rect 3976 14229 3985 14263
rect 3985 14229 4019 14263
rect 4019 14229 4028 14263
rect 3976 14220 4028 14229
rect 7840 14220 7892 14272
rect 8944 14220 8996 14272
rect 9220 14220 9272 14272
rect 12716 14288 12768 14340
rect 13176 14356 13228 14408
rect 13360 14288 13412 14340
rect 14648 14288 14700 14340
rect 15016 14288 15068 14340
rect 14096 14220 14148 14272
rect 15936 14424 15988 14476
rect 16212 14424 16264 14476
rect 17868 14492 17920 14544
rect 21456 14492 21508 14544
rect 19800 14424 19852 14476
rect 20720 14424 20772 14476
rect 22008 14424 22060 14476
rect 23388 14424 23440 14476
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 20444 14356 20496 14408
rect 22836 14356 22888 14408
rect 24032 14424 24084 14476
rect 25412 14356 25464 14408
rect 16580 14220 16632 14272
rect 17040 14288 17092 14340
rect 18328 14288 18380 14340
rect 24492 14288 24544 14340
rect 25320 14288 25372 14340
rect 17776 14220 17828 14272
rect 18420 14220 18472 14272
rect 19800 14263 19852 14272
rect 19800 14229 19809 14263
rect 19809 14229 19843 14263
rect 19843 14229 19852 14263
rect 19800 14220 19852 14229
rect 20444 14263 20496 14272
rect 20444 14229 20453 14263
rect 20453 14229 20487 14263
rect 20487 14229 20496 14263
rect 20444 14220 20496 14229
rect 21916 14220 21968 14272
rect 23020 14263 23072 14272
rect 23020 14229 23029 14263
rect 23029 14229 23063 14263
rect 23063 14229 23072 14263
rect 23020 14220 23072 14229
rect 23388 14263 23440 14272
rect 23388 14229 23397 14263
rect 23397 14229 23431 14263
rect 23431 14229 23440 14263
rect 23388 14220 23440 14229
rect 24124 14220 24176 14272
rect 24768 14220 24820 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 1308 14016 1360 14068
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 4160 13948 4212 14000
rect 8300 14016 8352 14068
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 4896 13923 4948 13932
rect 4896 13889 4905 13923
rect 4905 13889 4939 13923
rect 4939 13889 4948 13923
rect 4896 13880 4948 13889
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 9128 13948 9180 14000
rect 10600 14016 10652 14068
rect 10968 14016 11020 14068
rect 11244 14016 11296 14068
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 9220 13880 9272 13932
rect 10416 13948 10468 14000
rect 5724 13812 5776 13864
rect 6368 13812 6420 13864
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 10324 13812 10376 13864
rect 12624 13948 12676 14000
rect 11152 13880 11204 13932
rect 12348 13880 12400 13932
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 11428 13812 11480 13864
rect 13728 14016 13780 14068
rect 14280 14016 14332 14068
rect 14556 14016 14608 14068
rect 17868 14059 17920 14068
rect 17868 14025 17877 14059
rect 17877 14025 17911 14059
rect 17911 14025 17920 14059
rect 17868 14016 17920 14025
rect 18604 14016 18656 14068
rect 19340 14016 19392 14068
rect 20352 14059 20404 14068
rect 20352 14025 20361 14059
rect 20361 14025 20395 14059
rect 20395 14025 20404 14059
rect 20352 14016 20404 14025
rect 21824 14016 21876 14068
rect 24032 14059 24084 14068
rect 24032 14025 24041 14059
rect 24041 14025 24075 14059
rect 24075 14025 24084 14059
rect 24032 14016 24084 14025
rect 24216 14016 24268 14068
rect 25136 14059 25188 14068
rect 25136 14025 25145 14059
rect 25145 14025 25179 14059
rect 25179 14025 25188 14059
rect 25136 14016 25188 14025
rect 15660 13948 15712 14000
rect 18328 13948 18380 14000
rect 21364 13948 21416 14000
rect 21916 13948 21968 14000
rect 23572 13948 23624 14000
rect 15016 13880 15068 13932
rect 14556 13812 14608 13864
rect 15108 13812 15160 13864
rect 16304 13880 16356 13932
rect 16580 13880 16632 13932
rect 20720 13880 20772 13932
rect 17040 13812 17092 13864
rect 17684 13812 17736 13864
rect 18328 13812 18380 13864
rect 20076 13812 20128 13864
rect 21272 13855 21324 13864
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 21732 13812 21784 13864
rect 22284 13923 22336 13932
rect 22284 13889 22293 13923
rect 22293 13889 22327 13923
rect 22327 13889 22336 13923
rect 22284 13880 22336 13889
rect 23848 13880 23900 13932
rect 23756 13812 23808 13864
rect 25596 13812 25648 13864
rect 3332 13744 3384 13796
rect 4528 13744 4580 13796
rect 4712 13744 4764 13796
rect 7288 13744 7340 13796
rect 10784 13744 10836 13796
rect 11520 13744 11572 13796
rect 12624 13744 12676 13796
rect 13636 13744 13688 13796
rect 15844 13744 15896 13796
rect 18420 13744 18472 13796
rect 20904 13744 20956 13796
rect 21180 13744 21232 13796
rect 3976 13676 4028 13728
rect 6092 13676 6144 13728
rect 9312 13676 9364 13728
rect 11152 13676 11204 13728
rect 15108 13676 15160 13728
rect 15200 13676 15252 13728
rect 21364 13676 21416 13728
rect 25412 13676 25464 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 2412 13472 2464 13524
rect 2504 13472 2556 13524
rect 2964 13472 3016 13524
rect 3240 13515 3292 13524
rect 3240 13481 3249 13515
rect 3249 13481 3283 13515
rect 3283 13481 3292 13515
rect 3240 13472 3292 13481
rect 4160 13472 4212 13524
rect 4712 13472 4764 13524
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 4436 13404 4488 13456
rect 2136 13336 2188 13388
rect 4252 13379 4304 13388
rect 4252 13345 4261 13379
rect 4261 13345 4295 13379
rect 4295 13345 4304 13379
rect 4252 13336 4304 13345
rect 6736 13472 6788 13524
rect 7012 13472 7064 13524
rect 8944 13515 8996 13524
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 6092 13404 6144 13456
rect 1308 13268 1360 13320
rect 2872 13268 2924 13320
rect 2320 13200 2372 13252
rect 2964 13243 3016 13252
rect 2964 13209 2973 13243
rect 2973 13209 3007 13243
rect 3007 13209 3016 13243
rect 2964 13200 3016 13209
rect 3792 13200 3844 13252
rect 5632 13336 5684 13388
rect 9128 13404 9180 13456
rect 10140 13472 10192 13524
rect 10600 13472 10652 13524
rect 11520 13472 11572 13524
rect 12624 13472 12676 13524
rect 14832 13472 14884 13524
rect 17132 13472 17184 13524
rect 17868 13472 17920 13524
rect 6460 13268 6512 13320
rect 9956 13336 10008 13388
rect 10048 13336 10100 13388
rect 10600 13336 10652 13388
rect 7104 13268 7156 13320
rect 9588 13268 9640 13320
rect 5172 13200 5224 13252
rect 7196 13200 7248 13252
rect 11152 13200 11204 13252
rect 12256 13200 12308 13252
rect 18788 13404 18840 13456
rect 21180 13404 21232 13456
rect 21364 13404 21416 13456
rect 23480 13472 23532 13524
rect 23940 13472 23992 13524
rect 24676 13472 24728 13524
rect 26884 13472 26936 13524
rect 14464 13336 14516 13388
rect 15384 13336 15436 13388
rect 16672 13336 16724 13388
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 14740 13268 14792 13320
rect 15016 13268 15068 13320
rect 17040 13268 17092 13320
rect 6000 13132 6052 13184
rect 6644 13132 6696 13184
rect 7012 13132 7064 13184
rect 9496 13132 9548 13184
rect 11060 13132 11112 13184
rect 13268 13132 13320 13184
rect 13452 13132 13504 13184
rect 13912 13132 13964 13184
rect 16212 13200 16264 13252
rect 15384 13175 15436 13184
rect 15384 13141 15393 13175
rect 15393 13141 15427 13175
rect 15427 13141 15436 13175
rect 15384 13132 15436 13141
rect 15476 13132 15528 13184
rect 16672 13132 16724 13184
rect 19340 13336 19392 13388
rect 21916 13379 21968 13388
rect 21916 13345 21925 13379
rect 21925 13345 21959 13379
rect 21959 13345 21968 13379
rect 21916 13336 21968 13345
rect 23572 13336 23624 13388
rect 26240 13404 26292 13456
rect 25228 13336 25280 13388
rect 24952 13268 25004 13320
rect 18512 13200 18564 13252
rect 19524 13200 19576 13252
rect 19984 13243 20036 13252
rect 19984 13209 19993 13243
rect 19993 13209 20027 13243
rect 20027 13209 20036 13243
rect 19984 13200 20036 13209
rect 18328 13175 18380 13184
rect 18328 13141 18337 13175
rect 18337 13141 18371 13175
rect 18371 13141 18380 13175
rect 18328 13132 18380 13141
rect 18972 13175 19024 13184
rect 18972 13141 18981 13175
rect 18981 13141 19015 13175
rect 19015 13141 19024 13175
rect 18972 13132 19024 13141
rect 19708 13132 19760 13184
rect 19892 13132 19944 13184
rect 20720 13132 20772 13184
rect 21456 13175 21508 13184
rect 21456 13141 21465 13175
rect 21465 13141 21499 13175
rect 21499 13141 21508 13175
rect 21456 13132 21508 13141
rect 23664 13200 23716 13252
rect 24768 13200 24820 13252
rect 25596 13200 25648 13252
rect 24584 13132 24636 13184
rect 24952 13132 25004 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 4620 12928 4672 12980
rect 4804 12928 4856 12980
rect 5172 12928 5224 12980
rect 5816 12971 5868 12980
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 6828 12928 6880 12980
rect 4896 12860 4948 12912
rect 6184 12860 6236 12912
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 11704 12928 11756 12980
rect 13912 12928 13964 12980
rect 14280 12928 14332 12980
rect 7932 12860 7984 12912
rect 3608 12792 3660 12844
rect 6828 12792 6880 12844
rect 6920 12792 6972 12844
rect 8944 12792 8996 12844
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 10232 12792 10284 12844
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 11060 12860 11112 12912
rect 12440 12860 12492 12912
rect 15016 12971 15068 12980
rect 15016 12937 15025 12971
rect 15025 12937 15059 12971
rect 15059 12937 15068 12971
rect 15016 12928 15068 12937
rect 15384 12928 15436 12980
rect 15936 12928 15988 12980
rect 16580 12928 16632 12980
rect 18972 12928 19024 12980
rect 17132 12860 17184 12912
rect 19156 12860 19208 12912
rect 19524 12928 19576 12980
rect 11520 12792 11572 12844
rect 12164 12835 12216 12844
rect 12164 12801 12173 12835
rect 12173 12801 12207 12835
rect 12207 12801 12216 12835
rect 12164 12792 12216 12801
rect 12624 12792 12676 12844
rect 13176 12792 13228 12844
rect 14648 12792 14700 12844
rect 16304 12792 16356 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 2780 12724 2832 12776
rect 7472 12767 7524 12776
rect 7472 12733 7481 12767
rect 7481 12733 7515 12767
rect 7515 12733 7524 12767
rect 7472 12724 7524 12733
rect 10048 12724 10100 12776
rect 7288 12656 7340 12708
rect 11428 12656 11480 12708
rect 11520 12656 11572 12708
rect 12256 12656 12308 12708
rect 14648 12656 14700 12708
rect 15752 12724 15804 12776
rect 17684 12724 17736 12776
rect 18604 12767 18656 12776
rect 18604 12733 18613 12767
rect 18613 12733 18647 12767
rect 18647 12733 18656 12767
rect 20260 12860 20312 12912
rect 20628 12928 20680 12980
rect 21180 12928 21232 12980
rect 21732 12928 21784 12980
rect 22376 12928 22428 12980
rect 22836 12928 22888 12980
rect 23480 12928 23532 12980
rect 24492 12928 24544 12980
rect 20444 12860 20496 12912
rect 20996 12860 21048 12912
rect 22928 12860 22980 12912
rect 23664 12860 23716 12912
rect 18604 12724 18656 12733
rect 6092 12588 6144 12640
rect 6552 12588 6604 12640
rect 6828 12588 6880 12640
rect 15200 12588 15252 12640
rect 21732 12792 21784 12844
rect 21916 12792 21968 12844
rect 24032 12792 24084 12844
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 19156 12588 19208 12640
rect 21180 12724 21232 12776
rect 20536 12656 20588 12708
rect 26148 12724 26200 12776
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 20812 12588 20864 12640
rect 21456 12588 21508 12640
rect 21824 12588 21876 12640
rect 22008 12588 22060 12640
rect 22100 12588 22152 12640
rect 22376 12588 22428 12640
rect 22652 12631 22704 12640
rect 22652 12597 22676 12631
rect 22676 12597 22704 12631
rect 22652 12588 22704 12597
rect 25320 12588 25372 12640
rect 25964 12588 26016 12640
rect 26148 12588 26200 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 2780 12384 2832 12436
rect 10324 12384 10376 12436
rect 10508 12384 10560 12436
rect 12256 12384 12308 12436
rect 12532 12384 12584 12436
rect 13728 12384 13780 12436
rect 15108 12384 15160 12436
rect 21180 12427 21232 12436
rect 2228 12316 2280 12368
rect 848 12248 900 12300
rect 8392 12316 8444 12368
rect 9220 12316 9272 12368
rect 21180 12393 21189 12427
rect 21189 12393 21223 12427
rect 21223 12393 21232 12427
rect 21180 12384 21232 12393
rect 22100 12384 22152 12436
rect 24124 12384 24176 12436
rect 24492 12384 24544 12436
rect 25320 12384 25372 12436
rect 2504 12180 2556 12232
rect 4160 12180 4212 12232
rect 4620 12180 4672 12232
rect 5448 12180 5500 12232
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 5632 12112 5684 12164
rect 6460 12112 6512 12164
rect 5908 12044 5960 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 9404 12248 9456 12300
rect 7656 12180 7708 12232
rect 9128 12180 9180 12232
rect 7472 12112 7524 12164
rect 9588 12248 9640 12300
rect 10232 12180 10284 12232
rect 10968 12180 11020 12232
rect 11612 12248 11664 12300
rect 15292 12359 15344 12368
rect 15292 12325 15301 12359
rect 15301 12325 15335 12359
rect 15335 12325 15344 12359
rect 15292 12316 15344 12325
rect 15476 12316 15528 12368
rect 18328 12316 18380 12368
rect 18972 12316 19024 12368
rect 11796 12180 11848 12232
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 16764 12248 16816 12300
rect 16856 12248 16908 12300
rect 17040 12248 17092 12300
rect 20168 12248 20220 12300
rect 22836 12248 22888 12300
rect 24676 12248 24728 12300
rect 25044 12248 25096 12300
rect 25320 12248 25372 12300
rect 12992 12180 13044 12232
rect 13452 12180 13504 12232
rect 14556 12180 14608 12232
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 16672 12180 16724 12232
rect 18512 12180 18564 12232
rect 21272 12180 21324 12232
rect 21916 12180 21968 12232
rect 24124 12223 24176 12232
rect 24124 12189 24133 12223
rect 24133 12189 24167 12223
rect 24167 12189 24176 12223
rect 24124 12180 24176 12189
rect 24952 12180 25004 12232
rect 8392 12044 8444 12096
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 8852 12044 8904 12096
rect 11244 12044 11296 12096
rect 11612 12044 11664 12096
rect 13912 12044 13964 12096
rect 16120 12044 16172 12096
rect 16488 12044 16540 12096
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 19616 12112 19668 12164
rect 20720 12112 20772 12164
rect 23664 12112 23716 12164
rect 25596 12316 25648 12368
rect 25596 12112 25648 12164
rect 21548 12044 21600 12096
rect 23940 12044 23992 12096
rect 24124 12044 24176 12096
rect 24584 12044 24636 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 26332 11976 26384 12028
rect 2780 11840 2832 11892
rect 2872 11840 2924 11892
rect 664 11772 716 11824
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 2780 11704 2832 11756
rect 2872 11704 2924 11756
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 2228 11636 2280 11688
rect 8852 11840 8904 11892
rect 10140 11840 10192 11892
rect 10968 11883 11020 11892
rect 10968 11849 10977 11883
rect 10977 11849 11011 11883
rect 11011 11849 11020 11883
rect 10968 11840 11020 11849
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 11612 11840 11664 11892
rect 12164 11840 12216 11892
rect 14372 11840 14424 11892
rect 14924 11840 14976 11892
rect 16304 11883 16356 11892
rect 16304 11849 16313 11883
rect 16313 11849 16347 11883
rect 16347 11849 16356 11883
rect 16304 11840 16356 11849
rect 16488 11840 16540 11892
rect 17224 11840 17276 11892
rect 7656 11772 7708 11824
rect 8576 11772 8628 11824
rect 5908 11704 5960 11756
rect 1860 11611 1912 11620
rect 1860 11577 1869 11611
rect 1869 11577 1903 11611
rect 1903 11577 1912 11611
rect 1860 11568 1912 11577
rect 4344 11636 4396 11688
rect 5540 11636 5592 11688
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 10876 11704 10928 11756
rect 12348 11815 12400 11824
rect 12348 11781 12357 11815
rect 12357 11781 12391 11815
rect 12391 11781 12400 11815
rect 12348 11772 12400 11781
rect 21456 11840 21508 11892
rect 21640 11840 21692 11892
rect 9680 11636 9732 11688
rect 11796 11704 11848 11756
rect 18696 11772 18748 11824
rect 19892 11772 19944 11824
rect 13912 11747 13964 11756
rect 13912 11713 13921 11747
rect 13921 11713 13955 11747
rect 13955 11713 13964 11747
rect 13912 11704 13964 11713
rect 16028 11704 16080 11756
rect 16304 11704 16356 11756
rect 12992 11636 13044 11688
rect 15292 11568 15344 11620
rect 7748 11500 7800 11552
rect 8576 11543 8628 11552
rect 8576 11509 8585 11543
rect 8585 11509 8619 11543
rect 8619 11509 8628 11543
rect 8576 11500 8628 11509
rect 8852 11543 8904 11552
rect 8852 11509 8861 11543
rect 8861 11509 8895 11543
rect 8895 11509 8904 11543
rect 8852 11500 8904 11509
rect 9036 11500 9088 11552
rect 9588 11500 9640 11552
rect 16856 11636 16908 11688
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 18420 11704 18472 11756
rect 19340 11747 19392 11756
rect 19340 11713 19349 11747
rect 19349 11713 19383 11747
rect 19383 11713 19392 11747
rect 19340 11704 19392 11713
rect 20720 11704 20772 11756
rect 20904 11704 20956 11756
rect 21364 11704 21416 11756
rect 21640 11704 21692 11756
rect 25228 11840 25280 11892
rect 24860 11772 24912 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 22744 11704 22796 11756
rect 23940 11747 23992 11756
rect 23940 11713 23949 11747
rect 23949 11713 23983 11747
rect 23983 11713 23992 11747
rect 23940 11704 23992 11713
rect 24676 11704 24728 11756
rect 26700 11704 26752 11756
rect 16856 11500 16908 11552
rect 17684 11636 17736 11688
rect 18972 11636 19024 11688
rect 20352 11636 20404 11688
rect 18512 11568 18564 11620
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 19248 11500 19300 11552
rect 24952 11636 25004 11688
rect 20904 11568 20956 11620
rect 23480 11568 23532 11620
rect 21088 11543 21140 11552
rect 21088 11509 21097 11543
rect 21097 11509 21131 11543
rect 21131 11509 21140 11543
rect 21088 11500 21140 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 2780 11296 2832 11305
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 6736 11296 6788 11348
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 9864 11296 9916 11348
rect 7012 11228 7064 11280
rect 8576 11228 8628 11280
rect 9588 11228 9640 11280
rect 11980 11296 12032 11348
rect 13268 11296 13320 11348
rect 15660 11296 15712 11348
rect 19156 11296 19208 11348
rect 5816 11160 5868 11212
rect 7104 11160 7156 11212
rect 9680 11160 9732 11212
rect 10600 11160 10652 11212
rect 18512 11228 18564 11280
rect 13544 11160 13596 11212
rect 16948 11160 17000 11212
rect 1860 11092 1912 11144
rect 3792 11092 3844 11144
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 8852 11092 8904 11144
rect 10876 11092 10928 11144
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 2412 11067 2464 11076
rect 2412 11033 2421 11067
rect 2421 11033 2455 11067
rect 2455 11033 2464 11067
rect 2412 11024 2464 11033
rect 2504 11024 2556 11076
rect 9312 11024 9364 11076
rect 10600 11024 10652 11076
rect 12072 11067 12124 11076
rect 12072 11033 12081 11067
rect 12081 11033 12115 11067
rect 12115 11033 12124 11067
rect 12072 11024 12124 11033
rect 12624 11092 12676 11144
rect 13360 11092 13412 11144
rect 15016 11092 15068 11144
rect 17132 11160 17184 11212
rect 17408 11203 17460 11212
rect 17408 11169 17417 11203
rect 17417 11169 17451 11203
rect 17451 11169 17460 11203
rect 17408 11160 17460 11169
rect 17960 11160 18012 11212
rect 20536 11296 20588 11348
rect 21180 11339 21232 11348
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 19708 11228 19760 11280
rect 22560 11296 22612 11348
rect 21456 11228 21508 11280
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 20628 11092 20680 11144
rect 21456 11092 21508 11144
rect 14924 11024 14976 11076
rect 15108 11024 15160 11076
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 8760 10956 8812 11008
rect 11152 10956 11204 11008
rect 12164 10956 12216 11008
rect 12440 10956 12492 11008
rect 16856 10956 16908 11008
rect 16948 10956 17000 11008
rect 18420 11024 18472 11076
rect 19156 11024 19208 11076
rect 20168 11024 20220 11076
rect 20996 11024 21048 11076
rect 25044 11160 25096 11212
rect 21916 11135 21968 11144
rect 21916 11101 21925 11135
rect 21925 11101 21959 11135
rect 21959 11101 21968 11135
rect 21916 11092 21968 11101
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 25504 11092 25556 11144
rect 25228 11067 25280 11076
rect 25228 11033 25237 11067
rect 25237 11033 25271 11067
rect 25271 11033 25280 11067
rect 25228 11024 25280 11033
rect 17500 10956 17552 11008
rect 18052 10956 18104 11008
rect 18512 10999 18564 11008
rect 18512 10965 18521 10999
rect 18521 10965 18555 10999
rect 18555 10965 18564 10999
rect 18512 10956 18564 10965
rect 19248 10956 19300 11008
rect 24216 10956 24268 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 3700 10752 3752 10804
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 7656 10752 7708 10804
rect 12164 10752 12216 10804
rect 12256 10752 12308 10804
rect 3240 10684 3292 10736
rect 3976 10727 4028 10736
rect 3976 10693 3985 10727
rect 3985 10693 4019 10727
rect 4019 10693 4028 10727
rect 3976 10684 4028 10693
rect 11060 10684 11112 10736
rect 11152 10684 11204 10736
rect 13820 10752 13872 10804
rect 16672 10752 16724 10804
rect 17776 10752 17828 10804
rect 18972 10752 19024 10804
rect 1032 10548 1084 10600
rect 8944 10616 8996 10668
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 15476 10684 15528 10736
rect 17224 10684 17276 10736
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 17316 10616 17368 10668
rect 18512 10616 18564 10668
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 20444 10616 20496 10668
rect 21180 10752 21232 10804
rect 21732 10752 21784 10804
rect 26516 10752 26568 10804
rect 25136 10727 25188 10736
rect 25136 10693 25145 10727
rect 25145 10693 25179 10727
rect 25179 10693 25188 10727
rect 25136 10684 25188 10693
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 5172 10548 5224 10600
rect 940 10412 992 10464
rect 6460 10548 6512 10600
rect 14832 10548 14884 10600
rect 7840 10480 7892 10532
rect 8852 10480 8904 10532
rect 14464 10480 14516 10532
rect 16120 10480 16172 10532
rect 17776 10480 17828 10532
rect 20720 10480 20772 10532
rect 21548 10523 21600 10532
rect 21548 10489 21557 10523
rect 21557 10489 21591 10523
rect 21591 10489 21600 10523
rect 21548 10480 21600 10489
rect 21732 10548 21784 10600
rect 23664 10616 23716 10668
rect 24860 10548 24912 10600
rect 22100 10480 22152 10532
rect 3884 10412 3936 10464
rect 6460 10412 6512 10464
rect 11336 10412 11388 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 15660 10412 15712 10464
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 16948 10412 17000 10464
rect 18512 10412 18564 10464
rect 20076 10412 20128 10464
rect 21180 10412 21232 10464
rect 21824 10412 21876 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 1492 10208 1544 10260
rect 2320 10183 2372 10192
rect 2320 10149 2329 10183
rect 2329 10149 2363 10183
rect 2363 10149 2372 10183
rect 2320 10140 2372 10149
rect 4436 10140 4488 10192
rect 6552 10208 6604 10260
rect 9220 10208 9272 10260
rect 11612 10208 11664 10260
rect 12348 10208 12400 10260
rect 14004 10208 14056 10260
rect 18972 10251 19024 10260
rect 18972 10217 18981 10251
rect 18981 10217 19015 10251
rect 19015 10217 19024 10251
rect 18972 10208 19024 10217
rect 19340 10251 19392 10260
rect 19340 10217 19349 10251
rect 19349 10217 19383 10251
rect 19383 10217 19392 10251
rect 19340 10208 19392 10217
rect 23848 10208 23900 10260
rect 24216 10251 24268 10260
rect 24216 10217 24225 10251
rect 24225 10217 24259 10251
rect 24259 10217 24268 10251
rect 24216 10208 24268 10217
rect 10692 10140 10744 10192
rect 6460 10072 6512 10124
rect 2780 9979 2832 9988
rect 2780 9945 2789 9979
rect 2789 9945 2823 9979
rect 2823 9945 2832 9979
rect 2780 9936 2832 9945
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 6000 9936 6052 9988
rect 8392 9936 8444 9988
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 10416 10004 10468 10056
rect 10600 10004 10652 10056
rect 14004 10004 14056 10056
rect 16028 10072 16080 10124
rect 16212 10140 16264 10192
rect 21180 10140 21232 10192
rect 24124 10140 24176 10192
rect 16488 10072 16540 10124
rect 17132 10072 17184 10124
rect 20904 10072 20956 10124
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 25044 10115 25096 10124
rect 25044 10081 25053 10115
rect 25053 10081 25087 10115
rect 25087 10081 25096 10115
rect 25044 10072 25096 10081
rect 16580 10004 16632 10056
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 19248 10004 19300 10056
rect 20444 10004 20496 10056
rect 20720 10047 20772 10056
rect 20720 10013 20729 10047
rect 20729 10013 20763 10047
rect 20763 10013 20772 10047
rect 20720 10004 20772 10013
rect 5080 9868 5132 9920
rect 7748 9868 7800 9920
rect 8944 9868 8996 9920
rect 11336 9911 11388 9920
rect 11336 9877 11345 9911
rect 11345 9877 11379 9911
rect 11379 9877 11388 9911
rect 11336 9868 11388 9877
rect 19156 9936 19208 9988
rect 21824 9936 21876 9988
rect 13636 9868 13688 9920
rect 13728 9911 13780 9920
rect 13728 9877 13737 9911
rect 13737 9877 13771 9911
rect 13771 9877 13780 9911
rect 13728 9868 13780 9877
rect 17500 9868 17552 9920
rect 17868 9868 17920 9920
rect 21732 9868 21784 9920
rect 22928 9868 22980 9920
rect 23480 9936 23532 9988
rect 23756 9911 23808 9920
rect 23756 9877 23765 9911
rect 23765 9877 23799 9911
rect 23799 9877 23808 9911
rect 23756 9868 23808 9877
rect 24308 9868 24360 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 1124 9664 1176 9716
rect 7748 9664 7800 9716
rect 11796 9664 11848 9716
rect 14832 9664 14884 9716
rect 14924 9664 14976 9716
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 4620 9596 4672 9648
rect 4712 9639 4764 9648
rect 4712 9605 4721 9639
rect 4721 9605 4755 9639
rect 4755 9605 4764 9639
rect 4712 9596 4764 9605
rect 5172 9639 5224 9648
rect 5172 9605 5181 9639
rect 5181 9605 5215 9639
rect 5215 9605 5224 9639
rect 5172 9596 5224 9605
rect 8300 9596 8352 9648
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 14096 9596 14148 9648
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 11796 9528 11848 9580
rect 12348 9571 12400 9580
rect 12348 9537 12357 9571
rect 12357 9537 12391 9571
rect 12391 9537 12400 9571
rect 12348 9528 12400 9537
rect 14556 9571 14608 9580
rect 2136 9435 2188 9444
rect 2136 9401 2145 9435
rect 2145 9401 2179 9435
rect 2179 9401 2188 9435
rect 2136 9392 2188 9401
rect 2872 9392 2924 9444
rect 3516 9392 3568 9444
rect 7380 9460 7432 9512
rect 6368 9392 6420 9444
rect 10784 9460 10836 9512
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 14924 9528 14976 9580
rect 17684 9596 17736 9648
rect 16304 9528 16356 9580
rect 16948 9460 17000 9512
rect 17224 9528 17276 9580
rect 17868 9528 17920 9580
rect 17960 9528 18012 9580
rect 18604 9460 18656 9512
rect 19064 9664 19116 9716
rect 20168 9664 20220 9716
rect 20444 9707 20496 9716
rect 20444 9673 20453 9707
rect 20453 9673 20487 9707
rect 20487 9673 20496 9707
rect 20444 9664 20496 9673
rect 21180 9664 21232 9716
rect 19064 9528 19116 9580
rect 20628 9596 20680 9648
rect 20812 9528 20864 9580
rect 11612 9392 11664 9444
rect 11888 9392 11940 9444
rect 572 9324 624 9376
rect 3608 9324 3660 9376
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 5448 9324 5500 9376
rect 7564 9324 7616 9376
rect 12164 9324 12216 9376
rect 12716 9324 12768 9376
rect 16580 9324 16632 9376
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 17132 9324 17184 9376
rect 17316 9324 17368 9376
rect 18052 9392 18104 9444
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 24860 9596 24912 9648
rect 22652 9460 22704 9512
rect 22928 9460 22980 9512
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 21180 9435 21232 9444
rect 21180 9401 21189 9435
rect 21189 9401 21223 9435
rect 21223 9401 21232 9435
rect 21180 9392 21232 9401
rect 18604 9324 18656 9376
rect 19064 9367 19116 9376
rect 19064 9333 19073 9367
rect 19073 9333 19107 9367
rect 19107 9333 19116 9367
rect 19064 9324 19116 9333
rect 20444 9324 20496 9376
rect 20628 9324 20680 9376
rect 20812 9324 20864 9376
rect 23388 9324 23440 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 2504 9120 2556 9172
rect 3332 9120 3384 9172
rect 3608 9120 3660 9172
rect 5080 9052 5132 9104
rect 5724 9120 5776 9172
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 7840 9163 7892 9172
rect 7840 9129 7849 9163
rect 7849 9129 7883 9163
rect 7883 9129 7892 9163
rect 7840 9120 7892 9129
rect 7932 9120 7984 9172
rect 8668 9120 8720 9172
rect 8944 9163 8996 9172
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 11796 9120 11848 9172
rect 13268 9120 13320 9172
rect 13544 9120 13596 9172
rect 15108 9120 15160 9172
rect 16672 9120 16724 9172
rect 16856 9163 16908 9172
rect 16856 9129 16865 9163
rect 16865 9129 16899 9163
rect 16899 9129 16908 9163
rect 16856 9120 16908 9129
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 9496 9052 9548 9104
rect 756 8984 808 9036
rect 1584 8916 1636 8968
rect 2596 8916 2648 8968
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 2780 8916 2832 8925
rect 3608 8984 3660 9036
rect 4252 8984 4304 9036
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 7932 8984 7984 9036
rect 8484 8984 8536 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 14556 9052 14608 9104
rect 12624 8984 12676 9036
rect 15384 8984 15436 9036
rect 6276 8916 6328 8968
rect 6828 8916 6880 8968
rect 7840 8916 7892 8968
rect 8668 8916 8720 8968
rect 3884 8780 3936 8832
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 4712 8823 4764 8832
rect 4712 8789 4721 8823
rect 4721 8789 4755 8823
rect 4755 8789 4764 8823
rect 4712 8780 4764 8789
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 8852 8780 8904 8832
rect 11428 8916 11480 8968
rect 12164 8916 12216 8968
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 15108 8959 15160 8968
rect 15108 8925 15117 8959
rect 15117 8925 15151 8959
rect 15151 8925 15160 8959
rect 15108 8916 15160 8925
rect 15660 8916 15712 8968
rect 16672 8916 16724 8968
rect 17224 8916 17276 8968
rect 17316 8959 17368 8968
rect 17316 8925 17325 8959
rect 17325 8925 17359 8959
rect 17359 8925 17368 8959
rect 17316 8916 17368 8925
rect 10324 8891 10376 8900
rect 10324 8857 10333 8891
rect 10333 8857 10367 8891
rect 10367 8857 10376 8891
rect 10324 8848 10376 8857
rect 11612 8848 11664 8900
rect 18052 8848 18104 8900
rect 19064 9120 19116 9172
rect 19892 9120 19944 9172
rect 22100 9120 22152 9172
rect 25780 9120 25832 9172
rect 18604 9052 18656 9104
rect 19064 8984 19116 9036
rect 18604 8916 18656 8968
rect 19616 8984 19668 9036
rect 11704 8780 11756 8832
rect 13636 8780 13688 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 17592 8780 17644 8832
rect 21824 8823 21876 8832
rect 21824 8789 21833 8823
rect 21833 8789 21867 8823
rect 21867 8789 21876 8823
rect 21824 8780 21876 8789
rect 25228 8916 25280 8968
rect 24952 8848 25004 8900
rect 25596 8780 25648 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 2228 8576 2280 8628
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 4160 8576 4212 8628
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 8392 8576 8444 8628
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 3976 8508 4028 8560
rect 9036 8508 9088 8560
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 8760 8440 8812 8492
rect 10048 8440 10100 8492
rect 4804 8372 4856 8424
rect 15108 8576 15160 8628
rect 16764 8576 16816 8628
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 20996 8576 21048 8628
rect 12072 8508 12124 8560
rect 13268 8440 13320 8492
rect 14280 8440 14332 8492
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 10508 8372 10560 8424
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 12624 8372 12676 8424
rect 16672 8440 16724 8492
rect 16304 8415 16356 8424
rect 16304 8381 16313 8415
rect 16313 8381 16347 8415
rect 16347 8381 16356 8415
rect 16304 8372 16356 8381
rect 3792 8304 3844 8356
rect 14832 8304 14884 8356
rect 11152 8236 11204 8288
rect 13820 8236 13872 8288
rect 15844 8236 15896 8288
rect 19616 8508 19668 8560
rect 19800 8508 19852 8560
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 18788 8440 18840 8492
rect 20076 8440 20128 8492
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 17316 8372 17368 8424
rect 17592 8372 17644 8424
rect 18880 8372 18932 8424
rect 19340 8372 19392 8424
rect 22008 8372 22060 8424
rect 23388 8372 23440 8424
rect 24216 8304 24268 8356
rect 16856 8236 16908 8288
rect 19064 8236 19116 8288
rect 19432 8236 19484 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 1952 8032 2004 8084
rect 2780 8032 2832 8084
rect 3608 8075 3660 8084
rect 3608 8041 3617 8075
rect 3617 8041 3651 8075
rect 3651 8041 3660 8075
rect 3608 8032 3660 8041
rect 10324 8032 10376 8084
rect 12164 8032 12216 8084
rect 12532 8032 12584 8084
rect 13912 8032 13964 8084
rect 14280 8032 14332 8084
rect 2596 8007 2648 8016
rect 2596 7973 2605 8007
rect 2605 7973 2639 8007
rect 2639 7973 2648 8007
rect 2596 7964 2648 7973
rect 3884 7964 3936 8016
rect 16856 8032 16908 8084
rect 16948 8032 17000 8084
rect 17960 8032 18012 8084
rect 18880 8032 18932 8084
rect 19156 8032 19208 8084
rect 20076 8075 20128 8084
rect 20076 8041 20085 8075
rect 20085 8041 20119 8075
rect 20119 8041 20128 8075
rect 20076 8032 20128 8041
rect 15108 8007 15160 8016
rect 15108 7973 15117 8007
rect 15117 7973 15151 8007
rect 15151 7973 15160 8007
rect 15108 7964 15160 7973
rect 22192 7964 22244 8016
rect 20720 7896 20772 7948
rect 2596 7828 2648 7880
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 14004 7828 14056 7880
rect 15200 7828 15252 7880
rect 16396 7828 16448 7880
rect 6552 7760 6604 7812
rect 11612 7760 11664 7812
rect 13820 7760 13872 7812
rect 17408 7828 17460 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 20444 7828 20496 7880
rect 16764 7760 16816 7812
rect 23664 7896 23716 7948
rect 22376 7828 22428 7880
rect 22836 7871 22888 7880
rect 22836 7837 22845 7871
rect 22845 7837 22879 7871
rect 22879 7837 22888 7871
rect 22836 7828 22888 7837
rect 26240 7896 26292 7948
rect 24400 7828 24452 7880
rect 1676 7692 1728 7744
rect 11336 7692 11388 7744
rect 13728 7692 13780 7744
rect 16212 7735 16264 7744
rect 16212 7701 16221 7735
rect 16221 7701 16255 7735
rect 16255 7701 16264 7735
rect 16212 7692 16264 7701
rect 16672 7692 16724 7744
rect 24952 7760 25004 7812
rect 22192 7735 22244 7744
rect 22192 7701 22201 7735
rect 22201 7701 22235 7735
rect 22235 7701 22244 7735
rect 22192 7692 22244 7701
rect 25228 7735 25280 7744
rect 25228 7701 25237 7735
rect 25237 7701 25271 7735
rect 25271 7701 25280 7735
rect 25228 7692 25280 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 10508 7488 10560 7540
rect 12256 7488 12308 7540
rect 15016 7531 15068 7540
rect 15016 7497 15025 7531
rect 15025 7497 15059 7531
rect 15059 7497 15068 7531
rect 15016 7488 15068 7497
rect 15200 7488 15252 7540
rect 15936 7488 15988 7540
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 17408 7488 17460 7540
rect 18512 7488 18564 7540
rect 23848 7488 23900 7540
rect 6184 7420 6236 7472
rect 6736 7352 6788 7404
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 12900 7420 12952 7472
rect 12532 7284 12584 7336
rect 12900 7284 12952 7336
rect 13820 7284 13872 7336
rect 14648 7352 14700 7404
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 16580 7420 16632 7472
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 25872 7420 25924 7472
rect 20444 7352 20496 7404
rect 16764 7284 16816 7336
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 4528 7216 4580 7268
rect 16212 7216 16264 7268
rect 18052 7284 18104 7336
rect 23940 7395 23992 7404
rect 23940 7361 23949 7395
rect 23949 7361 23983 7395
rect 23983 7361 23992 7395
rect 23940 7352 23992 7361
rect 24676 7352 24728 7404
rect 23296 7327 23348 7336
rect 23296 7293 23305 7327
rect 23305 7293 23339 7327
rect 23339 7293 23348 7327
rect 23296 7284 23348 7293
rect 22744 7216 22796 7268
rect 10324 7191 10376 7200
rect 10324 7157 10333 7191
rect 10333 7157 10367 7191
rect 10367 7157 10376 7191
rect 10324 7148 10376 7157
rect 12256 7148 12308 7200
rect 20720 7148 20772 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 12624 6944 12676 6996
rect 14556 6944 14608 6996
rect 18052 6944 18104 6996
rect 18144 6944 18196 6996
rect 15200 6876 15252 6928
rect 26792 6944 26844 6996
rect 19248 6919 19300 6928
rect 19248 6885 19257 6919
rect 19257 6885 19291 6919
rect 19291 6885 19300 6919
rect 19248 6876 19300 6885
rect 22008 6876 22060 6928
rect 5356 6808 5408 6860
rect 10140 6808 10192 6860
rect 1400 6740 1452 6792
rect 11520 6740 11572 6792
rect 3424 6672 3476 6724
rect 8300 6672 8352 6724
rect 9588 6672 9640 6724
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 13268 6740 13320 6792
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 11152 6604 11204 6613
rect 13452 6672 13504 6724
rect 15108 6740 15160 6792
rect 15936 6740 15988 6792
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 16580 6783 16632 6792
rect 16580 6749 16589 6783
rect 16589 6749 16623 6783
rect 16623 6749 16632 6783
rect 16580 6740 16632 6749
rect 17500 6808 17552 6860
rect 19156 6808 19208 6860
rect 20352 6851 20404 6860
rect 20352 6817 20361 6851
rect 20361 6817 20395 6851
rect 20395 6817 20404 6851
rect 20352 6808 20404 6817
rect 17224 6740 17276 6792
rect 20720 6740 20772 6792
rect 22192 6808 22244 6860
rect 22560 6808 22612 6860
rect 22284 6740 22336 6792
rect 11888 6604 11940 6656
rect 14464 6647 14516 6656
rect 14464 6613 14473 6647
rect 14473 6613 14507 6647
rect 14507 6613 14516 6647
rect 14464 6604 14516 6613
rect 25228 6740 25280 6792
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 16028 6647 16080 6656
rect 16028 6613 16037 6647
rect 16037 6613 16071 6647
rect 16071 6613 16080 6647
rect 16028 6604 16080 6613
rect 16764 6604 16816 6656
rect 25688 6672 25740 6724
rect 19984 6604 20036 6656
rect 21548 6604 21600 6656
rect 25044 6604 25096 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 9864 6400 9916 6452
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 12900 6443 12952 6452
rect 12900 6409 12909 6443
rect 12909 6409 12943 6443
rect 12943 6409 12952 6443
rect 12900 6400 12952 6409
rect 14464 6400 14516 6452
rect 15108 6400 15160 6452
rect 15476 6443 15528 6452
rect 15476 6409 15485 6443
rect 15485 6409 15519 6443
rect 15519 6409 15528 6443
rect 15476 6400 15528 6409
rect 16120 6443 16172 6452
rect 16120 6409 16129 6443
rect 16129 6409 16163 6443
rect 16163 6409 16172 6443
rect 16120 6400 16172 6409
rect 7656 6332 7708 6384
rect 11888 6332 11940 6384
rect 12716 6332 12768 6384
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 13360 6264 13412 6316
rect 14188 6307 14240 6316
rect 14188 6273 14197 6307
rect 14197 6273 14231 6307
rect 14231 6273 14240 6307
rect 14188 6264 14240 6273
rect 15292 6264 15344 6316
rect 11980 6128 12032 6180
rect 14924 6196 14976 6248
rect 22008 6400 22060 6452
rect 22376 6400 22428 6452
rect 17040 6332 17092 6384
rect 18696 6332 18748 6384
rect 18880 6332 18932 6384
rect 23480 6332 23532 6384
rect 17224 6196 17276 6248
rect 17776 6264 17828 6316
rect 19616 6264 19668 6316
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 20812 6307 20864 6316
rect 20812 6273 20821 6307
rect 20821 6273 20855 6307
rect 20855 6273 20864 6307
rect 20812 6264 20864 6273
rect 24032 6332 24084 6384
rect 23940 6307 23992 6316
rect 23940 6273 23949 6307
rect 23949 6273 23983 6307
rect 23983 6273 23992 6307
rect 23940 6264 23992 6273
rect 19892 6196 19944 6248
rect 19984 6196 20036 6248
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 23940 6128 23992 6180
rect 9312 6060 9364 6112
rect 13268 6060 13320 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 15936 6060 15988 6112
rect 17592 6060 17644 6112
rect 18236 6060 18288 6112
rect 18604 6060 18656 6112
rect 19984 6060 20036 6112
rect 21640 6060 21692 6112
rect 22836 6060 22888 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 10600 5856 10652 5908
rect 16764 5856 16816 5908
rect 16948 5856 17000 5908
rect 18420 5856 18472 5908
rect 5632 5788 5684 5840
rect 21548 5788 21600 5840
rect 10232 5720 10284 5772
rect 21364 5763 21416 5772
rect 21364 5729 21373 5763
rect 21373 5729 21407 5763
rect 21407 5729 21416 5763
rect 21364 5720 21416 5729
rect 13728 5652 13780 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 17132 5652 17184 5704
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 17592 5627 17644 5636
rect 17592 5593 17601 5627
rect 17601 5593 17635 5627
rect 17635 5593 17644 5627
rect 17592 5584 17644 5593
rect 17776 5627 17828 5636
rect 17776 5593 17785 5627
rect 17785 5593 17819 5627
rect 17819 5593 17828 5627
rect 17776 5584 17828 5593
rect 13360 5516 13412 5568
rect 13728 5516 13780 5568
rect 15752 5516 15804 5568
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 18880 5627 18932 5636
rect 18880 5593 18889 5627
rect 18889 5593 18923 5627
rect 18923 5593 18932 5627
rect 18880 5584 18932 5593
rect 19156 5584 19208 5636
rect 18604 5516 18656 5568
rect 24952 5584 25004 5636
rect 25228 5559 25280 5568
rect 25228 5525 25237 5559
rect 25237 5525 25271 5559
rect 25271 5525 25280 5559
rect 25228 5516 25280 5525
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 13544 5355 13596 5364
rect 13544 5321 13553 5355
rect 13553 5321 13587 5355
rect 13587 5321 13596 5355
rect 13544 5312 13596 5321
rect 2412 5244 2464 5296
rect 12808 5176 12860 5228
rect 14096 5312 14148 5364
rect 14740 5312 14792 5364
rect 15568 5355 15620 5364
rect 15568 5321 15577 5355
rect 15577 5321 15611 5355
rect 15611 5321 15620 5355
rect 15568 5312 15620 5321
rect 17592 5312 17644 5364
rect 17960 5312 18012 5364
rect 18972 5312 19024 5364
rect 18512 5244 18564 5296
rect 20904 5312 20956 5364
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17592 5176 17644 5228
rect 17960 5176 18012 5228
rect 22836 5244 22888 5296
rect 19892 5176 19944 5228
rect 21088 5176 21140 5228
rect 25320 5312 25372 5364
rect 24860 5244 24912 5296
rect 23940 5219 23992 5228
rect 23940 5185 23949 5219
rect 23949 5185 23983 5219
rect 23983 5185 23992 5219
rect 23940 5176 23992 5185
rect 8484 5040 8536 5092
rect 12256 5040 12308 5092
rect 16396 5040 16448 5092
rect 16488 5083 16540 5092
rect 16488 5049 16497 5083
rect 16497 5049 16531 5083
rect 16531 5049 16540 5083
rect 16488 5040 16540 5049
rect 17500 5083 17552 5092
rect 17500 5049 17509 5083
rect 17509 5049 17543 5083
rect 17543 5049 17552 5083
rect 17500 5040 17552 5049
rect 17592 5040 17644 5092
rect 17868 5040 17920 5092
rect 18052 5108 18104 5160
rect 23388 5108 23440 5160
rect 24676 5151 24728 5160
rect 24676 5117 24685 5151
rect 24685 5117 24719 5151
rect 24719 5117 24728 5151
rect 24676 5108 24728 5117
rect 26056 5040 26108 5092
rect 14004 4972 14056 5024
rect 17132 4972 17184 5024
rect 19248 5015 19300 5024
rect 19248 4981 19257 5015
rect 19257 4981 19291 5015
rect 19291 4981 19300 5015
rect 19248 4972 19300 4981
rect 20444 4972 20496 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 8668 4768 8720 4820
rect 10784 4768 10836 4820
rect 16856 4768 16908 4820
rect 17132 4811 17184 4820
rect 17132 4777 17141 4811
rect 17141 4777 17175 4811
rect 17175 4777 17184 4811
rect 17132 4768 17184 4777
rect 19616 4768 19668 4820
rect 25412 4768 25464 4820
rect 16212 4700 16264 4752
rect 19248 4700 19300 4752
rect 17408 4632 17460 4684
rect 7840 4564 7892 4616
rect 15016 4607 15068 4616
rect 15016 4573 15025 4607
rect 15025 4573 15059 4607
rect 15059 4573 15068 4607
rect 15016 4564 15068 4573
rect 16304 4564 16356 4616
rect 16488 4564 16540 4616
rect 17132 4564 17184 4616
rect 26148 4700 26200 4752
rect 20444 4564 20496 4616
rect 23756 4632 23808 4684
rect 22468 4564 22520 4616
rect 25044 4564 25096 4616
rect 10048 4496 10100 4548
rect 18052 4496 18104 4548
rect 18696 4539 18748 4548
rect 18696 4505 18705 4539
rect 18705 4505 18739 4539
rect 18739 4505 18748 4539
rect 18696 4496 18748 4505
rect 14832 4428 14884 4480
rect 17868 4428 17920 4480
rect 17960 4471 18012 4480
rect 17960 4437 17969 4471
rect 17969 4437 18003 4471
rect 18003 4437 18012 4471
rect 17960 4428 18012 4437
rect 23388 4496 23440 4548
rect 24952 4496 25004 4548
rect 22652 4428 22704 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 16304 4267 16356 4276
rect 16304 4233 16313 4267
rect 16313 4233 16347 4267
rect 16347 4233 16356 4267
rect 16304 4224 16356 4233
rect 16396 4224 16448 4276
rect 26332 4224 26384 4276
rect 10324 4156 10376 4208
rect 18696 4156 18748 4208
rect 19156 4156 19208 4208
rect 26424 4156 26476 4208
rect 9128 4088 9180 4140
rect 10876 4088 10928 4140
rect 16948 4088 17000 4140
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 12440 4020 12492 4072
rect 13544 4020 13596 4072
rect 14280 4020 14332 4072
rect 18236 4088 18288 4140
rect 18604 4088 18656 4140
rect 19340 4088 19392 4140
rect 19984 4088 20036 4140
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 17500 4063 17552 4072
rect 17500 4029 17509 4063
rect 17509 4029 17543 4063
rect 17543 4029 17552 4063
rect 17500 4020 17552 4029
rect 17776 4020 17828 4072
rect 23480 4088 23532 4140
rect 22284 4020 22336 4072
rect 11704 3952 11756 4004
rect 16948 3952 17000 4004
rect 19156 3952 19208 4004
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 24952 3952 25004 4004
rect 7380 3884 7432 3936
rect 13544 3884 13596 3936
rect 18236 3884 18288 3936
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19432 3884 19484 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 7840 3680 7892 3732
rect 10692 3680 10744 3732
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 9404 3476 9456 3528
rect 18328 3680 18380 3732
rect 19708 3680 19760 3732
rect 20536 3680 20588 3732
rect 25596 3680 25648 3732
rect 17684 3612 17736 3664
rect 20076 3612 20128 3664
rect 19524 3544 19576 3596
rect 9772 3408 9824 3460
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 25136 3544 25188 3596
rect 21916 3476 21968 3528
rect 22652 3519 22704 3528
rect 22652 3485 22661 3519
rect 22661 3485 22695 3519
rect 22695 3485 22704 3519
rect 22652 3476 22704 3485
rect 25228 3476 25280 3528
rect 8484 3340 8536 3392
rect 19984 3408 20036 3460
rect 23388 3408 23440 3460
rect 25688 3408 25740 3460
rect 20444 3340 20496 3392
rect 24492 3340 24544 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 17592 3136 17644 3188
rect 20444 3136 20496 3188
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 22192 3068 22244 3120
rect 24860 3068 24912 3120
rect 21824 3000 21876 3052
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 26608 3000 26660 3052
rect 21180 2932 21232 2984
rect 6736 2864 6788 2916
rect 8668 2864 8720 2916
rect 10968 2864 11020 2916
rect 24584 2975 24636 2984
rect 24584 2941 24593 2975
rect 24593 2941 24627 2975
rect 24627 2941 24636 2975
rect 24584 2932 24636 2941
rect 25044 2864 25096 2916
rect 7196 2796 7248 2848
rect 20720 2796 20772 2848
rect 22560 2796 22612 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 7564 2592 7616 2644
rect 8668 2635 8720 2644
rect 8668 2601 8677 2635
rect 8677 2601 8711 2635
rect 8711 2601 8720 2635
rect 8668 2592 8720 2601
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 17408 2592 17460 2644
rect 7196 2524 7248 2576
rect 22100 2592 22152 2644
rect 25136 2592 25188 2644
rect 13636 2456 13688 2508
rect 19340 2456 19392 2508
rect 8668 2388 8720 2440
rect 19524 2388 19576 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 23480 2524 23532 2576
rect 24860 2456 24912 2508
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 19340 2252 19392 2304
rect 19432 2295 19484 2304
rect 19432 2261 19441 2295
rect 19441 2261 19475 2295
rect 19475 2261 19484 2295
rect 19432 2252 19484 2261
rect 20720 2320 20772 2372
rect 24952 2320 25004 2372
rect 20260 2252 20312 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 15016 2048 15068 2100
rect 22652 2048 22704 2100
rect 12532 1980 12584 2032
rect 19432 1980 19484 2032
rect 19524 1980 19576 2032
rect 24124 1980 24176 2032
rect 17316 1912 17368 1964
rect 24584 1912 24636 1964
rect 13728 1844 13780 1896
rect 19892 1844 19944 1896
rect 11612 1776 11664 1828
rect 20536 1776 20588 1828
<< metal2 >>
rect 1214 26888 1270 26897
rect 1214 26823 1270 26832
rect 1032 26376 1084 26382
rect 1032 26318 1084 26324
rect 938 25800 994 25809
rect 572 25764 624 25770
rect 938 25735 994 25744
rect 572 25706 624 25712
rect 478 25120 534 25129
rect 478 25055 534 25064
rect 492 15337 520 25055
rect 478 15328 534 15337
rect 478 15263 534 15272
rect 584 9382 612 25706
rect 952 25129 980 25735
rect 938 25120 994 25129
rect 938 25055 994 25064
rect 756 24948 808 24954
rect 756 24890 808 24896
rect 662 24304 718 24313
rect 662 24239 718 24248
rect 676 11830 704 24239
rect 664 11824 716 11830
rect 664 11766 716 11772
rect 572 9376 624 9382
rect 572 9318 624 9324
rect 768 9042 796 24890
rect 848 21616 900 21622
rect 848 21558 900 21564
rect 860 12306 888 21558
rect 938 21040 994 21049
rect 938 20975 994 20984
rect 848 12300 900 12306
rect 848 12242 900 12248
rect 952 10470 980 20975
rect 1044 10606 1072 26318
rect 1124 25016 1176 25022
rect 1124 24958 1176 24964
rect 1032 10600 1084 10606
rect 1032 10542 1084 10548
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 1136 9722 1164 24958
rect 1228 15473 1256 26823
rect 1674 26200 1730 27000
rect 2042 26200 2098 27000
rect 2410 26330 2466 27000
rect 2778 26330 2834 27000
rect 3146 26330 3202 27000
rect 2136 26308 2188 26314
rect 2136 26250 2188 26256
rect 2410 26302 2728 26330
rect 1584 26172 1636 26178
rect 1584 26114 1636 26120
rect 1596 24410 1624 26114
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1688 22692 1716 26200
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 1768 24064 1820 24070
rect 1766 24032 1768 24041
rect 1820 24032 1822 24041
rect 1766 23967 1822 23976
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1596 22664 1716 22692
rect 1308 21344 1360 21350
rect 1308 21286 1360 21292
rect 1214 15464 1270 15473
rect 1214 15399 1270 15408
rect 1320 14074 1348 21286
rect 1492 19440 1544 19446
rect 1492 19382 1544 19388
rect 1504 15586 1532 19382
rect 1596 19310 1624 22664
rect 1676 22432 1728 22438
rect 1676 22374 1728 22380
rect 1688 21554 1716 22374
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1780 19122 1808 23462
rect 1872 22234 1900 25842
rect 1950 23080 2006 23089
rect 1950 23015 2006 23024
rect 1860 22228 1912 22234
rect 1860 22170 1912 22176
rect 1872 22137 1900 22170
rect 1858 22128 1914 22137
rect 1858 22063 1914 22072
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1596 19094 1808 19122
rect 1596 16250 1624 19094
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1688 18426 1716 18702
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17678 1716 18022
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1688 16574 1716 17614
rect 1688 16546 1808 16574
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1504 15558 1624 15586
rect 1492 15428 1544 15434
rect 1492 15370 1544 15376
rect 1398 15328 1454 15337
rect 1398 15263 1454 15272
rect 1308 14068 1360 14074
rect 1308 14010 1360 14016
rect 1320 13326 1348 14010
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1124 9716 1176 9722
rect 1124 9658 1176 9664
rect 756 9036 808 9042
rect 756 8978 808 8984
rect 1412 6798 1440 15263
rect 1504 10266 1532 15370
rect 1596 14414 1624 15558
rect 1676 14884 1728 14890
rect 1676 14826 1728 14832
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 13938 1624 14214
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1582 9208 1638 9217
rect 1582 9143 1584 9152
rect 1636 9143 1638 9152
rect 1584 9114 1636 9120
rect 1596 8974 1624 9114
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1688 7750 1716 14826
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1780 6361 1808 16546
rect 1872 15094 1900 21966
rect 1964 19378 1992 23015
rect 2056 20806 2084 26200
rect 2148 21729 2176 26250
rect 2410 26200 2466 26302
rect 2412 25696 2464 25702
rect 2412 25638 2464 25644
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2226 23216 2282 23225
rect 2226 23151 2282 23160
rect 2240 23118 2268 23151
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2134 21720 2190 21729
rect 2134 21655 2190 21664
rect 2136 21548 2188 21554
rect 2136 21490 2188 21496
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2056 16574 2084 17478
rect 1964 16546 2084 16574
rect 1860 15088 1912 15094
rect 1860 15030 1912 15036
rect 1964 15042 1992 16546
rect 2148 15638 2176 21490
rect 2228 20936 2280 20942
rect 2226 20904 2228 20913
rect 2280 20904 2282 20913
rect 2226 20839 2282 20848
rect 2332 20330 2360 24142
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2424 18986 2452 25638
rect 2596 25628 2648 25634
rect 2596 25570 2648 25576
rect 2608 24041 2636 25570
rect 2594 24032 2650 24041
rect 2594 23967 2650 23976
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2516 22098 2544 22714
rect 2504 22092 2556 22098
rect 2504 22034 2556 22040
rect 2516 21457 2544 22034
rect 2502 21448 2558 21457
rect 2502 21383 2558 21392
rect 2504 20868 2556 20874
rect 2504 20810 2556 20816
rect 2516 19122 2544 20810
rect 2608 19310 2636 23666
rect 2700 23474 2728 26302
rect 2778 26302 2912 26330
rect 2778 26200 2834 26302
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2792 23769 2820 24550
rect 2778 23760 2834 23769
rect 2778 23695 2834 23704
rect 2700 23446 2820 23474
rect 2686 22536 2742 22545
rect 2686 22471 2742 22480
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2516 19094 2636 19122
rect 2424 18958 2544 18986
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 2240 15094 2268 18566
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2136 15088 2188 15094
rect 1964 15014 2084 15042
rect 2136 15030 2188 15036
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1872 13938 1900 14758
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1858 11656 1914 11665
rect 1858 11591 1860 11600
rect 1912 11591 1914 11600
rect 1860 11562 1912 11568
rect 1858 11384 1914 11393
rect 1858 11319 1860 11328
rect 1912 11319 1914 11328
rect 1860 11290 1912 11296
rect 1872 11150 1900 11290
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1964 8090 1992 14894
rect 2056 12986 2084 15014
rect 2148 14906 2176 15030
rect 2148 14878 2268 14906
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2056 11257 2084 11698
rect 2042 11248 2098 11257
rect 2042 11183 2098 11192
rect 2148 9450 2176 13330
rect 2240 12374 2268 14878
rect 2332 14482 2360 16390
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2332 13410 2360 14282
rect 2424 13530 2452 16390
rect 2516 13530 2544 18958
rect 2608 15638 2636 19094
rect 2700 17338 2728 22471
rect 2792 21010 2820 23446
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 2792 19922 2820 20742
rect 2884 20380 2912 26302
rect 3146 26302 3372 26330
rect 3146 26200 3202 26302
rect 3238 25936 3294 25945
rect 3238 25871 3294 25880
rect 3252 25226 3280 25871
rect 3240 25220 3292 25226
rect 3240 25162 3292 25168
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2962 23760 3018 23769
rect 2962 23695 2964 23704
rect 3016 23695 3018 23704
rect 2964 23666 3016 23672
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3148 23248 3200 23254
rect 3148 23190 3200 23196
rect 3160 22710 3188 23190
rect 3148 22704 3200 22710
rect 3148 22646 3200 22652
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3344 22098 3372 26302
rect 3514 26200 3570 27000
rect 3882 26330 3938 27000
rect 3882 26302 4108 26330
rect 3882 26200 3938 26302
rect 3424 25832 3476 25838
rect 3424 25774 3476 25780
rect 3436 22778 3464 25774
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3422 22672 3478 22681
rect 3422 22607 3478 22616
rect 3436 22438 3464 22607
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3528 21486 3556 26200
rect 3698 24848 3754 24857
rect 3698 24783 3754 24792
rect 3712 24682 3740 24783
rect 3700 24676 3752 24682
rect 3700 24618 3752 24624
rect 3712 23322 3740 24618
rect 3976 24336 4028 24342
rect 3974 24304 3976 24313
rect 4028 24304 4030 24313
rect 3974 24239 4030 24248
rect 3700 23316 3752 23322
rect 3700 23258 3752 23264
rect 3700 22976 3752 22982
rect 3700 22918 3752 22924
rect 3608 22636 3660 22642
rect 3608 22578 3660 22584
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 3332 21072 3384 21078
rect 3332 21014 3384 21020
rect 2964 20392 3016 20398
rect 2884 20352 2964 20380
rect 2964 20334 3016 20340
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 3344 19802 3372 21014
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 2792 19774 3372 19802
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2700 16182 2728 16526
rect 2688 16176 2740 16182
rect 2688 16118 2740 16124
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 15162 2636 15438
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2594 15056 2650 15065
rect 2594 14991 2650 15000
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2332 13382 2452 13410
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 2240 8634 2268 11630
rect 2332 10198 2360 13194
rect 2424 12050 2452 13382
rect 2608 12866 2636 14991
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2516 12838 2636 12866
rect 2516 12238 2544 12838
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2504 12232 2556 12238
rect 2608 12209 2636 12718
rect 2504 12174 2556 12180
rect 2594 12200 2650 12209
rect 2594 12135 2650 12144
rect 2424 12022 2636 12050
rect 2410 11112 2466 11121
rect 2410 11047 2412 11056
rect 2464 11047 2466 11056
rect 2504 11076 2556 11082
rect 2412 11018 2464 11024
rect 2504 11018 2556 11024
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 9489 2360 9522
rect 2318 9480 2374 9489
rect 2318 9415 2374 9424
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1766 6352 1822 6361
rect 1766 6287 1822 6296
rect 2424 5302 2452 10542
rect 2516 9178 2544 11018
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2608 8974 2636 12022
rect 2700 11914 2728 14350
rect 2792 13002 2820 19774
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3436 17746 3464 18566
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 3422 17640 3478 17649
rect 3422 17575 3424 17584
rect 3476 17575 3478 17584
rect 3424 17546 3476 17552
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2870 16688 2926 16697
rect 2870 16623 2926 16632
rect 2884 14074 2912 16623
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2884 13326 2912 14010
rect 3344 13802 3372 16050
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2976 13258 3004 13466
rect 3252 13297 3280 13466
rect 3238 13288 3294 13297
rect 2964 13252 3016 13258
rect 3238 13223 3294 13232
rect 2964 13194 3016 13200
rect 2792 12974 3372 13002
rect 2870 12880 2926 12889
rect 2870 12815 2926 12824
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2792 12442 2820 12718
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2700 11898 2820 11914
rect 2884 11898 2912 12815
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2700 11892 2832 11898
rect 2700 11886 2780 11892
rect 2780 11834 2832 11840
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2792 11354 2820 11698
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2778 10024 2834 10033
rect 2778 9959 2780 9968
rect 2832 9959 2834 9968
rect 2780 9930 2832 9936
rect 2884 9450 2912 11698
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3252 10742 3280 10950
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3344 9178 3372 12974
rect 3436 12730 3464 17138
rect 3528 16590 3556 20742
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3528 14346 3556 14758
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3620 12850 3648 22578
rect 3712 22273 3740 22918
rect 3698 22264 3754 22273
rect 3698 22199 3754 22208
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3712 13870 3740 20266
rect 3804 17762 3832 22034
rect 4080 21978 4108 26302
rect 4250 26200 4306 27000
rect 4618 26200 4674 27000
rect 4894 26616 4950 26625
rect 4894 26551 4950 26560
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4172 24206 4200 25230
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4264 23202 4292 26200
rect 4528 25492 4580 25498
rect 4528 25434 4580 25440
rect 4436 24200 4488 24206
rect 4436 24142 4488 24148
rect 4172 23174 4292 23202
rect 4172 22710 4200 23174
rect 4252 23112 4304 23118
rect 4252 23054 4304 23060
rect 4160 22704 4212 22710
rect 4160 22646 4212 22652
rect 3976 21956 4028 21962
rect 4080 21950 4200 21978
rect 3976 21898 4028 21904
rect 3882 21720 3938 21729
rect 3882 21655 3938 21664
rect 3896 20058 3924 21655
rect 3988 21146 4016 21898
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 4172 21010 4200 21950
rect 4264 21690 4292 23054
rect 4342 21992 4398 22001
rect 4342 21927 4398 21936
rect 4252 21684 4304 21690
rect 4252 21626 4304 21632
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4068 20936 4120 20942
rect 4120 20884 4200 20890
rect 4068 20878 4200 20884
rect 4080 20862 4200 20878
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3988 19938 4016 20266
rect 4172 19990 4200 20862
rect 4356 20380 4384 21927
rect 4448 20602 4476 24142
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4356 20352 4476 20380
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 3896 19910 4016 19938
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 3896 18290 3924 19910
rect 3976 19780 4028 19786
rect 3976 19722 4028 19728
rect 3988 18766 4016 19722
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4080 19417 4108 19450
rect 4066 19408 4122 19417
rect 4066 19343 4122 19352
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4172 19242 4200 19314
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4066 19000 4122 19009
rect 4066 18935 4122 18944
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3976 17808 4028 17814
rect 3974 17776 3976 17785
rect 4028 17776 4030 17785
rect 3804 17734 3924 17762
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 3804 17338 3832 17614
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3896 15994 3924 17734
rect 3974 17711 4030 17720
rect 4080 16658 4108 18935
rect 4158 18864 4214 18873
rect 4158 18799 4214 18808
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 3804 15966 3924 15994
rect 3804 14958 3832 15966
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3974 15872 4030 15881
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3790 14784 3846 14793
rect 3790 14719 3846 14728
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3804 13682 3832 14719
rect 3712 13654 3832 13682
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3436 12702 3648 12730
rect 3514 12336 3570 12345
rect 3514 12271 3570 12280
rect 3422 11248 3478 11257
rect 3422 11183 3478 11192
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2594 8664 2650 8673
rect 2594 8599 2596 8608
rect 2648 8599 2650 8608
rect 2596 8570 2648 8576
rect 2792 8090 2820 8910
rect 3238 8800 3294 8809
rect 3238 8735 3294 8744
rect 3252 8634 3280 8735
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2596 8016 2648 8022
rect 2594 7984 2596 7993
rect 2648 7984 2650 7993
rect 2594 7919 2650 7928
rect 2608 7886 2636 7919
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3436 6730 3464 11183
rect 3528 9450 3556 12271
rect 3620 9674 3648 12702
rect 3712 10810 3740 13654
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3804 11762 3832 13194
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3790 11520 3846 11529
rect 3790 11455 3846 11464
rect 3804 11354 3832 11455
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3804 11150 3832 11290
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3896 10470 3924 15846
rect 3974 15807 4030 15816
rect 3988 14618 4016 15807
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 4080 14414 4108 16458
rect 4172 15706 4200 18799
rect 4264 18290 4292 20198
rect 4344 19984 4396 19990
rect 4344 19926 4396 19932
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4264 16250 4292 17138
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4068 14408 4120 14414
rect 3974 14376 4030 14385
rect 4068 14350 4120 14356
rect 3974 14311 4030 14320
rect 3988 14278 4016 14311
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 4172 14006 4200 14962
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 10742 4016 13670
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4172 12238 4200 13466
rect 4264 13394 4292 15506
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4356 11694 4384 19926
rect 4448 16674 4476 20352
rect 4540 19854 4568 25434
rect 4632 23186 4660 26200
rect 4804 25356 4856 25362
rect 4804 25298 4856 25304
rect 4816 23730 4844 25298
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4802 23352 4858 23361
rect 4802 23287 4858 23296
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4632 22001 4660 22918
rect 4816 22642 4844 23287
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4710 22128 4766 22137
rect 4710 22063 4766 22072
rect 4618 21992 4674 22001
rect 4618 21927 4674 21936
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4632 21010 4660 21830
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4724 20874 4752 22063
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 4710 20632 4766 20641
rect 4710 20567 4712 20576
rect 4764 20567 4766 20576
rect 4712 20538 4764 20544
rect 4816 20482 4844 21626
rect 4724 20454 4844 20482
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4540 19718 4568 19790
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4540 16794 4568 19246
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4632 17882 4660 18702
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4448 16646 4568 16674
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4448 15366 4476 16526
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4434 15192 4490 15201
rect 4434 15127 4490 15136
rect 4448 14414 4476 15127
rect 4540 15026 4568 16646
rect 4618 16552 4674 16561
rect 4618 16487 4674 16496
rect 4632 15502 4660 16487
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4724 15434 4752 20454
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4710 14920 4766 14929
rect 4710 14855 4766 14864
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4448 13462 4476 14350
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4436 13456 4488 13462
rect 4436 13398 4488 13404
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4434 10976 4490 10985
rect 4434 10911 4490 10920
rect 4342 10840 4398 10849
rect 4342 10775 4398 10784
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 4250 10568 4306 10577
rect 4250 10503 4306 10512
rect 3884 10464 3936 10470
rect 3790 10432 3846 10441
rect 3884 10406 3936 10412
rect 3790 10367 3846 10376
rect 3620 9646 3740 9674
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9178 3648 9318
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3620 8090 3648 8978
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3712 7313 3740 9646
rect 3804 8362 3832 10367
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3896 8022 3924 8774
rect 3988 8566 4016 8774
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3698 7304 3754 7313
rect 3698 7239 3754 7248
rect 4080 6769 4108 9318
rect 4158 9072 4214 9081
rect 4264 9042 4292 10503
rect 4356 10062 4384 10775
rect 4448 10606 4476 10911
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4448 10198 4476 10542
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4158 9007 4214 9016
rect 4252 9036 4304 9042
rect 4172 8974 4200 9007
rect 4252 8978 4304 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4172 8634 4200 8910
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4158 8528 4214 8537
rect 4158 8463 4160 8472
rect 4212 8463 4214 8472
rect 4160 8434 4212 8440
rect 4540 7274 4568 13738
rect 4632 12986 4660 14350
rect 4724 14074 4752 14855
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4724 13530 4752 13738
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4816 13138 4844 18906
rect 4908 17218 4936 26551
rect 4986 26330 5042 27000
rect 5170 26480 5226 26489
rect 5170 26415 5226 26424
rect 4986 26302 5120 26330
rect 4986 26200 5042 26302
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 18737 5028 21830
rect 5092 21486 5120 26302
rect 5184 21729 5212 26415
rect 5354 26200 5410 27000
rect 5448 26240 5500 26246
rect 5264 25424 5316 25430
rect 5264 25366 5316 25372
rect 5170 21720 5226 21729
rect 5170 21655 5226 21664
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 5092 20262 5120 20402
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 4986 18728 5042 18737
rect 4986 18663 5042 18672
rect 4908 17190 5120 17218
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4908 15910 4936 16390
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4908 13938 4936 15302
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4724 13110 4844 13138
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12866 4752 13110
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4632 12838 4752 12866
rect 4632 12238 4660 12838
rect 4710 12744 4766 12753
rect 4710 12679 4766 12688
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4618 11520 4674 11529
rect 4618 11455 4674 11464
rect 4632 9654 4660 11455
rect 4724 9654 4752 12679
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4710 9208 4766 9217
rect 4710 9143 4766 9152
rect 4724 8838 4752 9143
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4816 8430 4844 12922
rect 4908 12918 4936 13874
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 5000 7857 5028 16390
rect 5092 9926 5120 17190
rect 5184 16522 5212 21490
rect 5276 19242 5304 25366
rect 5368 23662 5396 26200
rect 5722 26200 5778 27000
rect 6090 26200 6146 27000
rect 6458 26200 6514 27000
rect 6826 26200 6882 27000
rect 7194 26330 7250 27000
rect 7194 26302 7512 26330
rect 7194 26200 7250 26302
rect 5448 26182 5500 26188
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5460 23497 5488 26182
rect 5446 23488 5502 23497
rect 5446 23423 5502 23432
rect 5736 22710 5764 26200
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 5540 22500 5592 22506
rect 5540 22442 5592 22448
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5368 21690 5396 21830
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5368 19378 5396 19654
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5276 18358 5304 18566
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5368 17882 5396 18226
rect 5460 18034 5488 21966
rect 5552 20806 5580 22442
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5644 20398 5672 22170
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5736 21078 5764 21626
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5644 19514 5672 19858
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5736 18766 5764 19654
rect 5828 19281 5856 23462
rect 5920 21690 5948 24142
rect 6000 22772 6052 22778
rect 6000 22714 6052 22720
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5908 21480 5960 21486
rect 5908 21422 5960 21428
rect 5814 19272 5870 19281
rect 5814 19207 5870 19216
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5460 18006 5580 18034
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5354 17232 5410 17241
rect 5354 17167 5356 17176
rect 5408 17167 5410 17176
rect 5356 17138 5408 17144
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 5276 16250 5304 16526
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5172 16176 5224 16182
rect 5172 16118 5224 16124
rect 5184 14414 5212 16118
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5276 14550 5304 15302
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5184 12986 5212 13194
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5262 12472 5318 12481
rect 5262 12407 5318 12416
rect 5170 11792 5226 11801
rect 5170 11727 5226 11736
rect 5184 10606 5212 11727
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5276 9738 5304 12407
rect 5092 9710 5304 9738
rect 5092 9110 5120 9710
rect 5172 9648 5224 9654
rect 5170 9616 5172 9625
rect 5224 9616 5226 9625
rect 5170 9551 5226 9560
rect 5368 9466 5396 13874
rect 5460 13530 5488 14962
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5184 9438 5396 9466
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5184 7993 5212 9438
rect 5460 9382 5488 12174
rect 5552 11694 5580 18006
rect 5644 17066 5672 18634
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 5736 16182 5764 17614
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5644 13394 5672 15914
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5736 14618 5764 15438
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5828 14346 5856 18566
rect 5920 17542 5948 21422
rect 6012 20890 6040 22714
rect 6104 21962 6132 26200
rect 6276 24336 6328 24342
rect 6276 24278 6328 24284
rect 6184 22976 6236 22982
rect 6184 22918 6236 22924
rect 6092 21956 6144 21962
rect 6092 21898 6144 21904
rect 6092 21684 6144 21690
rect 6092 21626 6144 21632
rect 6104 21350 6132 21626
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 6012 20862 6132 20890
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 6012 20602 6040 20742
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6012 19514 6040 20402
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 6000 18692 6052 18698
rect 6000 18634 6052 18640
rect 6012 18426 6040 18634
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5920 15162 5948 17070
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 6012 15502 6040 16934
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5170 7984 5226 7993
rect 5170 7919 5226 7928
rect 4986 7848 5042 7857
rect 4986 7783 5042 7792
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 5368 6866 5396 9318
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 4066 6760 4122 6769
rect 3424 6724 3476 6730
rect 4066 6695 4122 6704
rect 3424 6666 3476 6672
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 5644 5846 5672 12106
rect 5736 9178 5764 13806
rect 6104 13734 6132 20862
rect 6196 18630 6224 22918
rect 6288 21486 6316 24278
rect 6472 24274 6500 26200
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6552 24404 6604 24410
rect 6552 24346 6604 24352
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6564 23118 6592 24346
rect 6644 24336 6696 24342
rect 6644 24278 6696 24284
rect 6656 23730 6684 24278
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6748 23633 6776 25094
rect 6840 24018 6868 26200
rect 7288 25560 7340 25566
rect 7288 25502 7340 25508
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 7012 24064 7064 24070
rect 6840 23990 6960 24018
rect 7012 24006 7064 24012
rect 6828 23724 6880 23730
rect 6828 23666 6880 23672
rect 6734 23624 6790 23633
rect 6734 23559 6790 23568
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6734 23488 6790 23497
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 6276 19440 6328 19446
rect 6276 19382 6328 19388
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6182 18456 6238 18465
rect 6182 18391 6184 18400
rect 6236 18391 6238 18400
rect 6184 18362 6236 18368
rect 6196 17678 6224 18362
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6288 16590 6316 19382
rect 6380 18766 6408 22510
rect 6656 22094 6684 23462
rect 6734 23423 6790 23432
rect 6748 22778 6776 23423
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6564 22066 6684 22094
rect 6458 21448 6514 21457
rect 6458 21383 6514 21392
rect 6472 21350 6500 21383
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6472 19122 6500 20878
rect 6564 20466 6592 22066
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6644 21344 6696 21350
rect 6642 21312 6644 21321
rect 6696 21312 6698 21321
rect 6642 21247 6698 21256
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6748 20380 6776 21898
rect 6840 21146 6868 23666
rect 6932 21486 6960 23990
rect 7024 22778 7052 24006
rect 7208 23594 7236 24142
rect 7300 23905 7328 25502
rect 7286 23896 7342 23905
rect 7286 23831 7342 23840
rect 7380 23860 7432 23866
rect 7380 23802 7432 23808
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 7288 23112 7340 23118
rect 7288 23054 7340 23060
rect 7300 22930 7328 23054
rect 7208 22902 7328 22930
rect 7012 22772 7064 22778
rect 7012 22714 7064 22720
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 7010 21176 7066 21185
rect 6828 21140 6880 21146
rect 7010 21111 7066 21120
rect 6828 21082 6880 21088
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 6840 20482 6868 20946
rect 7024 20913 7052 21111
rect 7010 20904 7066 20913
rect 7010 20839 7066 20848
rect 6840 20454 7052 20482
rect 6642 20360 6698 20369
rect 6748 20352 6868 20380
rect 6642 20295 6698 20304
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6564 19224 6592 20198
rect 6656 19378 6684 20295
rect 6840 19854 6868 20352
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6748 19514 6776 19790
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6564 19196 6776 19224
rect 6472 19094 6592 19122
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6380 18329 6408 18566
rect 6366 18320 6422 18329
rect 6366 18255 6422 18264
rect 6564 17490 6592 19094
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6380 17462 6592 17490
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 5814 13560 5870 13569
rect 5814 13495 5870 13504
rect 5828 12986 5856 13495
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5814 12608 5870 12617
rect 5814 12543 5870 12552
rect 5828 11218 5856 12543
rect 6012 12434 6040 13126
rect 6104 12646 6132 13398
rect 6196 12918 6224 16526
rect 6380 15994 6408 17462
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6472 16114 6500 17274
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6564 16153 6592 16186
rect 6550 16144 6606 16153
rect 6460 16108 6512 16114
rect 6550 16079 6606 16088
rect 6460 16050 6512 16056
rect 6380 15966 6500 15994
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6012 12406 6132 12434
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5920 11762 5948 12038
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 6012 9994 6040 12038
rect 6104 11642 6132 12406
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 11801 6224 12174
rect 6182 11792 6238 11801
rect 6182 11727 6238 11736
rect 6104 11614 6224 11642
rect 6090 10296 6146 10305
rect 6090 10231 6146 10240
rect 6104 10062 6132 10231
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 6196 7478 6224 11614
rect 6288 8974 6316 15098
rect 6366 14512 6422 14521
rect 6366 14447 6368 14456
rect 6420 14447 6422 14456
rect 6368 14418 6420 14424
rect 6472 13954 6500 15966
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6564 14074 6592 14282
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6472 13926 6592 13954
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6380 11506 6408 13806
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12170 6500 13262
rect 6564 13002 6592 13926
rect 6656 13190 6684 18702
rect 6748 18170 6776 19196
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6840 18426 6868 18702
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6932 18290 6960 19382
rect 7024 19242 7052 20454
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6748 18142 6868 18170
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6748 17270 6776 17750
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6748 16114 6776 16934
rect 6840 16114 6868 18142
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6932 17882 6960 18090
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7024 17202 7052 18566
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7116 16674 7144 22578
rect 7208 17218 7236 22902
rect 7392 22094 7420 23802
rect 7300 22066 7420 22094
rect 7300 22030 7328 22066
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 7300 21010 7328 21422
rect 7392 21146 7420 21966
rect 7484 21486 7512 26302
rect 7562 26200 7618 27000
rect 7930 26330 7986 27000
rect 7668 26302 7986 26330
rect 7576 23662 7604 26200
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7668 23186 7696 26302
rect 7930 26200 7986 26302
rect 8298 26200 8354 27000
rect 8666 26200 8722 27000
rect 9034 26330 9090 27000
rect 8772 26302 9090 26330
rect 7746 25800 7802 25809
rect 7746 25735 7802 25744
rect 7760 25401 7788 25735
rect 7746 25392 7802 25401
rect 7746 25327 7802 25336
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7760 22094 7788 24006
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7852 22098 7880 23666
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8208 22106 8260 22112
rect 7668 22066 7788 22094
rect 7840 22092 7892 22098
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7286 20904 7342 20913
rect 7286 20839 7342 20848
rect 7300 20534 7328 20839
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7378 19816 7434 19825
rect 7378 19751 7434 19760
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7300 17338 7328 19110
rect 7392 18222 7420 19751
rect 7484 19514 7512 19994
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7392 17882 7420 18022
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7484 17762 7512 19314
rect 7392 17734 7512 17762
rect 7392 17338 7420 17734
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7484 17270 7512 17478
rect 7472 17264 7524 17270
rect 7208 17190 7420 17218
rect 7472 17206 7524 17212
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7286 17096 7342 17105
rect 6932 16646 7144 16674
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6748 13530 6776 15914
rect 6932 15314 6960 16646
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6840 15286 6960 15314
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6564 12974 6776 13002
rect 6840 12986 6868 15286
rect 7024 13530 7052 15982
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7116 13326 7144 16458
rect 7208 15978 7236 17070
rect 7286 17031 7342 17040
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7208 13258 7236 15574
rect 7300 15162 7328 17031
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7300 13802 7328 14418
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7286 13424 7342 13433
rect 7286 13359 7342 13368
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6918 13016 6974 13025
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 6380 11478 6500 11506
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6380 9450 6408 11086
rect 6472 10606 6500 11478
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6472 10130 6500 10406
rect 6564 10266 6592 12582
rect 6748 11354 6776 12974
rect 6828 12980 6880 12986
rect 6918 12951 6974 12960
rect 6828 12922 6880 12928
rect 6826 12880 6882 12889
rect 6932 12850 6960 12951
rect 6826 12815 6828 12824
rect 6880 12815 6882 12824
rect 6920 12844 6972 12850
rect 6828 12786 6880 12792
rect 7024 12832 7052 13126
rect 7300 12832 7328 13359
rect 7024 12804 7144 12832
rect 6920 12786 6972 12792
rect 6826 12744 6882 12753
rect 7010 12744 7066 12753
rect 6882 12702 6960 12730
rect 6826 12679 6882 12688
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6840 9874 6868 12582
rect 6932 12481 6960 12702
rect 7010 12679 7066 12688
rect 6918 12472 6974 12481
rect 6918 12407 6974 12416
rect 7024 11286 7052 12679
rect 7012 11280 7064 11286
rect 6918 11248 6974 11257
rect 7012 11222 7064 11228
rect 7116 11218 7144 12804
rect 7208 12804 7328 12832
rect 6918 11183 6974 11192
rect 7104 11212 7156 11218
rect 6748 9846 6868 9874
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6564 7818 6592 8774
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6748 7410 6776 9846
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 8634 6868 8910
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 6932 5681 6960 11183
rect 7104 11154 7156 11160
rect 7102 10840 7158 10849
rect 7102 10775 7104 10784
rect 7156 10775 7158 10784
rect 7104 10746 7156 10752
rect 7208 9586 7236 12804
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7300 9178 7328 12650
rect 7392 9518 7420 17190
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 14464 7512 15846
rect 7576 15706 7604 21286
rect 7668 20641 7696 22066
rect 8312 22094 8340 26200
rect 8576 24880 8628 24886
rect 8576 24822 8628 24828
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8260 22066 8340 22094
rect 8208 22048 8260 22054
rect 7840 22034 7892 22040
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8390 21720 8446 21729
rect 8390 21655 8446 21664
rect 7748 20936 7800 20942
rect 7748 20878 7800 20884
rect 7654 20632 7710 20641
rect 7654 20567 7710 20576
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7668 19378 7696 19994
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7668 17338 7696 17614
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7654 16688 7710 16697
rect 7654 16623 7710 16632
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 14822 7604 15302
rect 7668 15162 7696 16623
rect 7760 15570 7788 20878
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 7838 20496 7894 20505
rect 7838 20431 7840 20440
rect 7892 20431 7894 20440
rect 7840 20402 7892 20408
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7852 19378 7880 20198
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7852 18290 7880 18566
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8220 17524 8248 17750
rect 8312 17746 8340 20334
rect 8404 20210 8432 21655
rect 8496 20602 8524 24346
rect 8588 21321 8616 24822
rect 8680 24138 8708 26200
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8666 22944 8722 22953
rect 8666 22879 8722 22888
rect 8574 21312 8630 21321
rect 8574 21247 8630 21256
rect 8574 21176 8630 21185
rect 8574 21111 8630 21120
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8404 20182 8524 20210
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8220 17496 8340 17524
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 17320 8340 17496
rect 8220 17292 8340 17320
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 7852 16232 7880 17002
rect 8128 16522 8156 17002
rect 8220 16522 8248 17292
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7932 16244 7984 16250
rect 7852 16204 7932 16232
rect 7932 16186 7984 16192
rect 8312 16114 8340 16390
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7838 15464 7894 15473
rect 7838 15399 7894 15408
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7484 14436 7696 14464
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7484 12170 7512 12718
rect 7562 12336 7618 12345
rect 7562 12271 7618 12280
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7576 12050 7604 12271
rect 7668 12238 7696 14436
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7484 12022 7604 12050
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7484 6225 7512 12022
rect 7760 11914 7788 14826
rect 7852 14278 7880 15399
rect 7944 15366 7972 15846
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8312 14414 8340 15302
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7840 13864 7892 13870
rect 8312 13841 8340 14010
rect 7840 13806 7892 13812
rect 8298 13832 8354 13841
rect 7852 12345 7880 13806
rect 8298 13767 8354 13776
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 7838 12336 7894 12345
rect 7838 12271 7894 12280
rect 7944 12186 7972 12854
rect 8404 12434 8432 19654
rect 8496 18306 8524 20182
rect 8588 19145 8616 21111
rect 8680 19922 8708 22879
rect 8772 22710 8800 26302
rect 9034 26200 9090 26302
rect 9402 26200 9458 27000
rect 9770 26330 9826 27000
rect 10138 26330 10194 27000
rect 9692 26302 9826 26330
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9232 23118 9260 23598
rect 9416 23338 9444 26200
rect 9496 25220 9548 25226
rect 9496 25162 9548 25168
rect 9508 23610 9536 25162
rect 9692 24274 9720 26302
rect 9770 26200 9826 26302
rect 9876 26302 10194 26330
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9588 23724 9640 23730
rect 9876 23712 9904 26302
rect 10138 26200 10194 26302
rect 10506 26330 10562 27000
rect 10506 26302 10824 26330
rect 10506 26200 10562 26302
rect 9640 23684 9904 23712
rect 9956 23724 10008 23730
rect 9588 23666 9640 23672
rect 9956 23666 10008 23672
rect 9508 23582 9628 23610
rect 9324 23310 9444 23338
rect 9324 23186 9352 23310
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 9034 22808 9090 22817
rect 9034 22743 9090 22752
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8944 22636 8996 22642
rect 8944 22578 8996 22584
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 8864 21894 8892 22034
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8956 21554 8984 22578
rect 9048 21894 9076 22743
rect 9218 22672 9274 22681
rect 9416 22642 9444 23122
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9218 22607 9274 22616
rect 9404 22636 9456 22642
rect 9232 22098 9260 22607
rect 9404 22578 9456 22584
rect 9404 22500 9456 22506
rect 9404 22442 9456 22448
rect 9416 22166 9444 22442
rect 9508 22409 9536 23054
rect 9494 22400 9550 22409
rect 9494 22335 9550 22344
rect 9404 22160 9456 22166
rect 9404 22102 9456 22108
rect 9220 22092 9272 22098
rect 9600 22094 9628 23582
rect 9680 23588 9732 23594
rect 9680 23530 9732 23536
rect 9692 23322 9720 23530
rect 9968 23497 9996 23666
rect 10796 23610 10824 26302
rect 10874 26200 10930 27000
rect 11242 26200 11298 27000
rect 11610 26200 11666 27000
rect 11978 26200 12034 27000
rect 12346 26200 12402 27000
rect 12714 26200 12770 27000
rect 13082 26200 13138 27000
rect 13450 26200 13506 27000
rect 13818 26200 13874 27000
rect 14186 26200 14242 27000
rect 14554 26330 14610 27000
rect 14292 26302 14610 26330
rect 10888 23730 10916 26200
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 10980 25401 11008 25910
rect 10966 25392 11022 25401
rect 10966 25327 11022 25336
rect 11256 24274 11284 26200
rect 11624 24954 11652 26200
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11886 24032 11942 24041
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10796 23582 11100 23610
rect 9954 23488 10010 23497
rect 9954 23423 10010 23432
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 10600 23044 10652 23050
rect 10600 22986 10652 22992
rect 9954 22808 10010 22817
rect 9220 22034 9272 22040
rect 9508 22066 9628 22094
rect 9692 22766 9954 22794
rect 9126 21992 9182 22001
rect 9126 21927 9182 21936
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 8772 20777 8800 20878
rect 8758 20768 8814 20777
rect 8758 20703 8814 20712
rect 8956 20466 8984 21490
rect 9048 21434 9076 21830
rect 9140 21593 9168 21927
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 9232 21690 9260 21830
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9126 21584 9182 21593
rect 9126 21519 9182 21528
rect 9048 21406 9168 21434
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 8864 20233 8892 20266
rect 8850 20224 8906 20233
rect 8850 20159 8906 20168
rect 8758 20088 8814 20097
rect 8758 20023 8814 20032
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8772 19242 8800 20023
rect 8956 19378 8984 20402
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8574 19136 8630 19145
rect 8574 19071 8630 19080
rect 8496 18278 8616 18306
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8496 17202 8524 18022
rect 8588 17921 8616 18278
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8574 17912 8630 17921
rect 8574 17847 8630 17856
rect 8680 17678 8708 18022
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8482 17096 8538 17105
rect 8482 17031 8538 17040
rect 8496 16833 8524 17031
rect 8482 16824 8538 16833
rect 8482 16759 8538 16768
rect 8588 16538 8616 17478
rect 8666 17368 8722 17377
rect 8666 17303 8722 17312
rect 8680 16658 8708 17303
rect 8772 16658 8800 19178
rect 8956 18290 8984 19314
rect 9034 18592 9090 18601
rect 9034 18527 9090 18536
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 17746 8984 18226
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8864 16810 8892 17682
rect 9048 17654 9076 18527
rect 9140 18193 9168 21406
rect 9218 21312 9274 21321
rect 9218 21247 9274 21256
rect 9232 19825 9260 21247
rect 9402 21176 9458 21185
rect 9402 21111 9458 21120
rect 9416 20058 9444 21111
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9218 19816 9274 19825
rect 9218 19751 9274 19760
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9402 19680 9458 19689
rect 9126 18184 9182 18193
rect 9126 18119 9182 18128
rect 9128 17808 9180 17814
rect 9232 17796 9260 19654
rect 9402 19615 9458 19624
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9324 18465 9352 18770
rect 9310 18456 9366 18465
rect 9310 18391 9366 18400
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9180 17768 9260 17796
rect 9128 17750 9180 17756
rect 9324 17728 9352 18022
rect 9416 17921 9444 19615
rect 9508 18970 9536 22066
rect 9692 21894 9720 22766
rect 9954 22743 10010 22752
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9600 21010 9628 21286
rect 9678 21040 9734 21049
rect 9588 21004 9640 21010
rect 9678 20975 9680 20984
rect 9588 20946 9640 20952
rect 9732 20975 9734 20984
rect 9680 20946 9732 20952
rect 9586 20632 9642 20641
rect 9586 20567 9642 20576
rect 9600 20369 9628 20567
rect 9680 20392 9732 20398
rect 9586 20360 9642 20369
rect 9680 20334 9732 20340
rect 9586 20295 9642 20304
rect 9692 19292 9720 20334
rect 9600 19264 9720 19292
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9402 17912 9458 17921
rect 9402 17847 9458 17856
rect 9508 17864 9536 18634
rect 9600 18601 9628 19264
rect 9586 18592 9642 18601
rect 9586 18527 9642 18536
rect 9678 17912 9734 17921
rect 9508 17836 9628 17864
rect 9678 17847 9734 17856
rect 9324 17700 9536 17728
rect 9036 17648 9088 17654
rect 9036 17590 9088 17596
rect 9220 17536 9272 17542
rect 9126 17504 9182 17513
rect 9220 17478 9272 17484
rect 9126 17439 9182 17448
rect 8864 16794 9076 16810
rect 8864 16788 9088 16794
rect 8864 16782 9036 16788
rect 9036 16730 9088 16736
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 9140 16674 9168 17439
rect 9232 17202 9260 17478
rect 9508 17252 9536 17700
rect 9600 17542 9628 17836
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9586 17368 9642 17377
rect 9692 17354 9720 17847
rect 9784 17377 9812 22510
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9876 17513 9904 21830
rect 10060 21078 10088 21966
rect 10612 21162 10640 22986
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10796 21978 10824 22918
rect 10796 21950 11008 21978
rect 11072 21962 11100 23582
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 10980 21706 11008 21950
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 11164 21894 11192 22578
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 10888 21678 11008 21706
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10428 21134 10640 21162
rect 10048 21072 10100 21078
rect 10048 21014 10100 21020
rect 9956 20800 10008 20806
rect 9954 20768 9956 20777
rect 10008 20768 10010 20777
rect 9954 20703 10010 20712
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9968 19718 9996 19994
rect 10428 19802 10456 21134
rect 10600 21004 10652 21010
rect 10704 20992 10732 21286
rect 10652 20964 10732 20992
rect 10600 20946 10652 20952
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10520 19825 10548 20198
rect 10244 19774 10456 19802
rect 10506 19816 10562 19825
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 10140 18760 10192 18766
rect 9954 18728 10010 18737
rect 10140 18702 10192 18708
rect 9954 18663 10010 18672
rect 9968 18329 9996 18663
rect 9954 18320 10010 18329
rect 9954 18255 10010 18264
rect 9862 17504 9918 17513
rect 9862 17439 9918 17448
rect 9642 17326 9720 17354
rect 9770 17368 9826 17377
rect 9586 17303 9642 17312
rect 9770 17303 9826 17312
rect 9416 17224 9536 17252
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9416 17116 9444 17224
rect 9496 17128 9548 17134
rect 9416 17088 9496 17116
rect 9496 17070 9548 17076
rect 9220 16992 9272 16998
rect 9272 16952 9536 16980
rect 9220 16934 9272 16940
rect 9508 16794 9536 16952
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9680 16720 9732 16726
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8484 16516 8536 16522
rect 8588 16510 8800 16538
rect 8484 16458 8536 16464
rect 7576 11886 7788 11914
rect 7852 12158 7972 12186
rect 8312 12406 8432 12434
rect 7576 9382 7604 11886
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7668 10810 7696 11766
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7760 11150 7788 11494
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7852 10690 7880 12158
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7668 10662 7880 10690
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7668 6390 7696 10662
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7760 9722 7788 9862
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7746 9616 7802 9625
rect 7746 9551 7748 9560
rect 7800 9551 7802 9560
rect 7748 9522 7800 9528
rect 7852 9178 7880 10474
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8312 9654 8340 12406
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8404 12102 8432 12310
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8390 11384 8446 11393
rect 8390 11319 8392 11328
rect 8444 11319 8446 11328
rect 8392 11290 8444 11296
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7852 8974 7880 9114
rect 7944 9042 7972 9114
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8404 8634 8432 9930
rect 8496 9042 8524 16458
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8588 15502 8616 16390
rect 8666 16280 8722 16289
rect 8666 16215 8668 16224
rect 8720 16215 8722 16224
rect 8668 16186 8720 16192
rect 8772 15978 8800 16510
rect 8864 16504 8892 16662
rect 9140 16646 9260 16674
rect 9680 16662 9732 16668
rect 9232 16522 9260 16646
rect 9692 16590 9720 16662
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9220 16516 9272 16522
rect 8864 16476 9168 16504
rect 9140 16402 9168 16476
rect 9220 16458 9272 16464
rect 9496 16448 9548 16454
rect 9402 16416 9458 16425
rect 9140 16374 9402 16402
rect 9496 16390 9548 16396
rect 9402 16351 9458 16360
rect 9508 16266 9536 16390
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 9416 16238 9536 16266
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8850 15736 8906 15745
rect 8850 15671 8906 15680
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8588 14618 8616 14962
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8574 13016 8630 13025
rect 8574 12951 8630 12960
rect 8588 12753 8616 12951
rect 8574 12744 8630 12753
rect 8574 12679 8630 12688
rect 8680 12696 8708 15370
rect 8680 12668 8800 12696
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8588 11830 8616 12038
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 11286 8616 11494
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8588 9489 8616 11086
rect 8772 11014 8800 12668
rect 8864 12186 8892 15671
rect 8956 14482 8984 16186
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9140 15473 9168 15506
rect 9126 15464 9182 15473
rect 9126 15399 9182 15408
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 9048 14657 9076 14894
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9034 14648 9090 14657
rect 9232 14618 9260 14826
rect 9034 14583 9036 14592
rect 9088 14583 9090 14592
rect 9220 14612 9272 14618
rect 9036 14554 9088 14560
rect 9220 14554 9272 14560
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 9232 14362 9260 14554
rect 9140 14334 9260 14362
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 13530 8984 14214
rect 9140 14006 9168 14334
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9232 13938 9260 14214
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9218 13560 9274 13569
rect 8944 13524 8996 13530
rect 9218 13495 9220 13504
rect 8944 13466 8996 13472
rect 9272 13495 9274 13504
rect 9220 13466 9272 13472
rect 8956 12850 8984 13466
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9140 12850 9168 13398
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9140 12238 9168 12786
rect 9232 12374 9260 13466
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 9128 12232 9180 12238
rect 8864 12158 8984 12186
rect 9128 12174 9180 12180
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11898 8892 12038
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11150 8892 11494
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8956 10792 8984 12158
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8864 10764 8984 10792
rect 8864 10538 8892 10764
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8956 9926 8984 10610
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8574 9480 8630 9489
rect 8574 9415 8630 9424
rect 8956 9178 8984 9862
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8680 8974 8708 9114
rect 8668 8968 8720 8974
rect 8482 8936 8538 8945
rect 8668 8910 8720 8916
rect 8482 8871 8538 8880
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7470 6216 7526 6225
rect 7470 6151 7526 6160
rect 6918 5672 6974 5681
rect 6918 5607 6974 5616
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 7392 3058 7420 3878
rect 7852 3738 7880 4558
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 6748 800 6776 2858
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7208 2582 7236 2790
rect 7576 2650 7604 3470
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8312 3097 8340 6666
rect 8496 5098 8524 8871
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8758 8528 8814 8537
rect 8758 8463 8760 8472
rect 8812 8463 8814 8472
rect 8760 8434 8812 8440
rect 8864 6905 8892 8774
rect 9048 8566 9076 11494
rect 9232 10826 9260 11698
rect 9324 11082 9352 13670
rect 9416 12306 9444 16238
rect 10152 16114 10180 18702
rect 10244 16697 10272 19774
rect 10506 19751 10562 19760
rect 10324 19712 10376 19718
rect 10416 19712 10468 19718
rect 10324 19654 10376 19660
rect 10414 19680 10416 19689
rect 10468 19680 10470 19689
rect 10336 19553 10364 19654
rect 10414 19615 10470 19624
rect 10322 19544 10378 19553
rect 10520 19530 10548 19751
rect 10322 19479 10378 19488
rect 10428 19502 10548 19530
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10336 18290 10364 19314
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10336 17610 10364 18226
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10230 16688 10286 16697
rect 10230 16623 10286 16632
rect 10428 16130 10456 19502
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10520 17542 10548 18226
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17270 10548 17478
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10612 16998 10640 20946
rect 10888 20346 10916 21678
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10980 20466 11008 21422
rect 11072 20534 11100 21490
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10888 20318 11008 20346
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10704 19514 10732 19790
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10782 17504 10838 17513
rect 10782 17439 10838 17448
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 9680 16108 9732 16114
rect 9600 16068 9680 16096
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9508 15473 9536 15982
rect 9494 15464 9550 15473
rect 9494 15399 9550 15408
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9508 13433 9536 14894
rect 9494 13424 9550 13433
rect 9494 13359 9550 13368
rect 9600 13326 9628 16068
rect 9680 16050 9732 16056
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10244 16102 10456 16130
rect 10520 16114 10548 16390
rect 10612 16250 10640 16390
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10508 16108 10560 16114
rect 9956 15904 10008 15910
rect 9954 15872 9956 15881
rect 10008 15872 10010 15881
rect 9954 15807 10010 15816
rect 9680 15632 9732 15638
rect 9680 15574 9732 15580
rect 9692 15473 9720 15574
rect 9678 15464 9734 15473
rect 9678 15399 9734 15408
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 10138 15056 10194 15065
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14550 9720 14758
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9968 13394 9996 15030
rect 10138 14991 10194 15000
rect 10152 13530 10180 14991
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10138 13424 10194 13433
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10048 13388 10100 13394
rect 10138 13359 10194 13368
rect 10048 13330 10100 13336
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9232 10798 9352 10826
rect 9218 10704 9274 10713
rect 9218 10639 9220 10648
rect 9272 10639 9274 10648
rect 9220 10610 9272 10616
rect 9232 10266 9260 10610
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8850 6896 8906 6905
rect 8850 6831 8906 6840
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8680 4826 8708 6258
rect 9324 6118 9352 10798
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8298 3088 8354 3097
rect 8496 3058 8524 3334
rect 9140 3194 9168 4082
rect 9416 3534 9444 9998
rect 9508 9110 9536 13126
rect 10060 12782 10088 13330
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9600 11558 9628 12242
rect 9678 11928 9734 11937
rect 9678 11863 9734 11872
rect 9692 11694 9720 11863
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9600 6730 9628 11222
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 8634 9720 11154
rect 9876 10674 9904 11290
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10060 9042 10088 12718
rect 10152 11898 10180 13359
rect 10244 12850 10272 16102
rect 10508 16050 10560 16056
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15706 10456 15846
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 15026 10548 15302
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10612 14482 10640 15506
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10612 14074 10640 14418
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10336 12442 10364 13806
rect 10428 13705 10456 13942
rect 10414 13696 10470 13705
rect 10414 13631 10470 13640
rect 10612 13530 10640 14010
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10612 13394 10640 13466
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10598 13152 10654 13161
rect 10598 13087 10654 13096
rect 10612 12889 10640 13087
rect 10598 12880 10654 12889
rect 10508 12844 10560 12850
rect 10598 12815 10654 12824
rect 10508 12786 10560 12792
rect 10520 12442 10548 12786
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9876 6458 9904 7822
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 10060 4554 10088 8434
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 8298 3023 8354 3032
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8680 2650 8708 2858
rect 9784 2650 9812 3402
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 8680 2446 8708 2586
rect 8668 2440 8720 2446
rect 10152 2417 10180 6802
rect 10244 5778 10272 12174
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10612 11082 10640 11154
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10598 10704 10654 10713
rect 10598 10639 10600 10648
rect 10652 10639 10654 10648
rect 10600 10610 10652 10616
rect 10704 10198 10732 17002
rect 10796 15337 10824 17439
rect 10888 17218 10916 19858
rect 10980 18834 11008 20318
rect 11164 20233 11192 20742
rect 11256 20534 11284 24006
rect 11716 23633 11744 24006
rect 11886 23967 11942 23976
rect 11900 23633 11928 23967
rect 11992 23662 12020 26200
rect 12360 24290 12388 26200
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12532 24676 12584 24682
rect 12532 24618 12584 24624
rect 12544 24313 12572 24618
rect 12530 24304 12586 24313
rect 12360 24274 12480 24290
rect 12360 24268 12492 24274
rect 12360 24262 12440 24268
rect 12530 24239 12586 24248
rect 12440 24210 12492 24216
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12360 24052 12388 24142
rect 12360 24041 12480 24052
rect 12360 24032 12494 24041
rect 12360 24024 12438 24032
rect 12438 23967 12494 23976
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12164 23792 12216 23798
rect 12164 23734 12216 23740
rect 11980 23656 12032 23662
rect 11702 23624 11758 23633
rect 11702 23559 11758 23568
rect 11886 23624 11942 23633
rect 11980 23598 12032 23604
rect 11886 23559 11942 23568
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11624 22982 11652 23462
rect 11716 23304 11744 23462
rect 11888 23316 11940 23322
rect 11716 23276 11888 23304
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11624 22710 11652 22918
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11716 22574 11744 23276
rect 11888 23258 11940 23264
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11348 21622 11376 22374
rect 11336 21616 11388 21622
rect 11336 21558 11388 21564
rect 11426 21584 11482 21593
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11348 20369 11376 21558
rect 11426 21519 11482 21528
rect 11334 20360 11390 20369
rect 11334 20295 11390 20304
rect 11244 20256 11296 20262
rect 11150 20224 11206 20233
rect 11244 20198 11296 20204
rect 11150 20159 11206 20168
rect 11256 19961 11284 20198
rect 11242 19952 11298 19961
rect 11242 19887 11298 19896
rect 11058 19408 11114 19417
rect 11058 19343 11114 19352
rect 11072 19310 11100 19343
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10888 17190 11008 17218
rect 10980 16998 11008 17190
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10874 16824 10930 16833
rect 10874 16759 10930 16768
rect 10782 15328 10838 15337
rect 10782 15263 10838 15272
rect 10888 15094 10916 16759
rect 10980 16182 11008 16934
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10692 10192 10744 10198
rect 10598 10160 10654 10169
rect 10692 10134 10744 10140
rect 10598 10095 10654 10104
rect 10612 10062 10640 10095
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10336 8090 10364 8842
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10428 7449 10456 9998
rect 10598 9616 10654 9625
rect 10796 9602 10824 13738
rect 10888 11762 10916 14758
rect 10966 14512 11022 14521
rect 10966 14447 10968 14456
rect 11020 14447 11022 14456
rect 10968 14418 11020 14424
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10980 12238 11008 14010
rect 11072 13190 11100 18158
rect 11164 16969 11192 18226
rect 11256 17882 11284 19887
rect 11440 19281 11468 21519
rect 11612 21480 11664 21486
rect 11612 21422 11664 21428
rect 11624 21350 11652 21422
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11532 19854 11560 20946
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11532 19514 11560 19790
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11426 19272 11482 19281
rect 11426 19207 11482 19216
rect 11518 18728 11574 18737
rect 11518 18663 11574 18672
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11426 18592 11482 18601
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11256 17066 11284 17478
rect 11348 17338 11376 18566
rect 11426 18527 11482 18536
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11150 16960 11206 16969
rect 11150 16895 11206 16904
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11164 16289 11192 16390
rect 11150 16280 11206 16289
rect 11150 16215 11206 16224
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11164 15094 11192 15982
rect 11242 15328 11298 15337
rect 11242 15263 11298 15272
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11256 14958 11284 15263
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11348 14464 11376 16594
rect 11256 14436 11376 14464
rect 11256 14074 11284 14436
rect 11334 14240 11390 14249
rect 11334 14175 11390 14184
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11242 13968 11298 13977
rect 11152 13932 11204 13938
rect 11242 13903 11298 13912
rect 11152 13874 11204 13880
rect 11164 13734 11192 13874
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11164 12986 11192 13194
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10966 12064 11022 12073
rect 10966 11999 11022 12008
rect 10980 11898 11008 11999
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10598 9551 10600 9560
rect 10652 9551 10654 9560
rect 10704 9574 10824 9602
rect 10600 9522 10652 9528
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10520 7546 10548 8366
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10414 7440 10470 7449
rect 10414 7375 10470 7384
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10336 4214 10364 7142
rect 10612 5914 10640 8366
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10704 3738 10732 9574
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10796 4826 10824 9454
rect 10888 8537 10916 11086
rect 10874 8528 10930 8537
rect 10874 8463 10930 8472
rect 10980 8412 11008 11086
rect 11072 10742 11100 12854
rect 11256 12102 11284 13903
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11242 11928 11298 11937
rect 11242 11863 11244 11872
rect 11296 11863 11298 11872
rect 11244 11834 11296 11840
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10742 11192 10950
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11348 10470 11376 14175
rect 11440 13954 11468 18527
rect 11532 18086 11560 18663
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11532 14521 11560 18022
rect 11518 14512 11574 14521
rect 11518 14447 11574 14456
rect 11440 13926 11560 13954
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11440 12714 11468 13806
rect 11532 13802 11560 13926
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11532 12850 11560 13466
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11532 12594 11560 12650
rect 11440 12566 11560 12594
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 10888 8384 11008 8412
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10888 4146 10916 8384
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10980 2922 11008 7822
rect 11164 7410 11192 8230
rect 11348 7750 11376 9862
rect 11440 8974 11468 12566
rect 11518 12472 11574 12481
rect 11518 12407 11574 12416
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11532 7698 11560 12407
rect 11624 12306 11652 21286
rect 11716 21185 11744 21286
rect 11702 21176 11758 21185
rect 11702 21111 11758 21120
rect 11704 20256 11756 20262
rect 11702 20224 11704 20233
rect 11756 20224 11758 20233
rect 11702 20159 11758 20168
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 17746 11744 18566
rect 11808 18222 11836 22714
rect 12176 22642 12204 23734
rect 12256 23044 12308 23050
rect 12256 22986 12308 22992
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12072 22568 12124 22574
rect 12268 22522 12296 22986
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12072 22510 12124 22516
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11992 20924 12020 21490
rect 12084 21486 12112 22510
rect 12176 22494 12296 22522
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 12084 21049 12112 21286
rect 12070 21040 12126 21049
rect 12070 20975 12126 20984
rect 12176 20924 12204 22494
rect 12360 22166 12388 22918
rect 12452 22574 12480 23802
rect 12636 23497 12664 25162
rect 12622 23488 12678 23497
rect 12622 23423 12678 23432
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12544 22710 12572 23258
rect 12636 22982 12664 23258
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12440 22568 12492 22574
rect 12636 22556 12664 22918
rect 12728 22642 12756 26200
rect 13096 25022 13124 26200
rect 13464 25537 13492 26200
rect 13728 25900 13780 25906
rect 13728 25842 13780 25848
rect 13450 25528 13506 25537
rect 13450 25463 13506 25472
rect 13084 25016 13136 25022
rect 13084 24958 13136 24964
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13360 23792 13412 23798
rect 13360 23734 13412 23740
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12992 23248 13044 23254
rect 12992 23190 13044 23196
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12440 22510 12492 22516
rect 12544 22528 12664 22556
rect 12348 22160 12400 22166
rect 12268 22120 12348 22148
rect 12268 21622 12296 22120
rect 12348 22102 12400 22108
rect 12440 22024 12492 22030
rect 12360 21984 12440 22012
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 11992 20896 12204 20924
rect 12176 20641 12204 20896
rect 12162 20632 12218 20641
rect 12162 20567 12218 20576
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11900 19281 11928 19314
rect 11886 19272 11942 19281
rect 11886 19207 11942 19216
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17134 11744 17682
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16114 11744 16526
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11716 15638 11744 16050
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11702 15328 11758 15337
rect 11702 15263 11758 15272
rect 11716 14113 11744 15263
rect 11702 14104 11758 14113
rect 11702 14039 11758 14048
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11716 12617 11744 12922
rect 11702 12608 11758 12617
rect 11702 12543 11758 12552
rect 11808 12434 11836 18022
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11900 16697 11928 17138
rect 11886 16688 11942 16697
rect 11886 16623 11942 16632
rect 11888 16516 11940 16522
rect 11992 16504 12020 20266
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 12162 20224 12218 20233
rect 12084 19417 12112 20198
rect 12162 20159 12218 20168
rect 12070 19408 12126 19417
rect 12070 19343 12126 19352
rect 12176 19292 12204 20159
rect 12360 19334 12388 21984
rect 12440 21966 12492 21972
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12452 20097 12480 21830
rect 12438 20088 12494 20097
rect 12438 20023 12494 20032
rect 12084 19264 12204 19292
rect 12256 19304 12308 19310
rect 12360 19306 12480 19334
rect 12084 18902 12112 19264
rect 12256 19246 12308 19252
rect 12268 18902 12296 19246
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12084 17882 12112 18838
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12268 18358 12296 18702
rect 12360 18630 12388 18906
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12348 18216 12400 18222
rect 12176 18176 12348 18204
rect 12176 17921 12204 18176
rect 12348 18158 12400 18164
rect 12256 18080 12308 18086
rect 12452 18057 12480 19306
rect 12256 18022 12308 18028
rect 12438 18048 12494 18057
rect 12162 17912 12218 17921
rect 12072 17876 12124 17882
rect 12162 17847 12218 17856
rect 12072 17818 12124 17824
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12084 17610 12112 17682
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 12072 17060 12124 17066
rect 12072 17002 12124 17008
rect 11940 16476 12020 16504
rect 11888 16458 11940 16464
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11900 15434 11928 16118
rect 11992 15434 12020 16476
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11900 14414 11928 15370
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11886 14104 11942 14113
rect 11886 14039 11942 14048
rect 11716 12406 11836 12434
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11898 11652 12038
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11624 9450 11652 10202
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11624 7818 11652 8842
rect 11716 8838 11744 12406
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11762 11836 12174
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 9722 11836 10610
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11808 9178 11836 9522
rect 11900 9450 11928 14039
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11992 11354 12020 12174
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12084 11234 12112 17002
rect 12176 16454 12204 17847
rect 12268 16640 12296 18022
rect 12438 17983 12494 17992
rect 12360 17882 12480 17898
rect 12348 17876 12492 17882
rect 12400 17870 12440 17876
rect 12348 17818 12400 17824
rect 12440 17818 12492 17824
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12452 17066 12480 17682
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12544 16833 12572 22528
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12636 21962 12664 22034
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12636 21010 12664 21422
rect 12728 21078 12756 21422
rect 12716 21072 12768 21078
rect 12716 21014 12768 21020
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12716 20868 12768 20874
rect 12716 20810 12768 20816
rect 12728 20641 12756 20810
rect 12714 20632 12770 20641
rect 12714 20567 12770 20576
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12714 20360 12770 20369
rect 12636 20233 12664 20334
rect 12714 20295 12770 20304
rect 12622 20224 12678 20233
rect 12622 20159 12678 20168
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12636 18222 12664 18770
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12530 16824 12586 16833
rect 12530 16759 12586 16768
rect 12530 16688 12586 16697
rect 12268 16612 12388 16640
rect 12530 16623 12586 16632
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12268 16250 12296 16458
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12360 16130 12388 16612
rect 12438 16552 12494 16561
rect 12438 16487 12494 16496
rect 12268 16102 12388 16130
rect 12268 15881 12296 16102
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12254 15872 12310 15881
rect 12254 15807 12310 15816
rect 12360 15745 12388 15982
rect 12346 15736 12402 15745
rect 12346 15671 12402 15680
rect 12256 15632 12308 15638
rect 12452 15609 12480 16487
rect 12544 16017 12572 16623
rect 12530 16008 12586 16017
rect 12530 15943 12586 15952
rect 12256 15574 12308 15580
rect 12438 15600 12494 15609
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 15094 12204 15438
rect 12164 15088 12216 15094
rect 12164 15030 12216 15036
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12176 14618 12204 14826
rect 12268 14793 12296 15574
rect 12438 15535 12494 15544
rect 12440 15360 12492 15366
rect 12346 15328 12402 15337
rect 12440 15302 12492 15308
rect 12346 15263 12402 15272
rect 12254 14784 12310 14793
rect 12254 14719 12310 14728
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12360 14550 12388 15263
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12268 13705 12296 14350
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12254 13696 12310 13705
rect 12254 13631 12310 13640
rect 12268 13258 12296 13631
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12176 11898 12204 12786
rect 12268 12714 12296 13194
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12360 12481 12388 13874
rect 12452 12918 12480 15302
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12544 14618 12572 14962
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12636 14006 12664 17682
rect 12728 15638 12756 20295
rect 12820 19446 12848 22918
rect 13004 22438 13032 23190
rect 13372 23118 13400 23734
rect 13464 23322 13492 24142
rect 13648 23866 13676 24754
rect 13740 24585 13768 25842
rect 13832 25673 13860 26200
rect 14200 25974 14228 26200
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 13818 25664 13874 25673
rect 13818 25599 13874 25608
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 13820 24676 13872 24682
rect 13820 24618 13872 24624
rect 13726 24576 13782 24585
rect 13726 24511 13782 24520
rect 13832 24449 13860 24618
rect 13818 24440 13874 24449
rect 13818 24375 13874 24384
rect 13924 23866 13952 25094
rect 14292 25090 14320 26302
rect 14554 26200 14610 26302
rect 14922 26200 14978 27000
rect 15290 26200 15346 27000
rect 15382 26344 15438 26353
rect 15658 26330 15714 27000
rect 15438 26302 15714 26330
rect 15382 26279 15438 26288
rect 15658 26200 15714 26302
rect 16026 26200 16082 27000
rect 16394 26200 16450 27000
rect 16762 26200 16818 27000
rect 17130 26200 17186 27000
rect 17498 26330 17554 27000
rect 17328 26302 17554 26330
rect 14280 25084 14332 25090
rect 14280 25026 14332 25032
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14464 24744 14516 24750
rect 14278 24712 14334 24721
rect 14464 24686 14516 24692
rect 14278 24647 14334 24656
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 14094 23624 14150 23633
rect 14094 23559 14096 23568
rect 14148 23559 14150 23568
rect 14096 23530 14148 23536
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13818 23488 13874 23497
rect 13452 23316 13504 23322
rect 13452 23258 13504 23264
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 13188 22817 13216 22986
rect 13174 22808 13230 22817
rect 13174 22743 13230 22752
rect 13556 22710 13584 23258
rect 13636 23112 13688 23118
rect 13636 23054 13688 23060
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 13648 22642 13676 23054
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13464 22234 13492 22578
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 13004 21622 13032 22034
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 13372 21321 13400 22170
rect 13648 21622 13676 22578
rect 13740 21622 13768 23462
rect 13818 23423 13874 23432
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13452 21412 13504 21418
rect 13452 21354 13504 21360
rect 13358 21312 13414 21321
rect 12950 21244 13258 21253
rect 13358 21247 13414 21256
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 13268 20868 13320 20874
rect 13268 20810 13320 20816
rect 13188 20466 13216 20810
rect 13280 20534 13308 20810
rect 13358 20768 13414 20777
rect 13358 20703 13414 20712
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19938 13400 20703
rect 13464 19990 13492 21354
rect 13648 21185 13676 21558
rect 13726 21312 13782 21321
rect 13726 21247 13782 21256
rect 13634 21176 13690 21185
rect 13634 21111 13690 21120
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13556 20777 13584 20878
rect 13542 20768 13598 20777
rect 13542 20703 13598 20712
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13556 20346 13584 20470
rect 13648 20466 13676 21111
rect 13740 20942 13768 21247
rect 13728 20936 13780 20942
rect 13832 20913 13860 23423
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13924 21690 13952 22374
rect 14016 21894 14044 22510
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13728 20878 13780 20884
rect 13818 20904 13874 20913
rect 13818 20839 13874 20848
rect 13818 20768 13874 20777
rect 13818 20703 13874 20712
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13832 20346 13860 20703
rect 13556 20318 13860 20346
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13726 20224 13782 20233
rect 12912 19910 13400 19938
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12912 19224 12940 19910
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13372 19310 13400 19790
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 12820 19196 12940 19224
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12728 14346 12756 15302
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12820 14226 12848 19196
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 13004 18193 13032 18838
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 13096 18290 13124 18702
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12990 18184 13046 18193
rect 12990 18119 13046 18128
rect 13188 18086 13216 18838
rect 13372 18816 13400 19110
rect 13464 18834 13492 19246
rect 13280 18788 13400 18816
rect 13452 18828 13504 18834
rect 13280 18222 13308 18788
rect 13452 18770 13504 18776
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17610 13400 18634
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13280 17490 13308 17546
rect 13280 17462 13400 17490
rect 13372 17134 13400 17462
rect 13464 17218 13492 18158
rect 13556 17882 13584 20198
rect 13726 20159 13782 20168
rect 13740 19990 13768 20159
rect 13924 19990 13952 21626
rect 14004 21616 14056 21622
rect 14004 21558 14056 21564
rect 14016 20874 14044 21558
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 20534 14044 20810
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 13740 19825 13768 19926
rect 13726 19816 13782 19825
rect 14016 19802 14044 20470
rect 13832 19786 14044 19802
rect 13726 19751 13782 19760
rect 13820 19780 14044 19786
rect 13872 19774 14044 19780
rect 13820 19722 13872 19728
rect 13818 19680 13874 19689
rect 13818 19615 13874 19624
rect 13832 19530 13860 19615
rect 13740 19502 13860 19530
rect 13740 18902 13768 19502
rect 13924 19378 13952 19774
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13648 17678 13676 18770
rect 13832 18290 13860 18770
rect 13924 18578 13952 19314
rect 14016 18766 14044 19654
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13924 18550 14044 18578
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13726 18184 13782 18193
rect 13726 18119 13782 18128
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13740 17513 13768 18119
rect 13726 17504 13782 17513
rect 13726 17439 13782 17448
rect 13464 17190 13676 17218
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13372 16590 13400 17070
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13464 16425 13492 17070
rect 13450 16416 13506 16425
rect 13450 16351 13506 16360
rect 13464 16250 13492 16351
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13268 15088 13320 15094
rect 13372 15076 13400 16118
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13320 15048 13400 15076
rect 13452 15088 13504 15094
rect 13268 15030 13320 15036
rect 13452 15030 13504 15036
rect 13464 14872 13492 15030
rect 13372 14844 13492 14872
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12728 14198 12848 14226
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12438 12608 12494 12617
rect 12438 12543 12494 12552
rect 12346 12472 12402 12481
rect 12256 12436 12308 12442
rect 12346 12407 12402 12416
rect 12256 12378 12308 12384
rect 12268 12186 12296 12378
rect 12268 12158 12388 12186
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12360 11830 12388 12158
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 11992 11206 12112 11234
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11532 7670 11652 7698
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 4185 11192 6598
rect 11532 6458 11560 6734
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11150 4176 11206 4185
rect 11150 4111 11206 4120
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 8668 2382 8720 2388
rect 10138 2408 10194 2417
rect 10138 2343 10194 2352
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 11624 1834 11652 7670
rect 11716 4010 11744 8366
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11900 6390 11928 6598
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11992 6186 12020 11206
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 8566 12112 11018
rect 12452 11014 12480 12543
rect 12544 12442 12572 13874
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12636 13530 12664 13738
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12636 12753 12664 12786
rect 12622 12744 12678 12753
rect 12622 12679 12678 12688
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12530 12336 12586 12345
rect 12530 12271 12586 12280
rect 12164 11008 12216 11014
rect 12440 11008 12492 11014
rect 12164 10950 12216 10956
rect 12346 10976 12402 10985
rect 12176 10810 12204 10950
rect 12440 10950 12492 10956
rect 12346 10911 12402 10920
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 8974 12204 9318
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12162 8120 12218 8129
rect 12162 8055 12164 8064
rect 12216 8055 12218 8064
rect 12164 8026 12216 8032
rect 12268 7546 12296 10746
rect 12360 10266 12388 10911
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 12268 5098 12296 7142
rect 12360 6497 12388 9522
rect 12452 8548 12480 10406
rect 12544 10305 12572 12271
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12530 10296 12586 10305
rect 12530 10231 12586 10240
rect 12636 9042 12664 11086
rect 12728 9466 12756 14198
rect 13188 14074 13216 14350
rect 13372 14346 13400 14844
rect 13556 14770 13584 16050
rect 13648 15722 13676 17190
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13740 16250 13768 16594
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13832 16114 13860 18226
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13924 16182 13952 18022
rect 14016 17184 14044 18550
rect 14108 18426 14136 19246
rect 14200 18601 14228 22170
rect 14292 21894 14320 24647
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14384 22681 14412 22986
rect 14370 22672 14426 22681
rect 14370 22607 14426 22616
rect 14476 22216 14504 24686
rect 14752 24274 14780 24890
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14648 23656 14700 23662
rect 14648 23598 14700 23604
rect 14660 23186 14688 23598
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14648 23180 14700 23186
rect 14648 23122 14700 23128
rect 14554 23080 14610 23089
rect 14554 23015 14556 23024
rect 14608 23015 14610 23024
rect 14556 22986 14608 22992
rect 14660 22438 14688 23122
rect 14844 23089 14872 23462
rect 14830 23080 14886 23089
rect 14740 23044 14792 23050
rect 14830 23015 14886 23024
rect 14740 22986 14792 22992
rect 14752 22778 14780 22986
rect 14936 22953 14964 26200
rect 15304 24562 15332 26200
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15856 24818 15884 25638
rect 16040 25106 16068 26200
rect 15948 25078 16068 25106
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15212 24534 15332 24562
rect 14922 22944 14978 22953
rect 14922 22879 14978 22888
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 15212 22234 15240 24534
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15304 23730 15332 24346
rect 15948 24154 15976 25078
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 15856 24126 15976 24154
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 14384 22188 14504 22216
rect 15200 22228 15252 22234
rect 14384 21962 14412 22188
rect 15200 22170 15252 22176
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14384 21486 14412 21898
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14278 21176 14334 21185
rect 14278 21111 14334 21120
rect 14292 19514 14320 21111
rect 14476 20942 14504 21966
rect 14646 21176 14702 21185
rect 14646 21111 14702 21120
rect 14372 20936 14424 20942
rect 14370 20904 14372 20913
rect 14464 20936 14516 20942
rect 14424 20904 14426 20913
rect 14464 20878 14516 20884
rect 14370 20839 14426 20848
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14292 18766 14320 19450
rect 14384 18970 14412 19722
rect 14476 19174 14504 20878
rect 14554 20088 14610 20097
rect 14554 20023 14610 20032
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14462 19000 14518 19009
rect 14372 18964 14424 18970
rect 14462 18935 14518 18944
rect 14372 18906 14424 18912
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14186 18592 14242 18601
rect 14186 18527 14242 18536
rect 14292 18426 14320 18702
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14200 17746 14228 18226
rect 14292 17746 14320 18362
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14096 17196 14148 17202
rect 14016 17156 14096 17184
rect 14096 17138 14148 17144
rect 14004 16992 14056 16998
rect 14002 16960 14004 16969
rect 14056 16960 14058 16969
rect 14002 16895 14058 16904
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13818 15736 13874 15745
rect 13648 15706 13768 15722
rect 13648 15700 13780 15706
rect 13648 15694 13728 15700
rect 13818 15671 13820 15680
rect 13728 15642 13780 15648
rect 13872 15671 13874 15680
rect 13820 15642 13872 15648
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13464 14742 13584 14770
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12806 13832 12862 13841
rect 12806 13767 12862 13776
rect 12820 12345 12848 13767
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13358 13560 13414 13569
rect 13358 13495 13414 13504
rect 13372 13410 13400 13495
rect 13188 13382 13400 13410
rect 13082 13016 13138 13025
rect 13082 12951 13138 12960
rect 13096 12753 13124 12951
rect 13188 12850 13216 13382
rect 13464 13274 13492 14742
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13372 13246 13492 13274
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13280 12753 13308 13126
rect 13082 12744 13138 12753
rect 13082 12679 13138 12688
rect 13266 12744 13322 12753
rect 13266 12679 13322 12688
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12806 12336 12862 12345
rect 12806 12271 12862 12280
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 11694 13032 12174
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13280 10520 13308 11290
rect 13372 11150 13400 13246
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13464 12238 13492 13126
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13450 11520 13506 11529
rect 13450 11455 13506 11464
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13464 11098 13492 11455
rect 13556 11218 13584 14554
rect 13648 13802 13676 15574
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13740 14074 13768 15302
rect 13832 15162 13860 15506
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13924 13682 13952 15846
rect 13648 13654 13952 13682
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13464 11070 13584 11098
rect 13280 10492 13400 10520
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12728 9438 12848 9466
rect 12716 9376 12768 9382
rect 12714 9344 12716 9353
rect 12768 9344 12770 9353
rect 12714 9279 12770 9288
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12452 8520 12756 8548
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12544 7886 12572 8026
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12346 6488 12402 6497
rect 12346 6423 12402 6432
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12452 4078 12480 6734
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 12544 2038 12572 7278
rect 12636 7002 12664 8366
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12728 6390 12756 8520
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12820 5234 12848 9438
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13280 8498 13308 9114
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12912 7342 12940 7414
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 12898 6624 12954 6633
rect 12898 6559 12954 6568
rect 12912 6458 12940 6559
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 13280 6118 13308 6734
rect 13372 6322 13400 10492
rect 13450 10432 13506 10441
rect 13450 10367 13506 10376
rect 13464 6730 13492 10367
rect 13556 9178 13584 11070
rect 13648 9926 13676 13654
rect 14016 13546 14044 16662
rect 14108 16658 14136 17138
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14094 16280 14150 16289
rect 14094 16215 14150 16224
rect 14108 16046 14136 16215
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14094 15872 14150 15881
rect 14094 15807 14150 15816
rect 14108 15502 14136 15807
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 14482 14136 14826
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 13740 13518 14044 13546
rect 13740 12442 13768 13518
rect 14108 13410 14136 14214
rect 13832 13382 14136 13410
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13832 11336 13860 13382
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13924 12986 13952 13126
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 14094 12744 14150 12753
rect 14094 12679 14150 12688
rect 14002 12472 14058 12481
rect 14002 12407 14058 12416
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11762 13952 12038
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13740 11308 13860 11336
rect 13740 10690 13768 11308
rect 13818 11248 13874 11257
rect 13818 11183 13874 11192
rect 13832 10810 13860 11183
rect 14016 10826 14044 12407
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13924 10798 14044 10826
rect 13740 10662 13860 10690
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13268 6112 13320 6118
rect 13544 6112 13596 6118
rect 13268 6054 13320 6060
rect 13542 6080 13544 6089
rect 13596 6080 13598 6089
rect 12950 6012 13258 6021
rect 13542 6015 13598 6024
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13372 3641 13400 5510
rect 13542 5400 13598 5409
rect 13542 5335 13544 5344
rect 13596 5335 13598 5344
rect 13544 5306 13596 5312
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13556 3942 13584 4014
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13358 3632 13414 3641
rect 13358 3567 13414 3576
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13648 2514 13676 8774
rect 13740 7834 13768 9862
rect 13832 8294 13860 10662
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13924 8090 13952 10798
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10266 14044 10610
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14002 10160 14058 10169
rect 14002 10095 14058 10104
rect 14016 10062 14044 10095
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14108 9654 14136 12679
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14002 8256 14058 8265
rect 14002 8191 14058 8200
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14016 7886 14044 8191
rect 14004 7880 14056 7886
rect 13740 7818 13860 7834
rect 14004 7822 14056 7828
rect 13740 7812 13872 7818
rect 13740 7806 13820 7812
rect 13820 7754 13872 7760
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13740 5710 13768 7686
rect 13820 7336 13872 7342
rect 13818 7304 13820 7313
rect 13872 7304 13874 7313
rect 13818 7239 13874 7248
rect 14200 6322 14228 17206
rect 14292 16658 14320 17682
rect 14370 17232 14426 17241
rect 14370 17167 14426 17176
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14292 14822 14320 15506
rect 14384 15366 14412 17167
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14370 14784 14426 14793
rect 14292 14482 14320 14758
rect 14370 14719 14426 14728
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14292 14074 14320 14418
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14384 13410 14412 14719
rect 14476 14385 14504 18935
rect 14568 15706 14596 20023
rect 14660 18086 14688 21111
rect 14844 20505 14872 22034
rect 15304 21978 15332 22714
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15212 21950 15332 21978
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 14830 20496 14886 20505
rect 14830 20431 14886 20440
rect 15120 20369 15148 21558
rect 15212 20777 15240 21950
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15304 21593 15332 21830
rect 15290 21584 15346 21593
rect 15346 21542 15424 21570
rect 15290 21519 15346 21528
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15198 20768 15254 20777
rect 15198 20703 15254 20712
rect 15106 20360 15162 20369
rect 15106 20295 15162 20304
rect 15108 19984 15160 19990
rect 15108 19926 15160 19932
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14752 19514 14780 19790
rect 15028 19718 15056 19858
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14844 18698 14872 19450
rect 14936 19417 14964 19654
rect 15120 19514 15148 19926
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 14922 19408 14978 19417
rect 14922 19343 14978 19352
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14832 18692 14884 18698
rect 14832 18634 14884 18640
rect 14844 18426 14872 18634
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14660 16998 14688 17274
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14462 14376 14518 14385
rect 14462 14311 14518 14320
rect 14568 14074 14596 15370
rect 14660 15065 14688 16390
rect 14752 15706 14780 17614
rect 14844 16182 14872 18362
rect 15028 17377 15056 19110
rect 15120 18873 15148 19314
rect 15106 18864 15162 18873
rect 15106 18799 15162 18808
rect 15212 18034 15240 20703
rect 15120 18006 15240 18034
rect 15014 17368 15070 17377
rect 15014 17303 15070 17312
rect 14832 16176 14884 16182
rect 14832 16118 14884 16124
rect 15120 16130 15148 18006
rect 15304 17746 15332 21286
rect 15396 20942 15424 21542
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15396 20505 15424 20538
rect 15382 20496 15438 20505
rect 15382 20431 15438 20440
rect 15488 20097 15516 22646
rect 15580 22094 15608 23802
rect 15856 23322 15884 24126
rect 15936 24064 15988 24070
rect 15936 24006 15988 24012
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15948 22642 15976 24006
rect 16040 23769 16068 24890
rect 16212 24132 16264 24138
rect 16212 24074 16264 24080
rect 16120 24064 16172 24070
rect 16120 24006 16172 24012
rect 16026 23760 16082 23769
rect 16026 23695 16082 23704
rect 16026 23216 16082 23225
rect 16026 23151 16082 23160
rect 16040 22642 16068 23151
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15750 22536 15806 22545
rect 15750 22471 15752 22480
rect 15804 22471 15806 22480
rect 15934 22536 15990 22545
rect 15934 22471 15990 22480
rect 15752 22442 15804 22448
rect 15764 22234 15792 22442
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 15580 22066 15792 22094
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15672 21146 15700 21966
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15658 20904 15714 20913
rect 15658 20839 15714 20848
rect 15474 20088 15530 20097
rect 15474 20023 15530 20032
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15474 19816 15530 19825
rect 15474 19751 15530 19760
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 14924 16108 14976 16114
rect 15120 16102 15332 16130
rect 14924 16050 14976 16056
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14646 15056 14702 15065
rect 14752 15026 14780 15642
rect 14646 14991 14702 15000
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14292 13382 14412 13410
rect 14464 13388 14516 13394
rect 14292 13161 14320 13382
rect 14464 13330 14516 13336
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14278 13152 14334 13161
rect 14278 13087 14334 13096
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14292 8498 14320 12922
rect 14384 11898 14412 13262
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14370 11384 14426 11393
rect 14370 11319 14426 11328
rect 14384 8974 14412 11319
rect 14476 10538 14504 13330
rect 14568 12238 14596 13806
rect 14660 12850 14688 14282
rect 14752 13326 14780 14758
rect 14844 13530 14872 14894
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14738 12880 14794 12889
rect 14648 12844 14700 12850
rect 14738 12815 14794 12824
rect 14648 12786 14700 12792
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14554 10568 14610 10577
rect 14464 10532 14516 10538
rect 14554 10503 14610 10512
rect 14464 10474 14516 10480
rect 14568 9586 14596 10503
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14462 8936 14518 8945
rect 14462 8871 14518 8880
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14292 8090 14320 8434
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14476 6662 14504 8871
rect 14568 8498 14596 9046
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14660 7410 14688 12650
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14476 6458 14504 6598
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14568 5710 14596 6938
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 12532 2032 12584 2038
rect 12532 1974 12584 1980
rect 13740 1902 13768 5510
rect 14096 5364 14148 5370
rect 14016 5324 14096 5352
rect 14016 5030 14044 5324
rect 14096 5306 14148 5312
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14292 4078 14320 5646
rect 14752 5370 14780 12815
rect 14936 11898 14964 16050
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 15028 13938 15056 14282
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15120 13870 15148 15982
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15212 13734 15240 14418
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15028 12986 15056 13262
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 15028 11150 15056 12922
rect 15120 12442 15148 13670
rect 15198 13152 15254 13161
rect 15198 13087 15254 13096
rect 15212 12646 15240 13087
rect 15200 12640 15252 12646
rect 15198 12608 15200 12617
rect 15252 12608 15254 12617
rect 15198 12543 15254 12552
rect 15108 12436 15160 12442
rect 15304 12434 15332 16102
rect 15396 13394 15424 19314
rect 15488 17338 15516 19751
rect 15580 19553 15608 19858
rect 15566 19544 15622 19553
rect 15566 19479 15622 19488
rect 15566 19000 15622 19009
rect 15566 18935 15622 18944
rect 15580 18902 15608 18935
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15672 18222 15700 20839
rect 15764 20233 15792 22066
rect 15856 20806 15884 22374
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15750 20224 15806 20233
rect 15750 20159 15806 20168
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15672 18086 15700 18158
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15764 17882 15792 18158
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15856 17610 15884 17818
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15488 13297 15516 17138
rect 15580 15162 15608 17274
rect 15856 17134 15884 17546
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 15658 16688 15714 16697
rect 15658 16623 15714 16632
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15672 15008 15700 16623
rect 15856 16522 15884 17070
rect 15948 16833 15976 22471
rect 16026 22128 16082 22137
rect 16026 22063 16082 22072
rect 16040 21486 16068 22063
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 16040 20942 16068 21422
rect 16132 21321 16160 24006
rect 16224 23225 16252 24074
rect 16304 23248 16356 23254
rect 16210 23216 16266 23225
rect 16304 23190 16356 23196
rect 16210 23151 16266 23160
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16224 21418 16252 22170
rect 16212 21412 16264 21418
rect 16212 21354 16264 21360
rect 16118 21312 16174 21321
rect 16118 21247 16174 21256
rect 16028 20936 16080 20942
rect 16080 20896 16160 20924
rect 16028 20878 16080 20884
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 17202 16068 19790
rect 16132 18426 16160 20896
rect 16210 19272 16266 19281
rect 16210 19207 16266 19216
rect 16224 19174 16252 19207
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16316 18834 16344 23190
rect 16408 21622 16436 26200
rect 16672 26172 16724 26178
rect 16672 26114 16724 26120
rect 16684 24614 16712 26114
rect 16776 26081 16804 26200
rect 16762 26072 16818 26081
rect 16762 26007 16818 26016
rect 16580 24608 16632 24614
rect 16580 24550 16632 24556
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16488 24336 16540 24342
rect 16488 24278 16540 24284
rect 16592 24290 16620 24550
rect 16500 24177 16528 24278
rect 16592 24262 16896 24290
rect 16580 24200 16632 24206
rect 16486 24168 16542 24177
rect 16580 24142 16632 24148
rect 16486 24103 16542 24112
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 16500 21690 16528 23462
rect 16592 23322 16620 24142
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 16500 21486 16528 21626
rect 16488 21480 16540 21486
rect 16394 21448 16450 21457
rect 16684 21457 16712 23054
rect 16488 21422 16540 21428
rect 16670 21448 16726 21457
rect 16394 21383 16450 21392
rect 16670 21383 16726 21392
rect 16408 19281 16436 21383
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16500 20534 16528 20878
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16500 19854 16528 20470
rect 16488 19848 16540 19854
rect 16540 19808 16620 19836
rect 16488 19790 16540 19796
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16500 19417 16528 19654
rect 16486 19408 16542 19417
rect 16486 19343 16542 19352
rect 16394 19272 16450 19281
rect 16394 19207 16450 19216
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16408 18680 16436 19110
rect 16592 18952 16620 19808
rect 16684 19174 16712 21383
rect 16776 20874 16804 24074
rect 16868 22817 16896 24262
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 16960 23050 16988 23598
rect 17040 23588 17092 23594
rect 17040 23530 17092 23536
rect 17052 23118 17080 23530
rect 17144 23497 17172 26200
rect 17328 26178 17356 26302
rect 17498 26200 17554 26302
rect 17866 26200 17922 27000
rect 18234 26330 18290 27000
rect 17972 26302 18290 26330
rect 17316 26172 17368 26178
rect 17316 26114 17368 26120
rect 17684 25016 17736 25022
rect 17684 24958 17736 24964
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17500 24676 17552 24682
rect 17500 24618 17552 24624
rect 17406 24304 17462 24313
rect 17406 24239 17408 24248
rect 17460 24239 17462 24248
rect 17408 24210 17460 24216
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17130 23488 17186 23497
rect 17130 23423 17186 23432
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 17236 23066 17264 24006
rect 17512 23882 17540 24618
rect 17604 24274 17632 24686
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17696 24041 17724 24958
rect 17682 24032 17738 24041
rect 17682 23967 17738 23976
rect 17328 23854 17540 23882
rect 17328 23730 17356 23854
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17500 23180 17552 23186
rect 17500 23122 17552 23128
rect 16948 23044 17000 23050
rect 17236 23038 17356 23066
rect 16948 22986 17000 22992
rect 16854 22808 16910 22817
rect 16960 22778 16988 22986
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17144 22778 17172 22918
rect 16854 22743 16910 22752
rect 16948 22772 17000 22778
rect 16868 22556 16896 22743
rect 16948 22714 17000 22720
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 16960 22658 16988 22714
rect 16960 22630 17172 22658
rect 16948 22568 17000 22574
rect 16868 22528 16948 22556
rect 16948 22510 17000 22516
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16960 20942 16988 21422
rect 17052 21418 17080 22034
rect 17144 22030 17172 22630
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17236 21706 17264 22918
rect 17144 21678 17264 21706
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16776 19922 16804 20810
rect 16856 20800 16908 20806
rect 16854 20768 16856 20777
rect 16908 20768 16910 20777
rect 16854 20703 16910 20712
rect 16960 20534 16988 20878
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 17052 20466 17080 21354
rect 17144 20482 17172 21678
rect 17328 21622 17356 23038
rect 17420 22166 17448 23122
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 17406 21992 17462 22001
rect 17406 21927 17462 21936
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17236 21078 17264 21490
rect 17420 21486 17448 21927
rect 17512 21894 17540 23122
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17590 22808 17646 22817
rect 17590 22743 17646 22752
rect 17604 22574 17632 22743
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17224 21072 17276 21078
rect 17512 21049 17540 21830
rect 17224 21014 17276 21020
rect 17498 21040 17554 21049
rect 17498 20975 17554 20984
rect 17498 20632 17554 20641
rect 17498 20567 17554 20576
rect 17040 20460 17092 20466
rect 17144 20454 17356 20482
rect 17040 20402 17092 20408
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16592 18924 16712 18952
rect 16316 18652 16436 18680
rect 16580 18692 16632 18698
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15934 16824 15990 16833
rect 15934 16759 15990 16768
rect 16040 16726 16068 17138
rect 16132 16969 16160 18158
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16118 16960 16174 16969
rect 16118 16895 16174 16904
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 16132 16538 16160 16662
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 16040 16510 16160 16538
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15580 14980 15700 15008
rect 15474 13288 15530 13297
rect 15474 13223 15530 13232
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15396 12986 15424 13126
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15488 12617 15516 13126
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15304 12406 15424 12434
rect 15108 12378 15160 12384
rect 15292 12368 15344 12374
rect 15290 12336 15292 12345
rect 15344 12336 15346 12345
rect 15290 12271 15346 12280
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15198 11112 15254 11121
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 15108 11076 15160 11082
rect 15198 11047 15254 11056
rect 15108 11018 15160 11024
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14844 9722 14872 10542
rect 14936 9722 14964 11018
rect 15120 10674 15148 11018
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15212 10520 15240 11047
rect 15028 10492 15240 10520
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14844 4486 14872 8298
rect 14936 6254 14964 9522
rect 15028 7546 15056 10492
rect 15198 10432 15254 10441
rect 15198 10367 15254 10376
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15120 8974 15148 9114
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15212 8650 15240 10367
rect 15304 10305 15332 11562
rect 15290 10296 15346 10305
rect 15290 10231 15346 10240
rect 15396 9042 15424 12406
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15488 10742 15516 12310
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15474 9752 15530 9761
rect 15474 9687 15530 9696
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15120 8634 15240 8650
rect 15108 8628 15240 8634
rect 15160 8622 15240 8628
rect 15108 8570 15160 8576
rect 15108 8016 15160 8022
rect 15106 7984 15108 7993
rect 15160 7984 15162 7993
rect 15106 7919 15162 7928
rect 15290 7984 15346 7993
rect 15290 7919 15346 7928
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15212 7546 15240 7822
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15212 6934 15240 7346
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15120 6458 15148 6734
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15304 6322 15332 7919
rect 15382 6760 15438 6769
rect 15382 6695 15438 6704
rect 15396 6662 15424 6695
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15488 6458 15516 9687
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 15580 5370 15608 14980
rect 15764 14618 15792 16050
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15842 15600 15898 15609
rect 15842 15535 15898 15544
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15672 12238 15700 13942
rect 15856 13920 15884 15535
rect 15948 15337 15976 15982
rect 15934 15328 15990 15337
rect 15934 15263 15990 15272
rect 16040 14906 16068 16510
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16132 15201 16160 15302
rect 16118 15192 16174 15201
rect 16118 15127 16174 15136
rect 16132 15094 16160 15127
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16040 14878 16160 14906
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15764 13892 15884 13920
rect 15764 12782 15792 13892
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15660 11348 15712 11354
rect 15856 11336 15884 13738
rect 15948 12986 15976 14418
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15712 11308 15884 11336
rect 15660 11290 15712 11296
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 8974 15700 10406
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15764 5574 15792 8774
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 5710 15884 8230
rect 15948 7546 15976 12922
rect 16040 11762 16068 14554
rect 16132 13818 16160 14878
rect 16224 14482 16252 17070
rect 16316 16726 16344 18652
rect 16580 18634 16632 18640
rect 16488 18216 16540 18222
rect 16486 18184 16488 18193
rect 16540 18184 16542 18193
rect 16396 18148 16448 18154
rect 16486 18119 16542 18128
rect 16396 18090 16448 18096
rect 16304 16720 16356 16726
rect 16304 16662 16356 16668
rect 16408 16561 16436 18090
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 16833 16528 18022
rect 16592 17882 16620 18634
rect 16684 18630 16712 18924
rect 16776 18816 16804 19110
rect 16856 18828 16908 18834
rect 16776 18788 16856 18816
rect 16672 18624 16724 18630
rect 16776 18601 16804 18788
rect 16856 18770 16908 18776
rect 16856 18624 16908 18630
rect 16672 18566 16724 18572
rect 16762 18592 16818 18601
rect 16684 18426 16712 18566
rect 16856 18566 16908 18572
rect 16762 18527 16818 18536
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16684 17610 16712 18362
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16684 17270 16712 17546
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16486 16824 16542 16833
rect 16486 16759 16542 16768
rect 16394 16552 16450 16561
rect 16394 16487 16450 16496
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16316 15978 16344 16118
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16316 13938 16344 15438
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16132 13790 16344 13818
rect 16118 13560 16174 13569
rect 16118 13495 16174 13504
rect 16132 13161 16160 13495
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16118 13152 16174 13161
rect 16118 13087 16174 13096
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16132 10538 16160 12038
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16040 10130 16068 10406
rect 16224 10198 16252 13194
rect 16316 13002 16344 13790
rect 16408 13161 16436 15982
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16500 15638 16528 15846
rect 16578 15736 16634 15745
rect 16578 15671 16580 15680
rect 16632 15671 16634 15680
rect 16580 15642 16632 15648
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16684 15434 16712 16934
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16394 13152 16450 13161
rect 16394 13087 16450 13096
rect 16316 12974 16436 13002
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16316 11898 16344 12786
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16316 9586 16344 11698
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16118 8664 16174 8673
rect 16118 8599 16174 8608
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15948 6118 15976 6734
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 16040 5817 16068 6598
rect 16132 6458 16160 8599
rect 16304 8424 16356 8430
rect 16302 8392 16304 8401
rect 16356 8392 16358 8401
rect 16302 8327 16358 8336
rect 16408 7886 16436 12974
rect 16500 12102 16528 14826
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 14278 16620 14758
rect 16670 14648 16726 14657
rect 16776 14618 16804 17682
rect 16868 17134 16896 18566
rect 16960 17882 16988 19382
rect 17052 19378 17080 20402
rect 17132 20324 17184 20330
rect 17132 20266 17184 20272
rect 17144 20058 17172 20266
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17038 19000 17094 19009
rect 17038 18935 17094 18944
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16960 16697 16988 17478
rect 16946 16688 17002 16697
rect 16856 16652 16908 16658
rect 16946 16623 17002 16632
rect 16856 16594 16908 16600
rect 16868 14822 16896 16594
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 15910 16988 16526
rect 17052 16289 17080 18935
rect 17144 18290 17172 19858
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17236 17882 17264 19790
rect 17328 19009 17356 20454
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17314 19000 17370 19009
rect 17314 18935 17370 18944
rect 17420 18465 17448 20334
rect 17512 20097 17540 20567
rect 17498 20088 17554 20097
rect 17498 20023 17554 20032
rect 17512 18986 17540 20023
rect 17604 19854 17632 22510
rect 17696 21690 17724 22918
rect 17788 22506 17816 23462
rect 17880 23322 17908 26200
rect 17972 25294 18000 26302
rect 18234 26200 18290 26302
rect 18602 26200 18658 27000
rect 18970 26330 19026 27000
rect 18970 26302 19288 26330
rect 18970 26200 19026 26302
rect 18616 25809 18644 26200
rect 18602 25800 18658 25809
rect 18602 25735 18658 25744
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 18142 24848 18198 24857
rect 18142 24783 18198 24792
rect 18156 24410 18184 24783
rect 19064 24676 19116 24682
rect 19064 24618 19116 24624
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23798 18368 24346
rect 18972 24336 19024 24342
rect 19076 24313 19104 24618
rect 18972 24278 19024 24284
rect 19062 24304 19118 24313
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18616 23866 18644 24006
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17776 22500 17828 22506
rect 17776 22442 17828 22448
rect 17776 22160 17828 22166
rect 17776 22102 17828 22108
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17788 21010 17816 22102
rect 17880 22030 17908 22646
rect 18236 22500 18288 22506
rect 18064 22460 18236 22488
rect 18064 22098 18092 22460
rect 18236 22442 18288 22448
rect 18142 22128 18198 22137
rect 18052 22092 18104 22098
rect 18142 22063 18198 22072
rect 18052 22034 18104 22040
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 18156 21894 18184 22063
rect 18236 22024 18288 22030
rect 18234 21992 18236 22001
rect 18288 21992 18290 22001
rect 18234 21927 18290 21936
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18340 21554 18368 23462
rect 18418 23216 18474 23225
rect 18418 23151 18474 23160
rect 18432 22778 18460 23151
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18432 22030 18460 22442
rect 18524 22094 18552 23802
rect 18694 23760 18750 23769
rect 18694 23695 18750 23704
rect 18708 23254 18736 23695
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18696 23248 18748 23254
rect 18696 23190 18748 23196
rect 18602 22808 18658 22817
rect 18602 22743 18658 22752
rect 18616 22642 18644 22743
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18524 22066 18736 22094
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18602 21720 18658 21729
rect 18602 21655 18658 21664
rect 18616 21622 18644 21655
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17592 19712 17644 19718
rect 17590 19680 17592 19689
rect 17644 19680 17646 19689
rect 17590 19615 17646 19624
rect 17696 19514 17724 20742
rect 17774 20224 17830 20233
rect 17774 20159 17830 20168
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 17512 18958 17632 18986
rect 17604 18902 17632 18958
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17406 18456 17462 18465
rect 17406 18391 17462 18400
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17222 17776 17278 17785
rect 17222 17711 17278 17720
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17038 16280 17094 16289
rect 17038 16215 17094 16224
rect 16948 15904 17000 15910
rect 16946 15872 16948 15881
rect 17040 15904 17092 15910
rect 17000 15872 17002 15881
rect 17040 15846 17092 15852
rect 16946 15807 17002 15816
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16670 14583 16726 14592
rect 16764 14612 16816 14618
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16684 14113 16712 14583
rect 16764 14554 16816 14560
rect 16670 14104 16726 14113
rect 16670 14039 16726 14048
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16592 12986 16620 13874
rect 16868 13410 16896 14758
rect 16684 13394 16896 13410
rect 16672 13388 16896 13394
rect 16724 13382 16896 13388
rect 16672 13330 16724 13336
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16684 12434 16712 13126
rect 16868 12850 16896 13382
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16592 12406 16712 12434
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16500 10130 16528 11834
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16592 10062 16620 12406
rect 16762 12336 16818 12345
rect 16868 12306 16896 12786
rect 16762 12271 16764 12280
rect 16816 12271 16818 12280
rect 16856 12300 16908 12306
rect 16764 12242 16816 12248
rect 16856 12242 16908 12248
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16684 10810 16712 12174
rect 16960 12102 16988 15438
rect 17052 15094 17080 15846
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 17052 13870 17080 14282
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17052 13326 17080 13806
rect 17144 13530 17172 17002
rect 17236 16969 17264 17711
rect 17420 16998 17448 17818
rect 17408 16992 17460 16998
rect 17222 16960 17278 16969
rect 17408 16934 17460 16940
rect 17222 16895 17278 16904
rect 17222 15600 17278 15609
rect 17222 15535 17224 15544
rect 17276 15535 17278 15544
rect 17224 15506 17276 15512
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17236 14770 17264 14894
rect 17236 14742 17356 14770
rect 17222 13696 17278 13705
rect 17222 13631 17278 13640
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17040 13320 17092 13326
rect 17092 13280 17172 13308
rect 17040 13262 17092 13268
rect 17144 12918 17172 13280
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 16948 12096 17000 12102
rect 16762 12064 16818 12073
rect 16948 12038 17000 12044
rect 16762 11999 16818 12008
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16224 7274 16252 7686
rect 16408 7546 16436 7822
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16592 7478 16620 9318
rect 16684 9178 16712 9318
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8498 16712 8910
rect 16776 8634 16804 11999
rect 16856 11688 16908 11694
rect 16854 11656 16856 11665
rect 16908 11656 16910 11665
rect 16854 11591 16910 11600
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11098 16896 11494
rect 16960 11218 16988 12038
rect 17052 11762 17080 12242
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17038 11248 17094 11257
rect 16948 11212 17000 11218
rect 17144 11218 17172 12854
rect 17236 11898 17264 13631
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17328 11608 17356 14742
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17236 11580 17356 11608
rect 17038 11183 17094 11192
rect 17132 11212 17184 11218
rect 16948 11154 17000 11160
rect 16868 11070 16988 11098
rect 16960 11014 16988 11070
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16868 9178 16896 10950
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16960 10062 16988 10406
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16868 8090 16896 8230
rect 16960 8090 16988 9454
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16578 7304 16634 7313
rect 16212 7268 16264 7274
rect 16578 7239 16634 7248
rect 16212 7210 16264 7216
rect 16592 6798 16620 7239
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16026 5808 16082 5817
rect 16026 5743 16082 5752
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 16224 4758 16252 6734
rect 16302 5808 16358 5817
rect 16302 5743 16358 5752
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 16316 4622 16344 5743
rect 16684 5409 16712 7686
rect 16776 7342 16804 7754
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16776 5914 16804 6598
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16670 5400 16726 5409
rect 16670 5335 16726 5344
rect 16486 5128 16542 5137
rect 16396 5092 16448 5098
rect 16486 5063 16488 5072
rect 16396 5034 16448 5040
rect 16540 5063 16542 5072
rect 16488 5034 16540 5040
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 15028 2106 15056 4558
rect 16316 4282 16344 4558
rect 16408 4282 16436 5034
rect 16500 4622 16528 5034
rect 16868 4826 16896 7278
rect 17052 6474 17080 11183
rect 17132 11154 17184 11160
rect 17236 10742 17264 11580
rect 17420 11506 17448 14554
rect 17328 11478 17448 11506
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17328 10674 17356 11478
rect 17512 11234 17540 18770
rect 17788 18630 17816 20159
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17604 18222 17632 18566
rect 17880 18222 17908 21286
rect 18248 20874 18276 21490
rect 18340 21418 18368 21490
rect 18328 21412 18380 21418
rect 18328 21354 18380 21360
rect 18340 21010 18368 21354
rect 18708 21146 18736 22066
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18326 19952 18382 19961
rect 18326 19887 18328 19896
rect 18380 19887 18382 19896
rect 18328 19858 18380 19864
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18432 19009 18460 20334
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18524 19786 18552 20198
rect 18512 19780 18564 19786
rect 18512 19722 18564 19728
rect 18418 19000 18474 19009
rect 18418 18935 18474 18944
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18432 18358 18460 18566
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17604 17202 17632 17818
rect 17682 17776 17738 17785
rect 17682 17711 17738 17720
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17590 16688 17646 16697
rect 17590 16623 17646 16632
rect 17604 15706 17632 16623
rect 17696 16522 17724 17711
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17604 14521 17632 15642
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17696 15094 17724 15370
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17590 14512 17646 14521
rect 17590 14447 17646 14456
rect 17590 14376 17646 14385
rect 17590 14311 17646 14320
rect 17604 13025 17632 14311
rect 17696 13870 17724 15030
rect 17788 14618 17816 18158
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17972 16833 18000 17070
rect 17958 16824 18014 16833
rect 17958 16759 18014 16768
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17880 14550 17908 16594
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18340 16250 18368 18294
rect 18420 18080 18472 18086
rect 18524 18057 18552 18566
rect 18420 18022 18472 18028
rect 18510 18048 18566 18057
rect 18432 17762 18460 18022
rect 18510 17983 18566 17992
rect 18432 17734 18552 17762
rect 18616 17746 18644 21082
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 19145 18736 19654
rect 18694 19136 18750 19145
rect 18694 19071 18750 19080
rect 18800 18766 18828 23598
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18892 23050 18920 23190
rect 18984 23118 19012 24278
rect 19062 24239 19118 24248
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 19062 23080 19118 23089
rect 18880 23044 18932 23050
rect 19062 23015 19118 23024
rect 18880 22986 18932 22992
rect 18892 22545 18920 22986
rect 18972 22568 19024 22574
rect 18878 22536 18934 22545
rect 18972 22510 19024 22516
rect 18878 22471 18934 22480
rect 18878 22128 18934 22137
rect 18878 22063 18934 22072
rect 18892 21962 18920 22063
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18984 21350 19012 22510
rect 19076 22166 19104 23015
rect 19156 22500 19208 22506
rect 19156 22442 19208 22448
rect 19064 22160 19116 22166
rect 19064 22102 19116 22108
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18984 20262 19012 21286
rect 19076 21010 19104 21966
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 19076 19922 19104 20742
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18420 17604 18472 17610
rect 18420 17546 18472 17552
rect 18432 17202 18460 17546
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17972 15065 18000 15098
rect 17958 15056 18014 15065
rect 17958 14991 18014 15000
rect 17868 14544 17920 14550
rect 17774 14512 17830 14521
rect 17868 14486 17920 14492
rect 17774 14447 17830 14456
rect 17788 14396 17816 14447
rect 17788 14368 17908 14396
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17590 13016 17646 13025
rect 17590 12951 17646 12960
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17696 12434 17724 12718
rect 17420 11218 17540 11234
rect 17408 11212 17540 11218
rect 17460 11206 17540 11212
rect 17604 12406 17724 12434
rect 17408 11154 17460 11160
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17144 9382 17172 10066
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17236 8974 17264 9522
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 8974 17356 9318
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17052 6446 17172 6474
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16946 5944 17002 5953
rect 16946 5879 16948 5888
rect 17000 5879 17002 5888
rect 16948 5850 17000 5856
rect 17052 5234 17080 6326
rect 17144 5710 17172 6446
rect 17236 6254 17264 6734
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17144 5030 17172 5646
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17130 4856 17186 4865
rect 16856 4820 16908 4826
rect 17130 4791 17132 4800
rect 16856 4762 16908 4768
rect 17184 4791 17186 4800
rect 17132 4762 17184 4768
rect 17144 4622 17172 4762
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16960 4010 16988 4082
rect 17052 4049 17080 4082
rect 17038 4040 17094 4049
rect 16948 4004 17000 4010
rect 17038 3975 17094 3984
rect 16948 3946 17000 3952
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 17328 1970 17356 8366
rect 17420 7886 17448 11154
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17512 10849 17540 10950
rect 17498 10840 17554 10849
rect 17498 10775 17554 10784
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17420 4808 17448 7482
rect 17512 6866 17540 9862
rect 17604 8838 17632 12406
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17696 9654 17724 11630
rect 17788 10810 17816 14214
rect 17880 14074 17908 14368
rect 18340 14346 18368 16186
rect 18432 16182 18460 16594
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 18432 16017 18460 16118
rect 18418 16008 18474 16017
rect 18418 15943 18474 15952
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 18340 14006 18368 14282
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18340 13682 18368 13806
rect 18432 13802 18460 14214
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18340 13654 18460 13682
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17880 12481 17908 13466
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17866 12472 17922 12481
rect 17866 12407 17922 12416
rect 18340 12374 18368 13126
rect 18328 12368 18380 12374
rect 18328 12310 18380 12316
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17866 11792 17922 11801
rect 17866 11727 17922 11736
rect 18050 11792 18106 11801
rect 18432 11762 18460 13654
rect 18524 13258 18552 17734
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18616 14618 18644 17206
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18616 13025 18644 14010
rect 18602 13016 18658 13025
rect 18602 12951 18658 12960
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18510 12336 18566 12345
rect 18510 12271 18566 12280
rect 18524 12238 18552 12271
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18050 11727 18106 11736
rect 18420 11756 18472 11762
rect 17880 11150 17908 11727
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17868 11144 17920 11150
rect 17972 11121 18000 11154
rect 17868 11086 17920 11092
rect 17958 11112 18014 11121
rect 17958 11047 18014 11056
rect 18064 11014 18092 11727
rect 18420 11698 18472 11704
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18524 11393 18552 11562
rect 18510 11384 18566 11393
rect 18510 11319 18566 11328
rect 18524 11286 18552 11319
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18326 11112 18382 11121
rect 18326 11047 18382 11056
rect 18420 11076 18472 11082
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17788 9432 17816 10474
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9586 17908 9862
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17696 9404 17816 9432
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17604 6118 17632 8366
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17604 5370 17632 5578
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17498 5264 17554 5273
rect 17498 5199 17554 5208
rect 17592 5228 17644 5234
rect 17512 5098 17540 5199
rect 17592 5170 17644 5176
rect 17604 5098 17632 5170
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 17592 5092 17644 5098
rect 17592 5034 17644 5040
rect 17420 4780 17632 4808
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17420 2650 17448 4626
rect 17498 4312 17554 4321
rect 17498 4247 17554 4256
rect 17512 4078 17540 4247
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17604 3194 17632 4780
rect 17696 3670 17724 9404
rect 17972 9178 18000 9522
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18064 8906 18092 9386
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17972 8090 18000 8434
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 7002 18092 7278
rect 18156 7002 18184 7346
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17774 6488 17830 6497
rect 17950 6491 18258 6500
rect 17774 6423 17830 6432
rect 17788 6322 17816 6423
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5710 18276 6054
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 17788 4078 17816 5578
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17960 5364 18012 5370
rect 17880 5324 17960 5352
rect 17880 5098 17908 5324
rect 17960 5306 18012 5312
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17972 4978 18000 5170
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17880 4950 18000 4978
rect 17880 4486 17908 4950
rect 17958 4584 18014 4593
rect 18064 4554 18092 5102
rect 17958 4519 18014 4528
rect 18052 4548 18104 4554
rect 17972 4486 18000 4519
rect 18052 4490 18104 4496
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 18248 3942 18276 4082
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18234 3768 18290 3777
rect 18340 3738 18368 11047
rect 18420 11018 18472 11024
rect 18432 7324 18460 11018
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18524 10674 18552 10950
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 7546 18552 10406
rect 18616 9518 18644 12718
rect 18708 11830 18736 17206
rect 18800 16658 18828 18566
rect 18892 18442 18920 19790
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18984 18873 19012 19654
rect 19076 18970 19104 19858
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18970 18864 19026 18873
rect 18970 18799 19026 18808
rect 19168 18698 19196 22442
rect 19260 22094 19288 26302
rect 19338 26200 19394 27000
rect 19614 26208 19670 26217
rect 19352 24818 19380 26200
rect 19706 26200 19762 27000
rect 20074 26200 20130 27000
rect 20350 26888 20406 26897
rect 20442 26874 20498 27000
rect 20406 26846 20498 26874
rect 20350 26823 20406 26832
rect 20442 26200 20498 26846
rect 20810 26200 20866 27000
rect 21178 26330 21234 27000
rect 21546 26330 21602 27000
rect 20916 26302 21234 26330
rect 19614 26143 19670 26152
rect 19628 26058 19656 26143
rect 19720 26058 19748 26200
rect 19628 26030 19748 26058
rect 20088 25945 20116 26200
rect 20074 25936 20130 25945
rect 20074 25871 20130 25880
rect 20536 25628 20588 25634
rect 20536 25570 20588 25576
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19444 24313 19472 24346
rect 19430 24304 19486 24313
rect 19430 24239 19486 24248
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19352 23633 19380 24006
rect 19338 23624 19394 23633
rect 19338 23559 19394 23568
rect 19536 22098 19564 25298
rect 19616 24948 19668 24954
rect 19616 24890 19668 24896
rect 19628 24410 19656 24890
rect 19984 24880 20036 24886
rect 19984 24822 20036 24828
rect 19996 24410 20024 24822
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19720 23662 19748 24210
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19812 23526 19840 24210
rect 19996 24138 20024 24346
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 19984 24132 20036 24138
rect 19984 24074 20036 24080
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19720 22681 19748 22986
rect 19706 22672 19762 22681
rect 19616 22636 19668 22642
rect 19706 22607 19762 22616
rect 19616 22578 19668 22584
rect 19628 22545 19656 22578
rect 19614 22536 19670 22545
rect 19614 22471 19670 22480
rect 19260 22066 19380 22094
rect 19248 21072 19300 21078
rect 19248 21014 19300 21020
rect 19260 20618 19288 21014
rect 19352 20754 19380 22066
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19524 22092 19576 22098
rect 19524 22034 19576 22040
rect 19444 21894 19472 22034
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19352 20726 19564 20754
rect 19260 20590 19472 20618
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19352 20262 19380 20402
rect 19444 20398 19472 20590
rect 19536 20505 19564 20726
rect 19522 20496 19578 20505
rect 19522 20431 19578 20440
rect 19432 20392 19484 20398
rect 19628 20369 19656 22471
rect 19812 22094 19840 23462
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 19996 22137 20024 22170
rect 19720 22066 19840 22094
rect 19982 22128 20038 22137
rect 19720 21418 19748 22066
rect 19982 22063 20038 22072
rect 20088 21894 20116 23462
rect 20180 23050 20208 23734
rect 20272 23322 20300 24278
rect 20548 24070 20576 25570
rect 20718 24168 20774 24177
rect 20718 24103 20774 24112
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20732 23798 20760 24103
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 20732 23322 20760 23598
rect 20824 23361 20852 26200
rect 20916 25770 20944 26302
rect 21178 26200 21234 26302
rect 21284 26302 21602 26330
rect 21284 26246 21312 26302
rect 21272 26240 21324 26246
rect 21546 26200 21602 26302
rect 21914 26200 21970 27000
rect 22282 26330 22338 27000
rect 22204 26314 22338 26330
rect 22560 26376 22612 26382
rect 22560 26318 22612 26324
rect 22192 26308 22338 26314
rect 22244 26302 22338 26308
rect 22192 26250 22244 26256
rect 22282 26200 22338 26302
rect 21272 26182 21324 26188
rect 21732 25832 21784 25838
rect 21732 25774 21784 25780
rect 20904 25764 20956 25770
rect 20904 25706 20956 25712
rect 20994 25392 21050 25401
rect 20994 25327 21050 25336
rect 21008 23662 21036 25327
rect 21638 25120 21694 25129
rect 21638 25055 21694 25064
rect 21180 24676 21232 24682
rect 21180 24618 21232 24624
rect 21192 24342 21220 24618
rect 21180 24336 21232 24342
rect 21180 24278 21232 24284
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20916 23497 20944 23598
rect 21088 23588 21140 23594
rect 21088 23530 21140 23536
rect 20902 23488 20958 23497
rect 20902 23423 20958 23432
rect 20810 23352 20866 23361
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 20720 23316 20772 23322
rect 20810 23287 20866 23296
rect 20720 23258 20772 23264
rect 20168 23044 20220 23050
rect 20168 22986 20220 22992
rect 20076 21888 20128 21894
rect 19798 21856 19854 21865
rect 20076 21830 20128 21836
rect 19798 21791 19854 21800
rect 19708 21412 19760 21418
rect 19708 21354 19760 21360
rect 19706 20904 19762 20913
rect 19706 20839 19708 20848
rect 19760 20839 19762 20848
rect 19708 20810 19760 20816
rect 19432 20334 19484 20340
rect 19614 20360 19670 20369
rect 19340 20256 19392 20262
rect 19338 20224 19340 20233
rect 19392 20224 19394 20233
rect 19338 20159 19394 20168
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19156 18692 19208 18698
rect 19156 18634 19208 18640
rect 18892 18414 19012 18442
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18892 17746 18920 18294
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18800 16250 18828 16390
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18892 15638 18920 16390
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18892 14414 18920 14826
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18696 11824 18748 11830
rect 18696 11766 18748 11772
rect 18800 11642 18828 13398
rect 18984 13274 19012 18414
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 19076 17134 19104 17614
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19076 15366 19104 16050
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 18892 13246 19012 13274
rect 18892 12866 18920 13246
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12986 19012 13126
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18892 12838 19012 12866
rect 18880 12640 18932 12646
rect 18878 12608 18880 12617
rect 18932 12608 18934 12617
rect 18878 12543 18934 12552
rect 18984 12434 19012 12838
rect 18708 11614 18828 11642
rect 18892 12406 19012 12434
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18616 9110 18644 9318
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18616 8634 18644 8910
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18432 7296 18644 7324
rect 18418 7168 18474 7177
rect 18418 7103 18474 7112
rect 18432 5914 18460 7103
rect 18616 6118 18644 7296
rect 18708 6390 18736 11614
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 8498 18828 11494
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18892 8430 18920 12406
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18984 11694 19012 12310
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 18984 10441 19012 10746
rect 18970 10432 19026 10441
rect 18970 10367 19026 10376
rect 18984 10266 19012 10367
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18970 10160 19026 10169
rect 18970 10095 19026 10104
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18892 6390 18920 8026
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18604 6112 18656 6118
rect 18510 6080 18566 6089
rect 18604 6054 18656 6060
rect 18510 6015 18566 6024
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18524 5302 18552 6015
rect 18616 5574 18644 6054
rect 18878 5672 18934 5681
rect 18878 5607 18880 5616
rect 18932 5607 18934 5616
rect 18880 5578 18932 5584
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18984 5370 19012 10095
rect 19076 9722 19104 15302
rect 19168 15076 19196 18090
rect 19260 15201 19288 19110
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19246 15192 19302 15201
rect 19246 15127 19302 15136
rect 19168 15048 19288 15076
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19168 12753 19196 12854
rect 19154 12744 19210 12753
rect 19154 12679 19210 12688
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 11354 19196 12582
rect 19260 11558 19288 15048
rect 19352 15042 19380 18838
rect 19444 18290 19472 20334
rect 19614 20295 19670 20304
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 17814 19472 18226
rect 19536 18086 19564 19654
rect 19628 19514 19656 20198
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19614 18864 19670 18873
rect 19614 18799 19670 18808
rect 19628 18766 19656 18799
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19524 18080 19576 18086
rect 19720 18057 19748 18566
rect 19524 18022 19576 18028
rect 19706 18048 19762 18057
rect 19706 17983 19762 17992
rect 19812 17898 19840 21791
rect 20180 21622 20208 22986
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20548 22778 20576 22918
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20810 22672 20866 22681
rect 20810 22607 20812 22616
rect 20864 22607 20866 22616
rect 20812 22578 20864 22584
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 20352 22160 20404 22166
rect 20350 22128 20352 22137
rect 20404 22128 20406 22137
rect 20350 22063 20406 22072
rect 20534 21992 20590 22001
rect 20732 21978 20760 22442
rect 20916 22234 21036 22250
rect 20916 22228 21048 22234
rect 20916 22222 20996 22228
rect 20732 21950 20852 21978
rect 20534 21927 20590 21936
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20168 21616 20220 21622
rect 20074 21584 20130 21593
rect 20168 21558 20220 21564
rect 20074 21519 20130 21528
rect 20088 21486 20116 21519
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 19904 20641 19932 21354
rect 20180 21350 20208 21558
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 19890 20632 19946 20641
rect 19890 20567 19946 20576
rect 20180 20534 20208 21286
rect 20456 21010 20484 21626
rect 20260 21004 20312 21010
rect 20260 20946 20312 20952
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 19996 19145 20024 19178
rect 19982 19136 20038 19145
rect 19982 19071 20038 19080
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19628 17870 19840 17898
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19524 16176 19576 16182
rect 19524 16118 19576 16124
rect 19430 15464 19486 15473
rect 19430 15399 19432 15408
rect 19484 15399 19486 15408
rect 19432 15370 19484 15376
rect 19536 15178 19564 16118
rect 19628 16046 19656 17870
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19720 16182 19748 16458
rect 19812 16454 19840 17138
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 19708 16176 19760 16182
rect 19708 16118 19760 16124
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19628 15570 19656 15982
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19616 15360 19668 15366
rect 19614 15328 19616 15337
rect 19800 15360 19852 15366
rect 19668 15328 19670 15337
rect 19800 15302 19852 15308
rect 19614 15263 19670 15272
rect 19536 15150 19656 15178
rect 19352 15014 19472 15042
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19352 14074 19380 14894
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19352 11762 19380 13330
rect 19444 13161 19472 15014
rect 19522 13288 19578 13297
rect 19522 13223 19524 13232
rect 19576 13223 19578 13232
rect 19524 13194 19576 13200
rect 19430 13152 19486 13161
rect 19430 13087 19486 13096
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19430 12608 19486 12617
rect 19430 12543 19486 12552
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19338 11248 19394 11257
rect 19338 11183 19394 11192
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19168 10674 19196 11018
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19260 10062 19288 10950
rect 19352 10305 19380 11183
rect 19444 10577 19472 12543
rect 19430 10568 19486 10577
rect 19430 10503 19486 10512
rect 19430 10432 19486 10441
rect 19430 10367 19486 10376
rect 19338 10296 19394 10305
rect 19338 10231 19340 10240
rect 19392 10231 19394 10240
rect 19340 10202 19392 10208
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19156 9988 19208 9994
rect 19156 9930 19208 9936
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19076 9382 19104 9522
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 9178 19104 9318
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 19076 8294 19104 8978
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19168 8090 19196 9930
rect 19444 9908 19472 10367
rect 19260 9880 19472 9908
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19260 7970 19288 9880
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19076 7942 19288 7970
rect 19076 5817 19104 7942
rect 19246 7848 19302 7857
rect 19246 7783 19302 7792
rect 19260 7410 19288 7783
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19260 6934 19288 7346
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19062 5808 19118 5817
rect 19062 5743 19118 5752
rect 19062 5672 19118 5681
rect 19168 5642 19196 6802
rect 19062 5607 19118 5616
rect 19156 5636 19208 5642
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18696 4548 18748 4554
rect 18696 4490 18748 4496
rect 18708 4214 18736 4490
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18616 3913 18644 4082
rect 18878 4040 18934 4049
rect 18878 3975 18934 3984
rect 18602 3904 18658 3913
rect 18602 3839 18658 3848
rect 18234 3703 18290 3712
rect 18328 3732 18380 3738
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 18248 3534 18276 3703
rect 18328 3674 18380 3680
rect 18892 3534 18920 3975
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 19076 3097 19104 5607
rect 19156 5578 19208 5584
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19260 4758 19288 4966
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19156 4208 19208 4214
rect 19156 4150 19208 4156
rect 19168 4010 19196 4150
rect 19352 4146 19380 8366
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19444 7886 19472 8230
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19062 3088 19118 3097
rect 19062 3023 19118 3032
rect 19444 2961 19472 3878
rect 19536 3602 19564 12922
rect 19628 12170 19656 15150
rect 19812 14482 19840 15302
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19720 12481 19748 13126
rect 19706 12472 19762 12481
rect 19706 12407 19762 12416
rect 19616 12164 19668 12170
rect 19616 12106 19668 12112
rect 19614 12064 19670 12073
rect 19614 11999 19670 12008
rect 19628 11393 19656 11999
rect 19614 11384 19670 11393
rect 19614 11319 19670 11328
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19628 8566 19656 8978
rect 19616 8560 19668 8566
rect 19616 8502 19668 8508
rect 19720 6440 19748 11222
rect 19812 8566 19840 14214
rect 19904 13190 19932 18906
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19996 15570 20024 17614
rect 20088 15570 20116 20198
rect 20180 17338 20208 20266
rect 20272 18834 20300 20946
rect 20442 20632 20498 20641
rect 20442 20567 20498 20576
rect 20456 19802 20484 20567
rect 20548 19854 20576 21927
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20626 21312 20682 21321
rect 20626 21247 20682 21256
rect 20640 20602 20668 21247
rect 20732 20874 20760 21830
rect 20720 20868 20772 20874
rect 20720 20810 20772 20816
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20364 19774 20484 19802
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20272 18358 20300 18770
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19996 15076 20024 15506
rect 20168 15428 20220 15434
rect 20168 15370 20220 15376
rect 20076 15088 20128 15094
rect 19996 15048 20076 15076
rect 20076 15030 20128 15036
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19892 11824 19944 11830
rect 19892 11766 19944 11772
rect 19904 9178 19932 11766
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19996 6662 20024 13194
rect 20088 10470 20116 13806
rect 20180 12889 20208 15370
rect 20272 13569 20300 16186
rect 20364 14657 20392 19774
rect 20732 19718 20760 20810
rect 20824 20097 20852 21950
rect 20916 21185 20944 22222
rect 20996 22170 21048 22176
rect 21100 22094 21128 23530
rect 21008 22066 21128 22094
rect 20902 21176 20958 21185
rect 20902 21111 20958 21120
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20810 20088 20866 20097
rect 20810 20023 20866 20032
rect 20916 19938 20944 20402
rect 20824 19910 20944 19938
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20456 19281 20484 19654
rect 20732 19378 20760 19654
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20442 19272 20498 19281
rect 20498 19230 20576 19258
rect 20442 19207 20498 19216
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20350 14648 20406 14657
rect 20350 14583 20406 14592
rect 20364 14074 20392 14583
rect 20456 14414 20484 19110
rect 20548 18834 20576 19230
rect 20824 19174 20852 19910
rect 21008 19514 21036 22066
rect 21180 21480 21232 21486
rect 21284 21457 21312 24074
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21376 21865 21404 23666
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21454 22808 21510 22817
rect 21454 22743 21510 22752
rect 21468 22642 21496 22743
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21560 22574 21588 23462
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21362 21856 21418 21865
rect 21362 21791 21418 21800
rect 21376 21486 21404 21791
rect 21652 21622 21680 25055
rect 21744 24410 21772 25774
rect 21928 24993 21956 26200
rect 22572 26058 22600 26318
rect 22650 26200 22706 27000
rect 23018 26330 23074 27000
rect 22756 26302 23074 26330
rect 22664 26058 22692 26200
rect 22572 26030 22692 26058
rect 22008 25560 22060 25566
rect 22008 25502 22060 25508
rect 21914 24984 21970 24993
rect 21914 24919 21970 24928
rect 22020 24721 22048 25502
rect 22006 24712 22062 24721
rect 22006 24647 22062 24656
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 22466 24576 22522 24585
rect 21822 24440 21878 24449
rect 21732 24404 21784 24410
rect 21822 24375 21878 24384
rect 21732 24346 21784 24352
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21364 21480 21416 21486
rect 21180 21422 21232 21428
rect 21270 21448 21326 21457
rect 21192 20466 21220 21422
rect 21364 21422 21416 21428
rect 21270 21383 21326 21392
rect 21284 21078 21312 21383
rect 21468 21321 21496 21490
rect 21548 21344 21600 21350
rect 21454 21312 21510 21321
rect 21548 21286 21600 21292
rect 21454 21247 21510 21256
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21272 21072 21324 21078
rect 21272 21014 21324 21020
rect 21376 20942 21404 21082
rect 21364 20936 21416 20942
rect 21270 20904 21326 20913
rect 21364 20878 21416 20884
rect 21270 20839 21326 20848
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21284 20398 21312 20839
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21100 19417 21128 20334
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 21086 19408 21142 19417
rect 21086 19343 21088 19352
rect 21140 19343 21142 19352
rect 21088 19314 21140 19320
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20548 18290 20576 18362
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20640 18170 20668 18770
rect 20824 18698 20852 19110
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20824 18290 20852 18634
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20548 18142 20668 18170
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20548 17921 20576 18142
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20534 17912 20590 17921
rect 20534 17847 20590 17856
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20444 14272 20496 14278
rect 20442 14240 20444 14249
rect 20496 14240 20498 14249
rect 20442 14175 20498 14184
rect 20442 14104 20498 14113
rect 20352 14068 20404 14074
rect 20442 14039 20498 14048
rect 20352 14010 20404 14016
rect 20258 13560 20314 13569
rect 20258 13495 20314 13504
rect 20258 13152 20314 13161
rect 20258 13087 20314 13096
rect 20272 12918 20300 13087
rect 20456 13002 20484 14039
rect 20364 12974 20484 13002
rect 20260 12912 20312 12918
rect 20166 12880 20222 12889
rect 20260 12854 20312 12860
rect 20166 12815 20222 12824
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 20180 11082 20208 12242
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20088 8090 20116 8434
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19720 6412 19840 6440
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19628 4826 19656 6258
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19720 3738 19748 6258
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19430 2952 19486 2961
rect 19430 2887 19486 2896
rect 19812 2774 19840 6412
rect 19892 6248 19944 6254
rect 19984 6248 20036 6254
rect 19892 6190 19944 6196
rect 19982 6216 19984 6225
rect 20036 6216 20038 6225
rect 19904 5234 19932 6190
rect 19982 6151 20038 6160
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19996 4146 20024 6054
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19996 3466 20024 4082
rect 20088 3670 20116 4082
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19812 2746 19932 2774
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 19614 2544 19670 2553
rect 19340 2508 19392 2514
rect 19614 2479 19670 2488
rect 19340 2450 19392 2456
rect 19352 2310 19380 2450
rect 19628 2446 19656 2479
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 19444 2038 19472 2246
rect 19536 2038 19564 2382
rect 19432 2032 19484 2038
rect 19432 1974 19484 1980
rect 19524 2032 19576 2038
rect 19524 1974 19576 1980
rect 17316 1964 17368 1970
rect 17316 1906 17368 1912
rect 19904 1902 19932 2746
rect 13728 1896 13780 1902
rect 13728 1838 13780 1844
rect 19892 1896 19944 1902
rect 19892 1838 19944 1844
rect 11612 1828 11664 1834
rect 11612 1770 11664 1776
rect 20180 800 20208 9658
rect 20272 2310 20300 12582
rect 20364 12345 20392 12974
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20548 12866 20576 17002
rect 20640 12986 20668 18022
rect 20732 17762 20760 18158
rect 20732 17734 20852 17762
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17202 20760 17614
rect 20824 17338 20852 17734
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20718 16824 20774 16833
rect 20718 16759 20774 16768
rect 20732 14929 20760 16759
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20824 16114 20852 16186
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20916 15706 20944 19246
rect 21100 18850 21128 19314
rect 21192 19009 21220 19722
rect 21178 19000 21234 19009
rect 21178 18935 21234 18944
rect 21100 18822 21220 18850
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 21100 18193 21128 18226
rect 21086 18184 21142 18193
rect 21086 18119 21142 18128
rect 20994 17640 21050 17649
rect 20994 17575 20996 17584
rect 21048 17575 21050 17584
rect 20996 17546 21048 17552
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20718 14920 20774 14929
rect 20718 14855 20774 14864
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14482 20760 14758
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13190 20760 13874
rect 20824 13705 20852 15438
rect 21008 15434 21036 16390
rect 21192 16250 21220 18822
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20810 13696 20866 13705
rect 20810 13631 20866 13640
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20350 12336 20406 12345
rect 20350 12271 20406 12280
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20364 6866 20392 11630
rect 20456 10674 20484 12854
rect 20548 12838 20668 12866
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20548 11354 20576 12650
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20640 11150 20668 12838
rect 20732 12170 20760 13126
rect 20916 12764 20944 13738
rect 21008 12918 21036 15370
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20916 12736 21036 12764
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20732 11762 20760 12106
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20534 10976 20590 10985
rect 20534 10911 20590 10920
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20456 9722 20484 9998
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 7886 20484 9318
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20456 7410 20484 7822
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20456 4622 20484 4966
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20548 3738 20576 10911
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20732 10062 20760 10474
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20640 9382 20668 9590
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20732 7954 20760 9998
rect 20824 9586 20852 12582
rect 21008 12220 21036 12736
rect 20916 12192 21036 12220
rect 20916 11762 20944 12192
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20904 11620 20956 11626
rect 20904 11562 20956 11568
rect 20916 10130 20944 11562
rect 21100 11558 21128 15982
rect 21192 13802 21220 15982
rect 21284 15570 21312 20198
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21376 14006 21404 19450
rect 21468 19446 21496 19654
rect 21456 19440 21508 19446
rect 21456 19382 21508 19388
rect 21468 18630 21496 19382
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21468 17610 21496 18566
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21468 17270 21496 17546
rect 21456 17264 21508 17270
rect 21456 17206 21508 17212
rect 21468 17134 21496 17206
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16250 21496 16934
rect 21560 16726 21588 21286
rect 21652 21078 21680 21558
rect 21744 21418 21772 22510
rect 21836 22094 21864 24375
rect 22204 23730 22232 24550
rect 22466 24511 22522 24520
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22388 23866 22416 24006
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22480 23798 22508 24511
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22572 24154 22600 24210
rect 22572 24126 22692 24154
rect 22468 23792 22520 23798
rect 22468 23734 22520 23740
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22664 23662 22692 24126
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21928 22273 21956 22986
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22296 22642 22324 22918
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 21914 22264 21970 22273
rect 21914 22199 21970 22208
rect 22190 22128 22246 22137
rect 21836 22066 21956 22094
rect 21732 21412 21784 21418
rect 21732 21354 21784 21360
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21640 21072 21692 21078
rect 21640 21014 21692 21020
rect 21652 20806 21680 21014
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21732 20800 21784 20806
rect 21732 20742 21784 20748
rect 21744 20641 21772 20742
rect 21730 20632 21786 20641
rect 21730 20567 21786 20576
rect 21732 20528 21784 20534
rect 21732 20470 21784 20476
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21652 19174 21680 19314
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21652 17746 21680 18838
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21468 15570 21496 15642
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21454 15192 21510 15201
rect 21454 15127 21510 15136
rect 21468 15094 21496 15127
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21560 14822 21588 14962
rect 21548 14816 21600 14822
rect 21546 14784 21548 14793
rect 21600 14784 21602 14793
rect 21546 14719 21602 14728
rect 21456 14544 21508 14550
rect 21456 14486 21508 14492
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21192 12986 21220 13398
rect 21284 13161 21312 13806
rect 21364 13728 21416 13734
rect 21362 13696 21364 13705
rect 21416 13696 21418 13705
rect 21362 13631 21418 13640
rect 21376 13462 21404 13631
rect 21364 13456 21416 13462
rect 21364 13398 21416 13404
rect 21468 13274 21496 14486
rect 21652 14464 21680 17682
rect 21744 16454 21772 20470
rect 21836 20244 21864 21354
rect 21928 20398 21956 22066
rect 22190 22063 22246 22072
rect 22204 22030 22232 22063
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 22020 21690 22048 21898
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21836 20216 21956 20244
rect 21824 20052 21876 20058
rect 21824 19994 21876 20000
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21732 16244 21784 16250
rect 21732 16186 21784 16192
rect 21376 13246 21496 13274
rect 21560 14436 21680 14464
rect 21270 13152 21326 13161
rect 21270 13087 21326 13096
rect 21376 13002 21404 13246
rect 21456 13184 21508 13190
rect 21454 13152 21456 13161
rect 21508 13152 21510 13161
rect 21454 13087 21510 13096
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21284 12974 21404 13002
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21192 12442 21220 12718
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21284 12322 21312 12974
rect 21362 12880 21418 12889
rect 21362 12815 21418 12824
rect 21192 12294 21312 12322
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20824 7834 20852 9318
rect 21008 8634 21036 11018
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20640 7806 20852 7834
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20456 3194 20484 3334
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20640 2774 20668 7806
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20732 6798 20760 7142
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20810 6352 20866 6361
rect 20810 6287 20812 6296
rect 20864 6287 20866 6296
rect 20812 6258 20864 6264
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 20916 5370 20944 5646
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 21100 5234 21128 11494
rect 21192 11354 21220 12294
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21178 11112 21234 11121
rect 21178 11047 21234 11056
rect 21192 10810 21220 11047
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21192 10198 21220 10406
rect 21180 10192 21232 10198
rect 21180 10134 21232 10140
rect 21192 9722 21220 10134
rect 21284 10130 21312 12174
rect 21376 12084 21404 12815
rect 21468 12646 21496 13087
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21560 12345 21588 14436
rect 21744 14396 21772 16186
rect 21836 14657 21864 19994
rect 21928 18902 21956 20216
rect 21916 18896 21968 18902
rect 21916 18838 21968 18844
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21928 16046 21956 18566
rect 22020 18306 22048 20402
rect 22112 18442 22140 21490
rect 22204 20913 22232 21966
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21486 22324 21830
rect 22480 21729 22508 23598
rect 22664 23186 22692 23598
rect 22652 23180 22704 23186
rect 22652 23122 22704 23128
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22572 22574 22600 22714
rect 22664 22710 22692 23122
rect 22652 22704 22704 22710
rect 22652 22646 22704 22652
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22756 22409 22784 26302
rect 23018 26200 23074 26302
rect 23386 26200 23442 27000
rect 24490 26200 24546 27000
rect 24858 26200 24914 27000
rect 25226 26200 25282 27000
rect 25870 26752 25926 26761
rect 25870 26687 25926 26696
rect 25686 26480 25742 26489
rect 25686 26415 25742 26424
rect 23400 25650 23428 26200
rect 23308 25622 23428 25650
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23308 23089 23336 25622
rect 23386 25528 23442 25537
rect 23386 25463 23442 25472
rect 24216 25492 24268 25498
rect 23400 24857 23428 25463
rect 24216 25434 24268 25440
rect 24032 25220 24084 25226
rect 24032 25162 24084 25168
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23386 24848 23442 24857
rect 23386 24783 23442 24792
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23400 23118 23428 23734
rect 23388 23112 23440 23118
rect 23294 23080 23350 23089
rect 23440 23072 23520 23100
rect 23388 23054 23440 23060
rect 23294 23015 23350 23024
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23124 22438 23152 22714
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23112 22432 23164 22438
rect 22742 22400 22798 22409
rect 23112 22374 23164 22380
rect 22742 22335 22798 22344
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 22466 21720 22522 21729
rect 22376 21684 22428 21690
rect 22466 21655 22522 21664
rect 22834 21720 22890 21729
rect 22834 21655 22890 21664
rect 22376 21626 22428 21632
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22190 20904 22246 20913
rect 22190 20839 22246 20848
rect 22296 20806 22324 21082
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22190 20632 22246 20641
rect 22190 20567 22246 20576
rect 22204 19417 22232 20567
rect 22296 20058 22324 20742
rect 22388 20602 22416 21626
rect 22742 21584 22798 21593
rect 22742 21519 22798 21528
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22572 21049 22600 21422
rect 22558 21040 22614 21049
rect 22468 21004 22520 21010
rect 22558 20975 22614 20984
rect 22468 20946 22520 20952
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22190 19408 22246 19417
rect 22296 19378 22324 19994
rect 22388 19990 22416 20538
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 22480 19938 22508 20946
rect 22650 20904 22706 20913
rect 22650 20839 22706 20848
rect 22664 20806 22692 20839
rect 22560 20800 22612 20806
rect 22558 20768 22560 20777
rect 22652 20800 22704 20806
rect 22612 20768 22614 20777
rect 22652 20742 22704 20748
rect 22558 20703 22614 20712
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22480 19910 22600 19938
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22480 19553 22508 19790
rect 22466 19544 22522 19553
rect 22572 19514 22600 19910
rect 22466 19479 22522 19488
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22664 19394 22692 20334
rect 22190 19343 22246 19352
rect 22284 19372 22336 19378
rect 22204 18698 22232 19343
rect 22284 19314 22336 19320
rect 22388 19366 22692 19394
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22112 18414 22232 18442
rect 22020 18278 22140 18306
rect 22112 17814 22140 18278
rect 22204 17814 22232 18414
rect 22100 17808 22152 17814
rect 22100 17750 22152 17756
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 22112 17218 22140 17750
rect 22204 17626 22232 17750
rect 22204 17598 22324 17626
rect 22296 17542 22324 17598
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22112 17190 22232 17218
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 22112 16998 22140 17070
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22100 16992 22152 16998
rect 22204 16969 22232 17190
rect 22100 16934 22152 16940
rect 22190 16960 22246 16969
rect 22020 16590 22048 16934
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 22020 16289 22048 16526
rect 22112 16425 22140 16934
rect 22190 16895 22246 16904
rect 22192 16720 22244 16726
rect 22192 16662 22244 16668
rect 22204 16454 22232 16662
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22192 16448 22244 16454
rect 22098 16416 22154 16425
rect 22192 16390 22244 16396
rect 22098 16351 22154 16360
rect 22006 16280 22062 16289
rect 22006 16215 22062 16224
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 22098 16008 22154 16017
rect 22098 15943 22154 15952
rect 22008 15904 22060 15910
rect 21914 15872 21970 15881
rect 22008 15846 22060 15852
rect 21914 15807 21970 15816
rect 21928 14929 21956 15807
rect 22020 15745 22048 15846
rect 22006 15736 22062 15745
rect 22006 15671 22062 15680
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21914 14920 21970 14929
rect 21914 14855 21970 14864
rect 21822 14648 21878 14657
rect 21822 14583 21878 14592
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21652 14368 21772 14396
rect 21546 12336 21602 12345
rect 21546 12271 21602 12280
rect 21548 12096 21600 12102
rect 21376 12056 21548 12084
rect 21548 12038 21600 12044
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 21192 2990 21220 9386
rect 21376 5778 21404 11698
rect 21468 11286 21496 11834
rect 21456 11280 21508 11286
rect 21456 11222 21508 11228
rect 21468 11150 21496 11222
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21560 10538 21588 12038
rect 21652 11898 21680 14368
rect 21928 14278 21956 14554
rect 22020 14482 22048 15438
rect 22112 14618 22140 15943
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21732 13864 21784 13870
rect 21730 13832 21732 13841
rect 21784 13832 21786 13841
rect 21730 13767 21786 13776
rect 21730 13424 21786 13433
rect 21730 13359 21786 13368
rect 21744 12986 21772 13359
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21730 12880 21786 12889
rect 21730 12815 21732 12824
rect 21784 12815 21786 12824
rect 21732 12786 21784 12792
rect 21836 12646 21864 14010
rect 21916 14000 21968 14006
rect 21916 13942 21968 13948
rect 21928 13394 21956 13942
rect 22204 13682 22232 15438
rect 22296 15026 22324 16594
rect 22388 15706 22416 19366
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22480 17202 22508 18362
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22572 17082 22600 19246
rect 22664 18902 22692 19246
rect 22756 19145 22784 21519
rect 22848 20913 22876 21655
rect 23032 21486 23060 21966
rect 23112 21956 23164 21962
rect 23112 21898 23164 21904
rect 23020 21480 23072 21486
rect 23020 21422 23072 21428
rect 23124 21418 23152 21898
rect 23308 21554 23336 22646
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22834 20904 22890 20913
rect 22834 20839 22890 20848
rect 22940 20244 22968 20946
rect 23110 20632 23166 20641
rect 23110 20567 23112 20576
rect 23164 20567 23166 20576
rect 23112 20538 23164 20544
rect 23308 20466 23336 21490
rect 23400 21434 23428 22918
rect 23492 22098 23520 23072
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23584 21622 23612 24890
rect 23940 24676 23992 24682
rect 23940 24618 23992 24624
rect 23952 24410 23980 24618
rect 23940 24404 23992 24410
rect 23940 24346 23992 24352
rect 23754 24304 23810 24313
rect 23754 24239 23810 24248
rect 23768 24206 23796 24239
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23768 21690 23796 24142
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23860 23202 23888 24006
rect 23860 23174 23980 23202
rect 23848 22976 23900 22982
rect 23848 22918 23900 22924
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23572 21480 23624 21486
rect 23400 21406 23520 21434
rect 23572 21422 23624 21428
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22848 20216 22968 20244
rect 22742 19136 22798 19145
rect 22742 19071 22798 19080
rect 22652 18896 22704 18902
rect 22652 18838 22704 18844
rect 22848 18850 22876 20216
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23112 19984 23164 19990
rect 23112 19926 23164 19932
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22940 19242 22968 19790
rect 23020 19712 23072 19718
rect 23018 19680 23020 19689
rect 23072 19680 23074 19689
rect 23018 19615 23074 19624
rect 23124 19378 23152 19926
rect 23216 19718 23244 19994
rect 23308 19922 23336 20402
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23308 19378 23336 19858
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23296 19372 23348 19378
rect 23400 19360 23428 21286
rect 23492 19990 23520 21406
rect 23584 21010 23612 21422
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23584 20777 23612 20946
rect 23664 20800 23716 20806
rect 23570 20768 23626 20777
rect 23664 20742 23716 20748
rect 23570 20703 23626 20712
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23480 19984 23532 19990
rect 23480 19926 23532 19932
rect 23400 19332 23520 19360
rect 23296 19314 23348 19320
rect 22928 19236 22980 19242
rect 22928 19178 22980 19184
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22848 18822 22968 18850
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22480 17054 22600 17082
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22480 15502 22508 17054
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22296 14618 22324 14962
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22296 13938 22324 14554
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22388 13841 22416 15030
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 22374 13832 22430 13841
rect 22374 13767 22430 13776
rect 22204 13654 22324 13682
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21928 12850 21956 13330
rect 22006 13152 22062 13161
rect 22006 13087 22062 13096
rect 22020 12889 22048 13087
rect 22006 12880 22062 12889
rect 21916 12844 21968 12850
rect 22006 12815 22062 12824
rect 21916 12786 21968 12792
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21822 12336 21878 12345
rect 21822 12271 21878 12280
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 5846 21588 6598
rect 21652 6118 21680 11698
rect 21730 11520 21786 11529
rect 21730 11455 21786 11464
rect 21744 10810 21772 11455
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 21732 10600 21784 10606
rect 21732 10542 21784 10548
rect 21744 9926 21772 10542
rect 21836 10470 21864 12271
rect 21928 12238 21956 12786
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22190 12608 22246 12617
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21836 9994 21864 10406
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21548 5840 21600 5846
rect 21548 5782 21600 5788
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 21836 3058 21864 8774
rect 21928 3534 21956 11086
rect 22020 8430 22048 12582
rect 22112 12442 22140 12582
rect 22190 12543 22246 12552
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22112 10538 22140 12378
rect 22100 10532 22152 10538
rect 22100 10474 22152 10480
rect 22204 9738 22232 12543
rect 22112 9710 22232 9738
rect 22112 9178 22140 9710
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22098 9072 22154 9081
rect 22098 9007 22154 9016
rect 22112 8498 22140 9007
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 22204 8022 22232 9522
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 22020 6458 22048 6870
rect 22204 6866 22232 7686
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 22296 6798 22324 13654
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22388 12646 22416 12922
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22388 6458 22416 7822
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22480 4622 22508 14826
rect 22572 11354 22600 16118
rect 22664 15178 22692 18566
rect 22756 18329 22784 18702
rect 22742 18320 22798 18329
rect 22742 18255 22798 18264
rect 22848 17814 22876 18702
rect 22940 18086 22968 18822
rect 23308 18426 23336 19314
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 22928 18080 22980 18086
rect 22928 18022 22980 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17808 22888 17814
rect 22836 17750 22888 17756
rect 22848 17649 22876 17750
rect 22834 17640 22890 17649
rect 22834 17575 22890 17584
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22756 16114 22784 16390
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22664 15150 22784 15178
rect 22650 15056 22706 15065
rect 22650 14991 22706 15000
rect 22664 14958 22692 14991
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22756 14890 22784 15150
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22848 14770 22876 17070
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23216 16697 23244 16730
rect 23202 16688 23258 16697
rect 23202 16623 23258 16632
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23032 14822 23060 15642
rect 22664 14742 22876 14770
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 22664 12753 22692 14742
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22742 13968 22798 13977
rect 22742 13903 22798 13912
rect 22650 12744 22706 12753
rect 22650 12679 22706 12688
rect 22652 12640 22704 12646
rect 22650 12608 22652 12617
rect 22704 12608 22706 12617
rect 22650 12543 22706 12552
rect 22756 12434 22784 13903
rect 22848 12986 22876 14350
rect 23020 14272 23072 14278
rect 23020 14214 23072 14220
rect 23032 14113 23060 14214
rect 23018 14104 23074 14113
rect 23018 14039 23074 14048
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22926 13424 22982 13433
rect 22926 13359 22982 13368
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22940 12918 22968 13359
rect 23018 13288 23074 13297
rect 23018 13223 23074 13232
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 23032 12730 23060 13223
rect 22664 12406 22784 12434
rect 22848 12702 23060 12730
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22664 11234 22692 12406
rect 22848 12306 22876 12702
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22572 11206 22692 11234
rect 22572 6866 22600 11206
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22664 9625 22692 11086
rect 22650 9616 22706 9625
rect 22650 9551 22706 9560
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 22664 6746 22692 9454
rect 22756 7274 22784 11698
rect 22848 7970 22876 12242
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 9518 22968 9862
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22848 7942 22968 7970
rect 22836 7880 22888 7886
rect 22834 7848 22836 7857
rect 22888 7848 22890 7857
rect 22834 7783 22890 7792
rect 22940 7698 22968 7942
rect 22848 7670 22968 7698
rect 22744 7268 22796 7274
rect 22744 7210 22796 7216
rect 22572 6718 22692 6746
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20548 2746 20668 2774
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 20548 1834 20576 2746
rect 20732 2378 20760 2790
rect 22112 2650 22140 2994
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 22204 2009 22232 3062
rect 22190 2000 22246 2009
rect 22190 1935 22246 1944
rect 20536 1828 20588 1834
rect 20536 1770 20588 1776
rect 22296 1601 22324 4014
rect 22572 2854 22600 6718
rect 22848 6118 22876 7670
rect 23308 7426 23336 17478
rect 23400 15994 23428 18838
rect 23492 16250 23520 19332
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23400 15966 23520 15994
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23400 15337 23428 15846
rect 23386 15328 23442 15337
rect 23386 15263 23442 15272
rect 23388 14952 23440 14958
rect 23388 14894 23440 14900
rect 23400 14482 23428 14894
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 13025 23428 14214
rect 23492 13530 23520 15966
rect 23584 15201 23612 20198
rect 23676 18970 23704 20742
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23768 19961 23796 20334
rect 23754 19952 23810 19961
rect 23754 19887 23810 19896
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23768 19417 23796 19654
rect 23754 19408 23810 19417
rect 23754 19343 23810 19352
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23860 17610 23888 22918
rect 23952 22710 23980 23174
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23952 21690 23980 22646
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 23848 17604 23900 17610
rect 23848 17546 23900 17552
rect 23952 17354 23980 19246
rect 24044 18873 24072 25162
rect 24228 22094 24256 25434
rect 24306 25256 24362 25265
rect 24306 25191 24362 25200
rect 24320 23322 24348 25191
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24308 23316 24360 23322
rect 24308 23258 24360 23264
rect 24228 22066 24348 22094
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24228 20534 24256 21626
rect 24216 20528 24268 20534
rect 24216 20470 24268 20476
rect 24320 19417 24348 22066
rect 24412 19922 24440 23462
rect 24504 22234 24532 26200
rect 24950 26072 25006 26081
rect 24950 26007 25006 26016
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24492 22228 24544 22234
rect 24492 22170 24544 22176
rect 24596 22094 24624 22918
rect 24504 22066 24624 22094
rect 24400 19916 24452 19922
rect 24400 19858 24452 19864
rect 24306 19408 24362 19417
rect 24306 19343 24362 19352
rect 24030 18864 24086 18873
rect 24030 18799 24086 18808
rect 24412 18465 24440 19858
rect 24398 18456 24454 18465
rect 24398 18391 24454 18400
rect 24400 18080 24452 18086
rect 24400 18022 24452 18028
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 23768 17326 23980 17354
rect 23662 16824 23718 16833
rect 23662 16759 23718 16768
rect 23676 16726 23704 16759
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23570 15192 23626 15201
rect 23570 15127 23626 15136
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23584 14006 23612 15030
rect 23676 14521 23704 15914
rect 23662 14512 23718 14521
rect 23662 14447 23718 14456
rect 23572 14000 23624 14006
rect 23624 13960 23704 13988
rect 23572 13942 23624 13948
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23386 13016 23442 13025
rect 23386 12951 23442 12960
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23492 11626 23520 12922
rect 23584 12050 23612 13330
rect 23676 13258 23704 13960
rect 23768 13870 23796 17326
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23860 16522 23888 17138
rect 24044 17134 24072 17682
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23952 15638 23980 16526
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 24044 16046 24072 16390
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23940 15632 23992 15638
rect 23940 15574 23992 15580
rect 24136 15366 24164 16050
rect 24228 15502 24256 16390
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 24136 15201 24164 15302
rect 24122 15192 24178 15201
rect 24122 15127 24178 15136
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 24044 14074 24072 14418
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23676 12918 23704 13194
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 23676 12170 23704 12854
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 23584 12022 23704 12050
rect 23570 11928 23626 11937
rect 23570 11863 23626 11872
rect 23480 11620 23532 11626
rect 23480 11562 23532 11568
rect 23480 9988 23532 9994
rect 23480 9930 23532 9936
rect 23492 9738 23520 9930
rect 23400 9710 23520 9738
rect 23400 9382 23428 9710
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23400 8129 23428 8366
rect 23386 8120 23442 8129
rect 23386 8055 23442 8064
rect 23308 7398 23428 7426
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23308 6905 23336 7278
rect 23294 6896 23350 6905
rect 23294 6831 23350 6840
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22848 5302 22876 6054
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22836 5296 22888 5302
rect 22836 5238 22888 5244
rect 23400 5166 23428 7398
rect 23480 6384 23532 6390
rect 23480 6326 23532 6332
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22664 3534 22692 4422
rect 23400 4049 23428 4490
rect 23492 4146 23520 6326
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23386 4040 23442 4049
rect 23386 3975 23442 3984
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 23388 3460 23440 3466
rect 23388 3402 23440 3408
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22664 2106 22692 2382
rect 22652 2100 22704 2106
rect 22652 2042 22704 2048
rect 22282 1592 22338 1601
rect 22282 1527 22338 1536
rect 23400 1193 23428 3402
rect 23584 2774 23612 11863
rect 23676 10792 23704 12022
rect 23860 10996 23888 13874
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 23952 12102 23980 13466
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23938 11792 23994 11801
rect 23938 11727 23940 11736
rect 23992 11727 23994 11736
rect 23940 11698 23992 11704
rect 24044 11121 24072 12786
rect 24136 12442 24164 14214
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24124 12232 24176 12238
rect 24122 12200 24124 12209
rect 24176 12200 24178 12209
rect 24122 12135 24178 12144
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 24030 11112 24086 11121
rect 24030 11047 24086 11056
rect 23860 10968 23980 10996
rect 23676 10764 23796 10792
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23676 7954 23704 10610
rect 23768 10010 23796 10764
rect 23952 10656 23980 10968
rect 23860 10628 23980 10656
rect 23860 10266 23888 10628
rect 24136 10588 24164 12038
rect 24228 11014 24256 14010
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 23952 10560 24164 10588
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23768 9982 23888 10010
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23768 4690 23796 9862
rect 23860 7546 23888 9982
rect 23952 8650 23980 10560
rect 24214 10432 24270 10441
rect 24214 10367 24270 10376
rect 24228 10266 24256 10367
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24124 10192 24176 10198
rect 24228 10169 24256 10202
rect 24124 10134 24176 10140
rect 24214 10160 24270 10169
rect 23952 8622 24072 8650
rect 23938 8528 23994 8537
rect 23938 8463 23940 8472
rect 23992 8463 23994 8472
rect 23940 8434 23992 8440
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23938 7440 23994 7449
rect 23938 7375 23940 7384
rect 23992 7375 23994 7384
rect 23940 7346 23992 7352
rect 23938 6624 23994 6633
rect 23938 6559 23994 6568
rect 23952 6322 23980 6559
rect 24044 6390 24072 8622
rect 24032 6384 24084 6390
rect 24032 6326 24084 6332
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 23952 5234 23980 6122
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23492 2746 23612 2774
rect 23492 2582 23520 2746
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 24136 2038 24164 10134
rect 24214 10095 24270 10104
rect 24320 10010 24348 15982
rect 24412 14958 24440 18022
rect 24504 17678 24532 22066
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24596 20942 24624 21830
rect 24676 21072 24728 21078
rect 24674 21040 24676 21049
rect 24728 21040 24730 21049
rect 24674 20975 24730 20984
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24582 19816 24638 19825
rect 24582 19751 24638 19760
rect 24596 19718 24624 19751
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24780 19310 24808 25366
rect 24964 23118 24992 26007
rect 25134 25664 25190 25673
rect 25134 25599 25190 25608
rect 25044 24336 25096 24342
rect 25044 24278 25096 24284
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 24860 22568 24912 22574
rect 24858 22536 24860 22545
rect 24912 22536 24914 22545
rect 24858 22471 24914 22480
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 24676 18692 24728 18698
rect 24676 18634 24728 18640
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18057 24624 18566
rect 24582 18048 24638 18057
rect 24582 17983 24638 17992
rect 24492 17672 24544 17678
rect 24492 17614 24544 17620
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24596 15706 24624 16050
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24228 9982 24348 10010
rect 24228 8362 24256 9982
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24320 7993 24348 9862
rect 24306 7984 24362 7993
rect 24306 7919 24362 7928
rect 24412 7886 24440 14894
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24504 12986 24532 14282
rect 24596 13190 24624 14758
rect 24688 13530 24716 18634
rect 24766 18184 24822 18193
rect 24766 18119 24768 18128
rect 24820 18119 24822 18128
rect 24768 18090 24820 18096
rect 24780 17202 24808 18090
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24780 14929 24808 16594
rect 24766 14920 24822 14929
rect 24766 14855 24822 14864
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 24780 13258 24808 14214
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 24584 13184 24636 13190
rect 24584 13126 24636 13132
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24674 12608 24730 12617
rect 24674 12543 24730 12552
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24504 3398 24532 12378
rect 24688 12306 24716 12543
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24674 12064 24730 12073
rect 24596 11150 24624 12038
rect 24674 11999 24730 12008
rect 24688 11762 24716 11999
rect 24872 11914 24900 21830
rect 24964 21078 24992 22714
rect 24952 21072 25004 21078
rect 24952 21014 25004 21020
rect 25056 18834 25084 24278
rect 25148 24206 25176 25599
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 25228 23588 25280 23594
rect 25228 23530 25280 23536
rect 25240 23497 25268 23530
rect 25226 23488 25282 23497
rect 25226 23423 25282 23432
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25148 20346 25176 23122
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25240 21146 25268 23054
rect 25332 21350 25360 24210
rect 25412 23724 25464 23730
rect 25412 23666 25464 23672
rect 25424 23633 25452 23666
rect 25410 23624 25466 23633
rect 25410 23559 25466 23568
rect 25516 22166 25544 24346
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25410 21448 25466 21457
rect 25608 21418 25636 24006
rect 25700 22030 25728 26415
rect 25778 22400 25834 22409
rect 25778 22335 25834 22344
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25410 21383 25466 21392
rect 25596 21412 25648 21418
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25424 21162 25452 21383
rect 25596 21354 25648 21360
rect 25504 21344 25556 21350
rect 25700 21298 25728 21966
rect 25504 21286 25556 21292
rect 25228 21140 25280 21146
rect 25228 21082 25280 21088
rect 25332 21134 25452 21162
rect 25332 20534 25360 21134
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25148 20318 25268 20346
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25148 18834 25176 20198
rect 25240 19514 25268 20318
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 25332 19417 25360 19654
rect 25318 19408 25374 19417
rect 25318 19343 25374 19352
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25148 18737 25176 18770
rect 25134 18728 25190 18737
rect 25134 18663 25190 18672
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24964 18057 24992 18566
rect 24950 18048 25006 18057
rect 24950 17983 25006 17992
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 13326 24992 17478
rect 25240 17105 25268 19246
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25332 18358 25360 18702
rect 25320 18352 25372 18358
rect 25320 18294 25372 18300
rect 25226 17096 25282 17105
rect 25226 17031 25282 17040
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25240 15609 25268 15846
rect 25226 15600 25282 15609
rect 25226 15535 25282 15544
rect 25226 15328 25282 15337
rect 25226 15263 25282 15272
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24964 12238 24992 13126
rect 25056 12306 25084 14758
rect 25148 14074 25176 15098
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25240 13394 25268 15263
rect 25332 14346 25360 18294
rect 25424 14414 25452 20742
rect 25516 18601 25544 21286
rect 25608 21270 25728 21298
rect 25608 20641 25636 21270
rect 25686 21176 25742 21185
rect 25686 21111 25742 21120
rect 25594 20632 25650 20641
rect 25594 20567 25650 20576
rect 25596 20528 25648 20534
rect 25596 20470 25648 20476
rect 25502 18592 25558 18601
rect 25502 18527 25558 18536
rect 25608 18290 25636 20470
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25594 16824 25650 16833
rect 25594 16759 25650 16768
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 25320 14340 25372 14346
rect 25320 14282 25372 14288
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25226 13016 25282 13025
rect 25226 12951 25282 12960
rect 25134 12608 25190 12617
rect 25134 12543 25190 12552
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 25042 12200 25098 12209
rect 25042 12135 25098 12144
rect 24872 11886 24992 11914
rect 24860 11824 24912 11830
rect 24766 11792 24822 11801
rect 24676 11756 24728 11762
rect 24860 11766 24912 11772
rect 24766 11727 24822 11736
rect 24676 11698 24728 11704
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24674 9616 24730 9625
rect 24674 9551 24730 9560
rect 24688 7410 24716 9551
rect 24780 9518 24808 11727
rect 24872 11393 24900 11766
rect 24964 11694 24992 11886
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 25056 11218 25084 12135
rect 25148 11830 25176 12543
rect 25240 11898 25268 12951
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25332 12442 25360 12582
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 25134 10976 25190 10985
rect 25134 10911 25190 10920
rect 25148 10742 25176 10911
rect 25136 10736 25188 10742
rect 25136 10678 25188 10684
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 25134 10568 25190 10577
rect 24872 10169 24900 10542
rect 25134 10503 25190 10512
rect 25042 10296 25098 10305
rect 25042 10231 25098 10240
rect 24858 10160 24914 10169
rect 25056 10130 25084 10231
rect 24858 10095 24914 10104
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24872 9353 24900 9590
rect 24858 9344 24914 9353
rect 24858 9279 24914 9288
rect 24950 8936 25006 8945
rect 24950 8871 24952 8880
rect 25004 8871 25006 8880
rect 24952 8842 25004 8848
rect 25148 8566 25176 10503
rect 25240 8974 25268 11018
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25136 8560 25188 8566
rect 24766 8528 24822 8537
rect 25136 8502 25188 8508
rect 24766 8463 24822 8472
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24674 7304 24730 7313
rect 24674 7239 24730 7248
rect 24582 5264 24638 5273
rect 24582 5199 24638 5208
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24596 2990 24624 5199
rect 24688 5166 24716 7239
rect 24780 6254 24808 8463
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24964 7721 24992 7754
rect 25228 7744 25280 7750
rect 24950 7712 25006 7721
rect 25228 7686 25280 7692
rect 24950 7647 25006 7656
rect 25240 6798 25268 7686
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24766 6080 24822 6089
rect 24766 6015 24822 6024
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24780 4078 24808 6015
rect 24950 5672 25006 5681
rect 24950 5607 24952 5616
rect 25004 5607 25006 5616
rect 24952 5578 25004 5584
rect 24860 5296 24912 5302
rect 24860 5238 24912 5244
rect 24872 4865 24900 5238
rect 24858 4856 24914 4865
rect 24858 4791 24914 4800
rect 25056 4622 25084 6598
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 25044 4616 25096 4622
rect 25044 4558 25096 4564
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24964 4457 24992 4490
rect 24950 4448 25006 4457
rect 24950 4383 25006 4392
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24952 4004 25004 4010
rect 24952 3946 25004 3952
rect 24964 3641 24992 3946
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 24584 2984 24636 2990
rect 24584 2926 24636 2932
rect 24872 2825 24900 3062
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 24858 2816 24914 2825
rect 24858 2751 24914 2760
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24124 2032 24176 2038
rect 24124 1974 24176 1980
rect 24596 1970 24624 2382
rect 24584 1964 24636 1970
rect 24584 1906 24636 1912
rect 23386 1184 23442 1193
rect 23386 1119 23442 1128
rect 6734 0 6790 800
rect 20166 0 20222 800
rect 24872 377 24900 2450
rect 24950 2408 25006 2417
rect 24950 2343 24952 2352
rect 25004 2343 25006 2352
rect 24952 2314 25004 2320
rect 25056 785 25084 2858
rect 25148 2650 25176 3538
rect 25240 3534 25268 5510
rect 25332 5370 25360 12242
rect 25320 5364 25372 5370
rect 25320 5306 25372 5312
rect 25424 4826 25452 13670
rect 25516 11150 25544 15302
rect 25608 15178 25636 16759
rect 25700 16658 25728 21111
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25688 16176 25740 16182
rect 25688 16118 25740 16124
rect 25700 15314 25728 16118
rect 25792 15745 25820 22335
rect 25884 18426 25912 26687
rect 26054 23624 26110 23633
rect 26110 23582 26280 23610
rect 26054 23559 26110 23568
rect 25962 23216 26018 23225
rect 25962 23151 26018 23160
rect 25976 21570 26004 23151
rect 26054 22808 26110 22817
rect 26054 22743 26110 22752
rect 26068 22438 26096 22743
rect 26056 22432 26108 22438
rect 26056 22374 26108 22380
rect 25976 21542 26188 21570
rect 26056 21412 26108 21418
rect 26056 21354 26108 21360
rect 25962 19952 26018 19961
rect 25962 19887 26018 19896
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 25778 15736 25834 15745
rect 25778 15671 25834 15680
rect 25778 15464 25834 15473
rect 25778 15399 25780 15408
rect 25832 15399 25834 15408
rect 25780 15370 25832 15376
rect 25700 15286 25820 15314
rect 25608 15150 25728 15178
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25608 13870 25636 14962
rect 25596 13864 25648 13870
rect 25594 13832 25596 13841
rect 25648 13832 25650 13841
rect 25594 13767 25650 13776
rect 25596 13252 25648 13258
rect 25596 13194 25648 13200
rect 25608 12374 25636 13194
rect 25596 12368 25648 12374
rect 25596 12310 25648 12316
rect 25596 12164 25648 12170
rect 25596 12106 25648 12112
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25608 8838 25636 12106
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25700 6916 25728 15150
rect 25792 9178 25820 15286
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25884 7478 25912 18226
rect 25976 12646 26004 19887
rect 26068 14385 26096 21354
rect 26160 15586 26188 21542
rect 26252 17270 26280 23582
rect 26884 23044 26936 23050
rect 26884 22986 26936 22992
rect 26700 22432 26752 22438
rect 26700 22374 26752 22380
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26240 17264 26292 17270
rect 26240 17206 26292 17212
rect 26160 15558 26280 15586
rect 26054 14376 26110 14385
rect 26054 14311 26110 14320
rect 26054 14240 26110 14249
rect 26054 14175 26110 14184
rect 25964 12640 26016 12646
rect 25964 12582 26016 12588
rect 26068 12152 26096 14175
rect 26252 13546 26280 15558
rect 26424 15428 26476 15434
rect 26424 15370 26476 15376
rect 26160 13518 26280 13546
rect 26160 12782 26188 13518
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26148 12640 26200 12646
rect 26148 12582 26200 12588
rect 25976 12124 26096 12152
rect 25976 11948 26004 12124
rect 25976 11920 26096 11948
rect 25872 7472 25924 7478
rect 25872 7414 25924 7420
rect 25608 6888 25728 6916
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25608 3738 25636 6888
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 25700 6497 25728 6666
rect 25686 6488 25742 6497
rect 25686 6423 25742 6432
rect 26068 5098 26096 11920
rect 26056 5092 26108 5098
rect 26056 5034 26108 5040
rect 26160 4758 26188 12582
rect 26252 7954 26280 13398
rect 26332 12028 26384 12034
rect 26332 11970 26384 11976
rect 26240 7948 26292 7954
rect 26240 7890 26292 7896
rect 26148 4752 26200 4758
rect 26148 4694 26200 4700
rect 26344 4282 26372 11970
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 26436 4214 26464 15370
rect 26528 10810 26556 19450
rect 26608 18896 26660 18902
rect 26608 18838 26660 18844
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26424 4208 26476 4214
rect 26424 4150 26476 4156
rect 25596 3732 25648 3738
rect 25596 3674 25648 3680
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25688 3460 25740 3466
rect 25688 3402 25740 3408
rect 25700 3233 25728 3402
rect 25686 3224 25742 3233
rect 25686 3159 25742 3168
rect 26620 3058 26648 18838
rect 26712 11762 26740 22374
rect 26792 17264 26844 17270
rect 26792 17206 26844 17212
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26804 7002 26832 17206
rect 26896 13530 26924 22986
rect 26884 13524 26936 13530
rect 26884 13466 26936 13472
rect 26792 6996 26844 7002
rect 26792 6938 26844 6944
rect 26608 3052 26660 3058
rect 26608 2994 26660 3000
rect 25136 2644 25188 2650
rect 25136 2586 25188 2592
rect 25042 776 25098 785
rect 25042 711 25098 720
rect 24858 368 24914 377
rect 24858 303 24914 312
<< via2 >>
rect 1214 26832 1270 26888
rect 938 25744 994 25800
rect 478 25064 534 25120
rect 478 15272 534 15328
rect 938 25064 994 25120
rect 662 24248 718 24304
rect 938 20984 994 21040
rect 1766 24012 1768 24032
rect 1768 24012 1820 24032
rect 1820 24012 1822 24032
rect 1766 23976 1822 24012
rect 1214 15408 1270 15464
rect 1950 23024 2006 23080
rect 1858 22072 1914 22128
rect 1398 15272 1454 15328
rect 1582 9172 1638 9208
rect 1582 9152 1584 9172
rect 1584 9152 1636 9172
rect 1636 9152 1638 9172
rect 2226 23160 2282 23216
rect 2134 21664 2190 21720
rect 2226 20884 2228 20904
rect 2228 20884 2280 20904
rect 2280 20884 2282 20904
rect 2226 20848 2282 20884
rect 2594 23976 2650 24032
rect 2502 21392 2558 21448
rect 2778 23704 2834 23760
rect 2686 22480 2742 22536
rect 1858 11620 1914 11656
rect 1858 11600 1860 11620
rect 1860 11600 1912 11620
rect 1912 11600 1914 11620
rect 1858 11348 1914 11384
rect 1858 11328 1860 11348
rect 1860 11328 1912 11348
rect 1912 11328 1914 11348
rect 2042 11192 2098 11248
rect 3238 25880 3294 25936
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2962 23724 3018 23760
rect 2962 23704 2964 23724
rect 2964 23704 3016 23724
rect 3016 23704 3018 23724
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3422 22616 3478 22672
rect 3698 24792 3754 24848
rect 3974 24284 3976 24304
rect 3976 24284 4028 24304
rect 4028 24284 4030 24304
rect 3974 24248 4030 24284
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2594 15000 2650 15056
rect 2594 12144 2650 12200
rect 2410 11076 2466 11112
rect 2410 11056 2412 11076
rect 2412 11056 2464 11076
rect 2464 11056 2466 11076
rect 2318 9424 2374 9480
rect 1766 6296 1822 6352
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 3422 17604 3478 17640
rect 3422 17584 3424 17604
rect 3424 17584 3476 17604
rect 3476 17584 3478 17604
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2870 16632 2926 16688
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3238 13232 3294 13288
rect 2870 12824 2926 12880
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2778 9988 2834 10024
rect 2778 9968 2780 9988
rect 2780 9968 2832 9988
rect 2832 9968 2834 9988
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3698 22208 3754 22264
rect 4894 26560 4950 26616
rect 3882 21664 3938 21720
rect 4342 21936 4398 21992
rect 4066 19352 4122 19408
rect 4066 18944 4122 19000
rect 3974 17756 3976 17776
rect 3976 17756 4028 17776
rect 4028 17756 4030 17776
rect 3974 17720 4030 17756
rect 4158 18808 4214 18864
rect 3790 14728 3846 14784
rect 3514 12280 3570 12336
rect 3422 11192 3478 11248
rect 2594 8628 2650 8664
rect 2594 8608 2596 8628
rect 2596 8608 2648 8628
rect 2648 8608 2650 8628
rect 3238 8744 3294 8800
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2594 7964 2596 7984
rect 2596 7964 2648 7984
rect 2648 7964 2650 7984
rect 2594 7928 2650 7964
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3790 11464 3846 11520
rect 3974 15816 4030 15872
rect 3974 14320 4030 14376
rect 4802 23296 4858 23352
rect 4710 22072 4766 22128
rect 4618 21936 4674 21992
rect 4710 20596 4766 20632
rect 4710 20576 4712 20596
rect 4712 20576 4764 20596
rect 4764 20576 4766 20596
rect 4434 15136 4490 15192
rect 4618 16496 4674 16552
rect 4710 14864 4766 14920
rect 4434 10920 4490 10976
rect 4342 10784 4398 10840
rect 4250 10512 4306 10568
rect 3790 10376 3846 10432
rect 3698 7248 3754 7304
rect 4158 9016 4214 9072
rect 4158 8492 4214 8528
rect 4158 8472 4160 8492
rect 4160 8472 4212 8492
rect 4212 8472 4214 8492
rect 5170 26424 5226 26480
rect 5170 21664 5226 21720
rect 4986 18672 5042 18728
rect 4710 12688 4766 12744
rect 4618 11464 4674 11520
rect 4710 9152 4766 9208
rect 5446 23432 5502 23488
rect 5814 19216 5870 19272
rect 5354 17196 5410 17232
rect 5354 17176 5356 17196
rect 5356 17176 5408 17196
rect 5408 17176 5410 17196
rect 5262 12416 5318 12472
rect 5170 11736 5226 11792
rect 5170 9596 5172 9616
rect 5172 9596 5224 9616
rect 5224 9596 5226 9616
rect 5170 9560 5226 9596
rect 5170 7928 5226 7984
rect 4986 7792 5042 7848
rect 4066 6704 4122 6760
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 6734 23568 6790 23624
rect 6182 18420 6238 18456
rect 6182 18400 6184 18420
rect 6184 18400 6236 18420
rect 6236 18400 6238 18420
rect 6734 23432 6790 23488
rect 6458 21392 6514 21448
rect 6642 21292 6644 21312
rect 6644 21292 6696 21312
rect 6696 21292 6698 21312
rect 6642 21256 6698 21292
rect 7286 23840 7342 23896
rect 7010 21120 7066 21176
rect 7010 20848 7066 20904
rect 6642 20304 6698 20360
rect 6366 18264 6422 18320
rect 5814 13504 5870 13560
rect 5814 12552 5870 12608
rect 6550 16088 6606 16144
rect 6182 11736 6238 11792
rect 6090 10240 6146 10296
rect 6366 14476 6422 14512
rect 6366 14456 6368 14476
rect 6368 14456 6420 14476
rect 6420 14456 6422 14476
rect 7746 25744 7802 25800
rect 7746 25336 7802 25392
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7286 20848 7342 20904
rect 7378 19760 7434 19816
rect 7286 17040 7342 17096
rect 7286 13368 7342 13424
rect 6918 12960 6974 13016
rect 6826 12844 6882 12880
rect 6826 12824 6828 12844
rect 6828 12824 6880 12844
rect 6880 12824 6882 12844
rect 6826 12688 6882 12744
rect 7010 12688 7066 12744
rect 6918 12416 6974 12472
rect 6918 11192 6974 11248
rect 7102 10804 7158 10840
rect 7102 10784 7104 10804
rect 7104 10784 7156 10804
rect 7156 10784 7158 10804
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8390 21664 8446 21720
rect 7654 20576 7710 20632
rect 7654 16632 7710 16688
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7838 20460 7894 20496
rect 7838 20440 7840 20460
rect 7840 20440 7892 20460
rect 7892 20440 7894 20460
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8666 22888 8722 22944
rect 8574 21256 8630 21312
rect 8574 21120 8630 21176
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7838 15408 7894 15464
rect 7562 12280 7618 12336
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 8298 13776 8354 13832
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7838 12280 7894 12336
rect 9034 22752 9090 22808
rect 9218 22616 9274 22672
rect 9494 22344 9550 22400
rect 10966 25336 11022 25392
rect 9954 23432 10010 23488
rect 9126 21936 9182 21992
rect 8758 20712 8814 20768
rect 9126 21528 9182 21584
rect 8850 20168 8906 20224
rect 8758 20032 8814 20088
rect 8574 19080 8630 19136
rect 8574 17856 8630 17912
rect 8482 17040 8538 17096
rect 8482 16768 8538 16824
rect 8666 17312 8722 17368
rect 9034 18536 9090 18592
rect 9218 21256 9274 21312
rect 9402 21120 9458 21176
rect 9218 19760 9274 19816
rect 9126 18128 9182 18184
rect 9402 19624 9458 19680
rect 9310 18400 9366 18456
rect 9954 22752 10010 22808
rect 9678 21004 9734 21040
rect 9678 20984 9680 21004
rect 9680 20984 9732 21004
rect 9732 20984 9734 21004
rect 9586 20576 9642 20632
rect 9586 20304 9642 20360
rect 9402 17856 9458 17912
rect 9586 18536 9642 18592
rect 9678 17856 9734 17912
rect 9126 17448 9182 17504
rect 9586 17312 9642 17368
rect 9954 20748 9956 20768
rect 9956 20748 10008 20768
rect 10008 20748 10010 20768
rect 9954 20712 10010 20748
rect 9954 18672 10010 18728
rect 9954 18264 10010 18320
rect 9862 17448 9918 17504
rect 9770 17312 9826 17368
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7746 9580 7802 9616
rect 7746 9560 7748 9580
rect 7748 9560 7800 9580
rect 7800 9560 7802 9580
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 8390 11348 8446 11384
rect 8390 11328 8392 11348
rect 8392 11328 8444 11348
rect 8444 11328 8446 11348
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 8666 16244 8722 16280
rect 8666 16224 8668 16244
rect 8668 16224 8720 16244
rect 8720 16224 8722 16244
rect 9402 16360 9458 16416
rect 8850 15680 8906 15736
rect 8574 12960 8630 13016
rect 8574 12688 8630 12744
rect 9126 15408 9182 15464
rect 9034 14612 9090 14648
rect 9034 14592 9036 14612
rect 9036 14592 9088 14612
rect 9088 14592 9090 14612
rect 9218 13524 9274 13560
rect 9218 13504 9220 13524
rect 9220 13504 9272 13524
rect 9272 13504 9274 13524
rect 8574 9424 8630 9480
rect 8482 8880 8538 8936
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7470 6160 7526 6216
rect 6918 5616 6974 5672
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 8758 8492 8814 8528
rect 8758 8472 8760 8492
rect 8760 8472 8812 8492
rect 8812 8472 8814 8492
rect 10506 19760 10562 19816
rect 10414 19660 10416 19680
rect 10416 19660 10468 19680
rect 10468 19660 10470 19680
rect 10414 19624 10470 19660
rect 10322 19488 10378 19544
rect 10230 16632 10286 16688
rect 10782 17448 10838 17504
rect 9494 15408 9550 15464
rect 9494 13368 9550 13424
rect 9954 15852 9956 15872
rect 9956 15852 10008 15872
rect 10008 15852 10010 15872
rect 9954 15816 10010 15852
rect 9678 15408 9734 15464
rect 10138 15000 10194 15056
rect 10138 13368 10194 13424
rect 9218 10668 9274 10704
rect 9218 10648 9220 10668
rect 9220 10648 9272 10668
rect 9272 10648 9274 10668
rect 8850 6840 8906 6896
rect 8298 3032 8354 3088
rect 9678 11872 9734 11928
rect 10414 13640 10470 13696
rect 10598 13096 10654 13152
rect 10598 12824 10654 12880
rect 10598 10668 10654 10704
rect 10598 10648 10600 10668
rect 10600 10648 10652 10668
rect 10652 10648 10654 10668
rect 11886 23976 11942 24032
rect 12530 24248 12586 24304
rect 12438 23976 12494 24032
rect 11702 23568 11758 23624
rect 11886 23568 11942 23624
rect 11426 21528 11482 21584
rect 11334 20304 11390 20360
rect 11150 20168 11206 20224
rect 11242 19896 11298 19952
rect 11058 19352 11114 19408
rect 10874 16768 10930 16824
rect 10782 15272 10838 15328
rect 10598 10104 10654 10160
rect 10598 9580 10654 9616
rect 10966 14476 11022 14512
rect 10966 14456 10968 14476
rect 10968 14456 11020 14476
rect 11020 14456 11022 14476
rect 11426 19216 11482 19272
rect 11518 18672 11574 18728
rect 11426 18536 11482 18592
rect 11150 16904 11206 16960
rect 11150 16224 11206 16280
rect 11242 15272 11298 15328
rect 11334 14184 11390 14240
rect 11242 13912 11298 13968
rect 10966 12008 11022 12064
rect 10598 9560 10600 9580
rect 10600 9560 10652 9580
rect 10652 9560 10654 9580
rect 10414 7384 10470 7440
rect 10874 8472 10930 8528
rect 11242 11892 11298 11928
rect 11242 11872 11244 11892
rect 11244 11872 11296 11892
rect 11296 11872 11298 11892
rect 11518 14456 11574 14512
rect 11518 12416 11574 12472
rect 11702 21120 11758 21176
rect 11702 20204 11704 20224
rect 11704 20204 11756 20224
rect 11756 20204 11758 20224
rect 11702 20168 11758 20204
rect 12070 20984 12126 21040
rect 12622 23432 12678 23488
rect 13450 25472 13506 25528
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12162 20576 12218 20632
rect 11886 19216 11942 19272
rect 11702 15272 11758 15328
rect 11702 14048 11758 14104
rect 11702 12552 11758 12608
rect 11886 16632 11942 16688
rect 12162 20168 12218 20224
rect 12070 19352 12126 19408
rect 12438 20032 12494 20088
rect 12162 17856 12218 17912
rect 11886 14048 11942 14104
rect 12438 17992 12494 18048
rect 12714 20576 12770 20632
rect 12714 20304 12770 20360
rect 12622 20168 12678 20224
rect 12530 16768 12586 16824
rect 12530 16632 12586 16688
rect 12438 16496 12494 16552
rect 12254 15816 12310 15872
rect 12346 15680 12402 15736
rect 12530 15952 12586 16008
rect 12438 15544 12494 15600
rect 12346 15272 12402 15328
rect 12254 14728 12310 14784
rect 12254 13640 12310 13696
rect 13818 25608 13874 25664
rect 13726 24520 13782 24576
rect 13818 24384 13874 24440
rect 15382 26288 15438 26344
rect 14278 24656 14334 24712
rect 14094 23588 14150 23624
rect 14094 23568 14096 23588
rect 14096 23568 14148 23588
rect 14148 23568 14150 23588
rect 13174 22752 13230 22808
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 13818 23432 13874 23488
rect 13358 21256 13414 21312
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 13358 20712 13414 20768
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 13726 21256 13782 21312
rect 13634 21120 13690 21176
rect 13542 20712 13598 20768
rect 13818 20848 13874 20904
rect 13818 20712 13874 20768
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12990 18128 13046 18184
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13726 20168 13782 20224
rect 13726 19760 13782 19816
rect 13818 19624 13874 19680
rect 13726 18128 13782 18184
rect 13726 17448 13782 17504
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13450 16360 13506 16416
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12438 12552 12494 12608
rect 12346 12416 12402 12472
rect 11150 4120 11206 4176
rect 10138 2352 10194 2408
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12622 12688 12678 12744
rect 12530 12280 12586 12336
rect 12346 10920 12402 10976
rect 12162 8084 12218 8120
rect 12162 8064 12164 8084
rect 12164 8064 12216 8084
rect 12216 8064 12218 8084
rect 12530 10240 12586 10296
rect 14370 22616 14426 22672
rect 14554 23044 14610 23080
rect 14554 23024 14556 23044
rect 14556 23024 14608 23044
rect 14608 23024 14610 23044
rect 14830 23024 14886 23080
rect 14922 22888 14978 22944
rect 14278 21120 14334 21176
rect 14646 21120 14702 21176
rect 14370 20884 14372 20904
rect 14372 20884 14424 20904
rect 14424 20884 14426 20904
rect 14370 20848 14426 20884
rect 14554 20032 14610 20088
rect 14462 18944 14518 19000
rect 14186 18536 14242 18592
rect 14002 16940 14004 16960
rect 14004 16940 14056 16960
rect 14056 16940 14058 16960
rect 14002 16904 14058 16940
rect 13818 15700 13874 15736
rect 13818 15680 13820 15700
rect 13820 15680 13872 15700
rect 13872 15680 13874 15700
rect 12806 13776 12862 13832
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13358 13504 13414 13560
rect 13082 12960 13138 13016
rect 13082 12688 13138 12744
rect 13266 12688 13322 12744
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12806 12280 12862 12336
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 13450 11464 13506 11520
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12714 9324 12716 9344
rect 12716 9324 12768 9344
rect 12768 9324 12770 9344
rect 12714 9288 12770 9324
rect 12346 6432 12402 6488
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12898 6568 12954 6624
rect 13450 10376 13506 10432
rect 14094 16224 14150 16280
rect 14094 15816 14150 15872
rect 14094 12688 14150 12744
rect 14002 12416 14058 12472
rect 13818 11192 13874 11248
rect 13542 6060 13544 6080
rect 13544 6060 13596 6080
rect 13596 6060 13598 6080
rect 13542 6024 13598 6060
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 13542 5364 13598 5400
rect 13542 5344 13544 5364
rect 13544 5344 13596 5364
rect 13596 5344 13598 5364
rect 13358 3576 13414 3632
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14002 10104 14058 10160
rect 14002 8200 14058 8256
rect 13818 7284 13820 7304
rect 13820 7284 13872 7304
rect 13872 7284 13874 7304
rect 13818 7248 13874 7284
rect 14370 17176 14426 17232
rect 14370 14728 14426 14784
rect 14830 20440 14886 20496
rect 15290 21528 15346 21584
rect 15198 20712 15254 20768
rect 15106 20304 15162 20360
rect 14922 19352 14978 19408
rect 14462 14320 14518 14376
rect 15106 18808 15162 18864
rect 15014 17312 15070 17368
rect 15382 20440 15438 20496
rect 16026 23704 16082 23760
rect 16026 23160 16082 23216
rect 15750 22500 15806 22536
rect 15750 22480 15752 22500
rect 15752 22480 15804 22500
rect 15804 22480 15806 22500
rect 15934 22480 15990 22536
rect 15658 20848 15714 20904
rect 15474 20032 15530 20088
rect 15474 19760 15530 19816
rect 14646 15000 14702 15056
rect 14278 13096 14334 13152
rect 14370 11328 14426 11384
rect 14738 12824 14794 12880
rect 14554 10512 14610 10568
rect 14462 8880 14518 8936
rect 15198 13096 15254 13152
rect 15198 12588 15200 12608
rect 15200 12588 15252 12608
rect 15252 12588 15254 12608
rect 15198 12552 15254 12588
rect 15566 19488 15622 19544
rect 15566 18944 15622 19000
rect 15750 20168 15806 20224
rect 15658 16632 15714 16688
rect 16026 22072 16082 22128
rect 16210 23160 16266 23216
rect 16118 21256 16174 21312
rect 16210 19216 16266 19272
rect 16762 26016 16818 26072
rect 16486 24112 16542 24168
rect 16394 21392 16450 21448
rect 16670 21392 16726 21448
rect 16486 19352 16542 19408
rect 16394 19216 16450 19272
rect 17406 24268 17462 24304
rect 17406 24248 17408 24268
rect 17408 24248 17460 24268
rect 17460 24248 17462 24268
rect 17130 23432 17186 23488
rect 17682 23976 17738 24032
rect 16854 22752 16910 22808
rect 16854 20748 16856 20768
rect 16856 20748 16908 20768
rect 16908 20748 16910 20768
rect 16854 20712 16910 20748
rect 17406 21936 17462 21992
rect 17590 22752 17646 22808
rect 17498 20984 17554 21040
rect 17498 20576 17554 20632
rect 15934 16768 15990 16824
rect 16118 16904 16174 16960
rect 15474 13232 15530 13288
rect 15474 12552 15530 12608
rect 15290 12316 15292 12336
rect 15292 12316 15344 12336
rect 15344 12316 15346 12336
rect 15290 12280 15346 12316
rect 15198 11056 15254 11112
rect 15198 10376 15254 10432
rect 15290 10240 15346 10296
rect 15474 9696 15530 9752
rect 15106 7964 15108 7984
rect 15108 7964 15160 7984
rect 15160 7964 15162 7984
rect 15106 7928 15162 7964
rect 15290 7928 15346 7984
rect 15382 6704 15438 6760
rect 15842 15544 15898 15600
rect 15934 15272 15990 15328
rect 16118 15136 16174 15192
rect 16486 18164 16488 18184
rect 16488 18164 16540 18184
rect 16540 18164 16542 18184
rect 16486 18128 16542 18164
rect 16762 18536 16818 18592
rect 16486 16768 16542 16824
rect 16394 16496 16450 16552
rect 16118 13504 16174 13560
rect 16118 13096 16174 13152
rect 16578 15700 16634 15736
rect 16578 15680 16580 15700
rect 16580 15680 16632 15700
rect 16632 15680 16634 15700
rect 16394 13096 16450 13152
rect 16118 8608 16174 8664
rect 16302 8372 16304 8392
rect 16304 8372 16356 8392
rect 16356 8372 16358 8392
rect 16302 8336 16358 8372
rect 16670 14592 16726 14648
rect 17038 18944 17094 19000
rect 16946 16632 17002 16688
rect 17314 18944 17370 19000
rect 17498 20032 17554 20088
rect 18602 25744 18658 25800
rect 18142 24792 18198 24848
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 18142 22072 18198 22128
rect 18234 21972 18236 21992
rect 18236 21972 18288 21992
rect 18288 21972 18290 21992
rect 18234 21936 18290 21972
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 18418 23160 18474 23216
rect 18694 23704 18750 23760
rect 18602 22752 18658 22808
rect 18602 21664 18658 21720
rect 17590 19660 17592 19680
rect 17592 19660 17644 19680
rect 17644 19660 17646 19680
rect 17590 19624 17646 19660
rect 17774 20168 17830 20224
rect 17406 18400 17462 18456
rect 17222 17720 17278 17776
rect 17038 16224 17094 16280
rect 16946 15852 16948 15872
rect 16948 15852 17000 15872
rect 17000 15852 17002 15872
rect 16946 15816 17002 15852
rect 16670 14048 16726 14104
rect 16762 12300 16818 12336
rect 16762 12280 16764 12300
rect 16764 12280 16816 12300
rect 16816 12280 16818 12300
rect 17222 16904 17278 16960
rect 17222 15564 17278 15600
rect 17222 15544 17224 15564
rect 17224 15544 17276 15564
rect 17276 15544 17278 15564
rect 17222 13640 17278 13696
rect 16762 12008 16818 12064
rect 16854 11636 16856 11656
rect 16856 11636 16908 11656
rect 16908 11636 16910 11656
rect 16854 11600 16910 11636
rect 17038 11192 17094 11248
rect 16578 7248 16634 7304
rect 16026 5752 16082 5808
rect 16302 5752 16358 5808
rect 16670 5344 16726 5400
rect 16486 5092 16542 5128
rect 16486 5072 16488 5092
rect 16488 5072 16540 5092
rect 16540 5072 16542 5092
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18326 19916 18382 19952
rect 18326 19896 18328 19916
rect 18328 19896 18380 19916
rect 18380 19896 18382 19916
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18418 18944 18474 19000
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17682 17720 17738 17776
rect 17590 16632 17646 16688
rect 17590 14456 17646 14512
rect 17590 14320 17646 14376
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17958 16768 18014 16824
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18510 17992 18566 18048
rect 18694 19080 18750 19136
rect 19062 24248 19118 24304
rect 19062 23024 19118 23080
rect 18878 22480 18934 22536
rect 18878 22072 18934 22128
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17958 15000 18014 15056
rect 17774 14456 17830 14512
rect 17590 12960 17646 13016
rect 16946 5908 17002 5944
rect 16946 5888 16948 5908
rect 16948 5888 17000 5908
rect 17000 5888 17002 5908
rect 17130 4820 17186 4856
rect 17130 4800 17132 4820
rect 17132 4800 17184 4820
rect 17184 4800 17186 4820
rect 17038 3984 17094 4040
rect 17498 10784 17554 10840
rect 18418 15952 18474 16008
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17866 12416 17922 12472
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17866 11736 17922 11792
rect 18050 11736 18106 11792
rect 18602 12960 18658 13016
rect 18510 12280 18566 12336
rect 17958 11056 18014 11112
rect 18510 11328 18566 11384
rect 18326 11056 18382 11112
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17498 5208 17554 5264
rect 17498 4256 17554 4312
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17774 6432 17830 6488
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17958 4528 18014 4584
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18234 3712 18290 3768
rect 18970 18808 19026 18864
rect 19614 26152 19670 26208
rect 20350 26832 20406 26888
rect 20074 25880 20130 25936
rect 19430 24248 19486 24304
rect 19338 23568 19394 23624
rect 19706 22616 19762 22672
rect 19614 22480 19670 22536
rect 19522 20440 19578 20496
rect 19982 22072 20038 22128
rect 20718 24112 20774 24168
rect 20994 25336 21050 25392
rect 21638 25064 21694 25120
rect 20902 23432 20958 23488
rect 20810 23296 20866 23352
rect 19798 21800 19854 21856
rect 19706 20868 19762 20904
rect 19706 20848 19708 20868
rect 19708 20848 19760 20868
rect 19760 20848 19762 20868
rect 19338 20204 19340 20224
rect 19340 20204 19392 20224
rect 19392 20204 19394 20224
rect 19338 20168 19394 20204
rect 18878 12588 18880 12608
rect 18880 12588 18932 12608
rect 18932 12588 18934 12608
rect 18878 12552 18934 12588
rect 18418 7112 18474 7168
rect 18970 10376 19026 10432
rect 18970 10104 19026 10160
rect 18510 6024 18566 6080
rect 18878 5636 18934 5672
rect 18878 5616 18880 5636
rect 18880 5616 18932 5636
rect 18932 5616 18934 5636
rect 19246 15136 19302 15192
rect 19154 12688 19210 12744
rect 19614 20304 19670 20360
rect 19614 18808 19670 18864
rect 19706 17992 19762 18048
rect 20810 22636 20866 22672
rect 20810 22616 20812 22636
rect 20812 22616 20864 22636
rect 20864 22616 20866 22636
rect 20350 22108 20352 22128
rect 20352 22108 20404 22128
rect 20404 22108 20406 22128
rect 20350 22072 20406 22108
rect 20534 21936 20590 21992
rect 20074 21528 20130 21584
rect 19890 20576 19946 20632
rect 19982 19080 20038 19136
rect 19430 15428 19486 15464
rect 19430 15408 19432 15428
rect 19432 15408 19484 15428
rect 19484 15408 19486 15428
rect 19614 15308 19616 15328
rect 19616 15308 19668 15328
rect 19668 15308 19670 15328
rect 19614 15272 19670 15308
rect 19522 13252 19578 13288
rect 19522 13232 19524 13252
rect 19524 13232 19576 13252
rect 19576 13232 19578 13252
rect 19430 13096 19486 13152
rect 19430 12552 19486 12608
rect 19338 11192 19394 11248
rect 19430 10512 19486 10568
rect 19430 10376 19486 10432
rect 19338 10260 19394 10296
rect 19338 10240 19340 10260
rect 19340 10240 19392 10260
rect 19392 10240 19394 10260
rect 19246 7792 19302 7848
rect 19062 5752 19118 5808
rect 19062 5616 19118 5672
rect 18878 3984 18934 4040
rect 18602 3848 18658 3904
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 19062 3032 19118 3088
rect 19706 12416 19762 12472
rect 19614 12008 19670 12064
rect 19614 11328 19670 11384
rect 20442 20576 20498 20632
rect 20626 21256 20682 21312
rect 20902 21120 20958 21176
rect 20810 20032 20866 20088
rect 20442 19216 20498 19272
rect 20350 14592 20406 14648
rect 21454 22752 21510 22808
rect 21362 21800 21418 21856
rect 21914 24928 21970 24984
rect 22006 24656 22062 24712
rect 21822 24384 21878 24440
rect 21270 21392 21326 21448
rect 21454 21256 21510 21312
rect 21270 20848 21326 20904
rect 21086 19372 21142 19408
rect 21086 19352 21088 19372
rect 21088 19352 21140 19372
rect 21140 19352 21142 19372
rect 20534 17856 20590 17912
rect 20442 14220 20444 14240
rect 20444 14220 20496 14240
rect 20496 14220 20498 14240
rect 20442 14184 20498 14220
rect 20442 14048 20498 14104
rect 20258 13504 20314 13560
rect 20258 13096 20314 13152
rect 20166 12824 20222 12880
rect 19430 2896 19486 2952
rect 19982 6196 19984 6216
rect 19984 6196 20036 6216
rect 20036 6196 20038 6216
rect 19982 6160 20038 6196
rect 19614 2488 19670 2544
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 20718 16768 20774 16824
rect 21178 18944 21234 19000
rect 21086 18128 21142 18184
rect 20994 17604 21050 17640
rect 20994 17584 20996 17604
rect 20996 17584 21048 17604
rect 21048 17584 21050 17604
rect 20718 14864 20774 14920
rect 20810 13640 20866 13696
rect 20350 12280 20406 12336
rect 20534 10920 20590 10976
rect 22466 24520 22522 24576
rect 21914 22208 21970 22264
rect 21730 20576 21786 20632
rect 21454 15136 21510 15192
rect 21546 14764 21548 14784
rect 21548 14764 21600 14784
rect 21600 14764 21602 14784
rect 21546 14728 21602 14764
rect 21362 13676 21364 13696
rect 21364 13676 21416 13696
rect 21416 13676 21418 13696
rect 21362 13640 21418 13676
rect 22190 22072 22246 22128
rect 21270 13096 21326 13152
rect 21454 13132 21456 13152
rect 21456 13132 21508 13152
rect 21508 13132 21510 13152
rect 21454 13096 21510 13132
rect 21362 12824 21418 12880
rect 20810 6316 20866 6352
rect 20810 6296 20812 6316
rect 20812 6296 20864 6316
rect 20864 6296 20866 6316
rect 21178 11056 21234 11112
rect 25870 26696 25926 26752
rect 25686 26424 25742 26480
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 23386 25472 23442 25528
rect 23386 24792 23442 24848
rect 23294 23024 23350 23080
rect 22742 22344 22798 22400
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22466 21664 22522 21720
rect 22834 21664 22890 21720
rect 22190 20848 22246 20904
rect 22190 20576 22246 20632
rect 22742 21528 22798 21584
rect 22558 20984 22614 21040
rect 22190 19352 22246 19408
rect 22650 20848 22706 20904
rect 22558 20748 22560 20768
rect 22560 20748 22612 20768
rect 22612 20748 22614 20768
rect 22558 20712 22614 20748
rect 22466 19488 22522 19544
rect 22190 16904 22246 16960
rect 22098 16360 22154 16416
rect 22006 16224 22062 16280
rect 22098 15952 22154 16008
rect 21914 15816 21970 15872
rect 22006 15680 22062 15736
rect 21914 14864 21970 14920
rect 21822 14592 21878 14648
rect 21546 12280 21602 12336
rect 21730 13812 21732 13832
rect 21732 13812 21784 13832
rect 21784 13812 21786 13832
rect 21730 13776 21786 13812
rect 21730 13368 21786 13424
rect 21730 12844 21786 12880
rect 21730 12824 21732 12844
rect 21732 12824 21784 12844
rect 21784 12824 21786 12844
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22834 20848 22890 20904
rect 23110 20596 23166 20632
rect 23110 20576 23112 20596
rect 23112 20576 23164 20596
rect 23164 20576 23166 20596
rect 23754 24248 23810 24304
rect 22742 19080 22798 19136
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23018 19660 23020 19680
rect 23020 19660 23072 19680
rect 23072 19660 23074 19680
rect 23018 19624 23074 19660
rect 23570 20712 23626 20768
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22374 13776 22430 13832
rect 22006 13096 22062 13152
rect 22006 12824 22062 12880
rect 21822 12280 21878 12336
rect 21730 11464 21786 11520
rect 22190 12552 22246 12608
rect 22098 9016 22154 9072
rect 22742 18264 22798 18320
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22834 17584 22890 17640
rect 22650 15000 22706 15056
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23202 16632 23258 16688
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22742 13912 22798 13968
rect 22650 12688 22706 12744
rect 22650 12588 22652 12608
rect 22652 12588 22704 12608
rect 22704 12588 22706 12608
rect 22650 12552 22706 12588
rect 23018 14048 23074 14104
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22926 13368 22982 13424
rect 23018 13232 23074 13288
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22650 9560 22706 9616
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22834 7828 22836 7848
rect 22836 7828 22888 7848
rect 22888 7828 22890 7848
rect 22834 7792 22890 7828
rect 22190 1944 22246 2000
rect 23386 15272 23442 15328
rect 23754 19896 23810 19952
rect 23754 19352 23810 19408
rect 24306 25200 24362 25256
rect 24950 26016 25006 26072
rect 24306 19352 24362 19408
rect 24030 18808 24086 18864
rect 24398 18400 24454 18456
rect 23662 16768 23718 16824
rect 23570 15136 23626 15192
rect 23662 14456 23718 14512
rect 23386 12960 23442 13016
rect 24122 15136 24178 15192
rect 23570 11872 23626 11928
rect 23386 8064 23442 8120
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 23294 6840 23350 6896
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 23386 3984 23442 4040
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 22282 1536 22338 1592
rect 23938 11756 23994 11792
rect 23938 11736 23940 11756
rect 23940 11736 23992 11756
rect 23992 11736 23994 11756
rect 24122 12180 24124 12200
rect 24124 12180 24176 12200
rect 24176 12180 24178 12200
rect 24122 12144 24178 12180
rect 24030 11056 24086 11112
rect 24214 10376 24270 10432
rect 23938 8492 23994 8528
rect 23938 8472 23940 8492
rect 23940 8472 23992 8492
rect 23992 8472 23994 8492
rect 23938 7404 23994 7440
rect 23938 7384 23940 7404
rect 23940 7384 23992 7404
rect 23992 7384 23994 7404
rect 23938 6568 23994 6624
rect 24214 10104 24270 10160
rect 24674 21020 24676 21040
rect 24676 21020 24728 21040
rect 24728 21020 24730 21040
rect 24674 20984 24730 21020
rect 24582 19760 24638 19816
rect 25134 25608 25190 25664
rect 24858 22516 24860 22536
rect 24860 22516 24912 22536
rect 24912 22516 24914 22536
rect 24858 22480 24914 22516
rect 24582 17992 24638 18048
rect 24306 7928 24362 7984
rect 24766 18148 24822 18184
rect 24766 18128 24768 18148
rect 24768 18128 24820 18148
rect 24820 18128 24822 18148
rect 24766 14864 24822 14920
rect 24674 12552 24730 12608
rect 24674 12008 24730 12064
rect 25226 23432 25282 23488
rect 25410 23568 25466 23624
rect 25410 21392 25466 21448
rect 25778 22344 25834 22400
rect 25318 19352 25374 19408
rect 25134 18672 25190 18728
rect 24950 17992 25006 18048
rect 25226 17040 25282 17096
rect 25226 15544 25282 15600
rect 25226 15272 25282 15328
rect 25686 21120 25742 21176
rect 25594 20576 25650 20632
rect 25502 18536 25558 18592
rect 25594 16768 25650 16824
rect 25226 12960 25282 13016
rect 25134 12552 25190 12608
rect 25042 12144 25098 12200
rect 24766 11736 24822 11792
rect 24674 9560 24730 9616
rect 24858 11328 24914 11384
rect 25134 10920 25190 10976
rect 25134 10512 25190 10568
rect 25042 10240 25098 10296
rect 24858 10104 24914 10160
rect 24858 9288 24914 9344
rect 24950 8900 25006 8936
rect 24950 8880 24952 8900
rect 24952 8880 25004 8900
rect 25004 8880 25006 8900
rect 24766 8472 24822 8528
rect 24674 7248 24730 7304
rect 24582 5208 24638 5264
rect 24950 7656 25006 7712
rect 24766 6024 24822 6080
rect 24950 5636 25006 5672
rect 24950 5616 24952 5636
rect 24952 5616 25004 5636
rect 25004 5616 25006 5636
rect 24858 4800 24914 4856
rect 24950 4392 25006 4448
rect 24950 3576 25006 3632
rect 24858 2760 24914 2816
rect 23386 1128 23442 1184
rect 24950 2372 25006 2408
rect 24950 2352 24952 2372
rect 24952 2352 25004 2372
rect 25004 2352 25006 2372
rect 26054 23568 26110 23624
rect 25962 23160 26018 23216
rect 26054 22752 26110 22808
rect 25962 19896 26018 19952
rect 25778 15680 25834 15736
rect 25778 15428 25834 15464
rect 25778 15408 25780 15428
rect 25780 15408 25832 15428
rect 25832 15408 25834 15428
rect 25594 13812 25596 13832
rect 25596 13812 25648 13832
rect 25648 13812 25650 13832
rect 25594 13776 25650 13812
rect 26054 14320 26110 14376
rect 26054 14184 26110 14240
rect 25686 6432 25742 6488
rect 25686 3168 25742 3224
rect 25042 720 25098 776
rect 24858 312 24914 368
<< metal3 >>
rect 1209 26890 1275 26893
rect 20345 26890 20411 26893
rect 1209 26888 20411 26890
rect 1209 26832 1214 26888
rect 1270 26832 20350 26888
rect 20406 26832 20411 26888
rect 1209 26830 20411 26832
rect 1209 26827 1275 26830
rect 20345 26827 20411 26830
rect 9254 26692 9260 26756
rect 9324 26754 9330 26756
rect 25865 26754 25931 26757
rect 9324 26752 25931 26754
rect 9324 26696 25870 26752
rect 25926 26696 25931 26752
rect 9324 26694 25931 26696
rect 9324 26692 9330 26694
rect 25865 26691 25931 26694
rect 4889 26618 4955 26621
rect 18454 26618 18460 26620
rect 4889 26616 18460 26618
rect 4889 26560 4894 26616
rect 4950 26560 18460 26616
rect 4889 26558 18460 26560
rect 4889 26555 4955 26558
rect 18454 26556 18460 26558
rect 18524 26556 18530 26620
rect 5165 26482 5231 26485
rect 18822 26482 18828 26484
rect 5165 26480 18828 26482
rect 5165 26424 5170 26480
rect 5226 26424 18828 26480
rect 5165 26422 18828 26424
rect 5165 26419 5231 26422
rect 18822 26420 18828 26422
rect 18892 26420 18898 26484
rect 25681 26482 25747 26485
rect 26200 26482 27000 26512
rect 25681 26480 27000 26482
rect 25681 26424 25686 26480
rect 25742 26424 27000 26480
rect 25681 26422 27000 26424
rect 25681 26419 25747 26422
rect 26200 26392 27000 26422
rect 6126 26284 6132 26348
rect 6196 26346 6202 26348
rect 15377 26346 15443 26349
rect 6196 26344 15443 26346
rect 6196 26288 15382 26344
rect 15438 26288 15443 26344
rect 6196 26286 15443 26288
rect 6196 26284 6202 26286
rect 15377 26283 15443 26286
rect 790 26148 796 26212
rect 860 26210 866 26212
rect 19609 26210 19675 26213
rect 860 26150 1042 26210
rect 860 26148 866 26150
rect 982 26074 1042 26150
rect 2730 26208 19675 26210
rect 2730 26152 19614 26208
rect 19670 26152 19675 26208
rect 2730 26150 19675 26152
rect 2730 26074 2790 26150
rect 19609 26147 19675 26150
rect 16757 26074 16823 26077
rect 982 26014 2790 26074
rect 5030 26072 16823 26074
rect 5030 26016 16762 26072
rect 16818 26016 16823 26072
rect 5030 26014 16823 26016
rect 0 25938 800 25968
rect 3233 25938 3299 25941
rect 0 25936 3299 25938
rect 0 25880 3238 25936
rect 3294 25880 3299 25936
rect 0 25878 3299 25880
rect 0 25848 800 25878
rect 3233 25875 3299 25878
rect 933 25802 999 25805
rect 5030 25802 5090 26014
rect 16757 26011 16823 26014
rect 24945 26074 25011 26077
rect 26200 26074 27000 26104
rect 24945 26072 27000 26074
rect 24945 26016 24950 26072
rect 25006 26016 27000 26072
rect 24945 26014 27000 26016
rect 24945 26011 25011 26014
rect 26200 25984 27000 26014
rect 5206 25876 5212 25940
rect 5276 25938 5282 25940
rect 20069 25938 20135 25941
rect 5276 25936 20135 25938
rect 5276 25880 20074 25936
rect 20130 25880 20135 25936
rect 5276 25878 20135 25880
rect 5276 25876 5282 25878
rect 20069 25875 20135 25878
rect 933 25800 5090 25802
rect 933 25744 938 25800
rect 994 25744 5090 25800
rect 933 25742 5090 25744
rect 7741 25802 7807 25805
rect 18597 25802 18663 25805
rect 7741 25800 18663 25802
rect 7741 25744 7746 25800
rect 7802 25744 18602 25800
rect 18658 25744 18663 25800
rect 7741 25742 18663 25744
rect 933 25739 999 25742
rect 7741 25739 7807 25742
rect 18597 25739 18663 25742
rect 790 25604 796 25668
rect 860 25666 866 25668
rect 13813 25666 13879 25669
rect 860 25664 13879 25666
rect 860 25608 13818 25664
rect 13874 25608 13879 25664
rect 860 25606 13879 25608
rect 860 25604 866 25606
rect 13813 25603 13879 25606
rect 25129 25666 25195 25669
rect 26200 25666 27000 25696
rect 25129 25664 27000 25666
rect 25129 25608 25134 25664
rect 25190 25608 27000 25664
rect 25129 25606 27000 25608
rect 25129 25603 25195 25606
rect 26200 25576 27000 25606
rect 974 25468 980 25532
rect 1044 25530 1050 25532
rect 13445 25530 13511 25533
rect 1044 25528 13511 25530
rect 1044 25472 13450 25528
rect 13506 25472 13511 25528
rect 1044 25470 13511 25472
rect 1044 25468 1050 25470
rect 13445 25467 13511 25470
rect 15142 25468 15148 25532
rect 15212 25530 15218 25532
rect 23381 25530 23447 25533
rect 15212 25528 23447 25530
rect 15212 25472 23386 25528
rect 23442 25472 23447 25528
rect 15212 25470 23447 25472
rect 15212 25468 15218 25470
rect 23381 25467 23447 25470
rect 4654 25332 4660 25396
rect 4724 25394 4730 25396
rect 7741 25394 7807 25397
rect 4724 25392 7807 25394
rect 4724 25336 7746 25392
rect 7802 25336 7807 25392
rect 4724 25334 7807 25336
rect 4724 25332 4730 25334
rect 7741 25331 7807 25334
rect 8334 25332 8340 25396
rect 8404 25394 8410 25396
rect 10961 25394 11027 25397
rect 8404 25392 11027 25394
rect 8404 25336 10966 25392
rect 11022 25336 11027 25392
rect 8404 25334 11027 25336
rect 8404 25332 8410 25334
rect 10961 25331 11027 25334
rect 11094 25332 11100 25396
rect 11164 25394 11170 25396
rect 20989 25394 21055 25397
rect 11164 25392 21055 25394
rect 11164 25336 20994 25392
rect 21050 25336 21055 25392
rect 11164 25334 21055 25336
rect 11164 25332 11170 25334
rect 20989 25331 21055 25334
rect 9438 25196 9444 25260
rect 9508 25258 9514 25260
rect 24301 25258 24367 25261
rect 26200 25258 27000 25288
rect 9508 25256 24367 25258
rect 9508 25200 24306 25256
rect 24362 25200 24367 25256
rect 9508 25198 24367 25200
rect 9508 25196 9514 25198
rect 24301 25195 24367 25198
rect 24534 25198 27000 25258
rect 473 25122 539 25125
rect 933 25122 999 25125
rect 473 25120 999 25122
rect 473 25064 478 25120
rect 534 25064 938 25120
rect 994 25064 999 25120
rect 473 25062 999 25064
rect 473 25059 539 25062
rect 933 25059 999 25062
rect 9806 25060 9812 25124
rect 9876 25122 9882 25124
rect 20662 25122 20668 25124
rect 9876 25062 20668 25122
rect 9876 25060 9882 25062
rect 20662 25060 20668 25062
rect 20732 25060 20738 25124
rect 21633 25122 21699 25125
rect 24534 25122 24594 25198
rect 26200 25168 27000 25198
rect 21633 25120 24594 25122
rect 21633 25064 21638 25120
rect 21694 25064 24594 25120
rect 21633 25062 24594 25064
rect 21633 25059 21699 25062
rect 9622 24924 9628 24988
rect 9692 24986 9698 24988
rect 21909 24986 21975 24989
rect 9692 24984 21975 24986
rect 9692 24928 21914 24984
rect 21970 24928 21975 24984
rect 9692 24926 21975 24928
rect 9692 24924 9698 24926
rect 21909 24923 21975 24926
rect 0 24850 800 24880
rect 3693 24850 3759 24853
rect 0 24848 3759 24850
rect 0 24792 3698 24848
rect 3754 24792 3759 24848
rect 0 24790 3759 24792
rect 0 24760 800 24790
rect 3693 24787 3759 24790
rect 10542 24788 10548 24852
rect 10612 24850 10618 24852
rect 18137 24850 18203 24853
rect 10612 24848 18203 24850
rect 10612 24792 18142 24848
rect 18198 24792 18203 24848
rect 10612 24790 18203 24792
rect 10612 24788 10618 24790
rect 18137 24787 18203 24790
rect 23381 24850 23447 24853
rect 26200 24850 27000 24880
rect 23381 24848 27000 24850
rect 23381 24792 23386 24848
rect 23442 24792 27000 24848
rect 23381 24790 27000 24792
rect 23381 24787 23447 24790
rect 26200 24760 27000 24790
rect 14273 24714 14339 24717
rect 2730 24712 14339 24714
rect 2730 24656 14278 24712
rect 14334 24656 14339 24712
rect 2730 24654 14339 24656
rect 657 24306 723 24309
rect 2730 24306 2790 24654
rect 14273 24651 14339 24654
rect 22001 24714 22067 24717
rect 22001 24712 24226 24714
rect 22001 24656 22006 24712
rect 22062 24656 24226 24712
rect 22001 24654 24226 24656
rect 22001 24651 22067 24654
rect 13721 24578 13787 24581
rect 22461 24578 22527 24581
rect 13721 24576 22527 24578
rect 13721 24520 13726 24576
rect 13782 24520 22466 24576
rect 22522 24520 22527 24576
rect 13721 24518 22527 24520
rect 13721 24515 13787 24518
rect 22461 24515 22527 24518
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 7230 24380 7236 24444
rect 7300 24442 7306 24444
rect 13813 24442 13879 24445
rect 21817 24442 21883 24445
rect 7300 24382 12818 24442
rect 7300 24380 7306 24382
rect 657 24304 2790 24306
rect 657 24248 662 24304
rect 718 24248 2790 24304
rect 657 24246 2790 24248
rect 3969 24306 4035 24309
rect 12525 24306 12591 24309
rect 3969 24304 12591 24306
rect 3969 24248 3974 24304
rect 4030 24248 12530 24304
rect 12586 24248 12591 24304
rect 3969 24246 12591 24248
rect 12758 24306 12818 24382
rect 13813 24440 21883 24442
rect 13813 24384 13818 24440
rect 13874 24384 21822 24440
rect 21878 24384 21883 24440
rect 13813 24382 21883 24384
rect 24166 24442 24226 24654
rect 26200 24442 27000 24472
rect 24166 24382 27000 24442
rect 13813 24379 13879 24382
rect 21817 24379 21883 24382
rect 26200 24352 27000 24382
rect 17401 24306 17467 24309
rect 19057 24308 19123 24309
rect 19006 24306 19012 24308
rect 12758 24304 17467 24306
rect 12758 24248 17406 24304
rect 17462 24248 17467 24304
rect 12758 24246 17467 24248
rect 18966 24246 19012 24306
rect 19076 24304 19123 24308
rect 19118 24248 19123 24304
rect 657 24243 723 24246
rect 3969 24243 4035 24246
rect 12525 24243 12591 24246
rect 17401 24243 17467 24246
rect 19006 24244 19012 24246
rect 19076 24244 19123 24248
rect 19057 24243 19123 24244
rect 19425 24306 19491 24309
rect 23749 24306 23815 24309
rect 19425 24304 23815 24306
rect 19425 24248 19430 24304
rect 19486 24248 23754 24304
rect 23810 24248 23815 24304
rect 19425 24246 23815 24248
rect 19425 24243 19491 24246
rect 23749 24243 23815 24246
rect 3550 24108 3556 24172
rect 3620 24170 3626 24172
rect 3620 24110 8402 24170
rect 3620 24108 3626 24110
rect 1761 24034 1827 24037
rect 2589 24036 2655 24037
rect 2589 24034 2636 24036
rect 1761 24032 2636 24034
rect 1761 23976 1766 24032
rect 1822 23976 2594 24032
rect 1761 23974 2636 23976
rect 1761 23971 1827 23974
rect 2589 23972 2636 23974
rect 2700 23972 2706 24036
rect 8342 24034 8402 24110
rect 11646 24108 11652 24172
rect 11716 24170 11722 24172
rect 16481 24170 16547 24173
rect 11716 24168 16547 24170
rect 11716 24112 16486 24168
rect 16542 24112 16547 24168
rect 11716 24110 16547 24112
rect 11716 24108 11722 24110
rect 16481 24107 16547 24110
rect 16614 24108 16620 24172
rect 16684 24170 16690 24172
rect 20713 24170 20779 24173
rect 16684 24168 20779 24170
rect 16684 24112 20718 24168
rect 20774 24112 20779 24168
rect 16684 24110 20779 24112
rect 16684 24108 16690 24110
rect 20713 24107 20779 24110
rect 11881 24034 11947 24037
rect 8342 24032 11947 24034
rect 8342 23976 11886 24032
rect 11942 23976 11947 24032
rect 8342 23974 11947 23976
rect 2589 23971 2655 23972
rect 11881 23971 11947 23974
rect 12198 23972 12204 24036
rect 12268 24034 12274 24036
rect 12433 24034 12499 24037
rect 12268 24032 12499 24034
rect 12268 23976 12438 24032
rect 12494 23976 12499 24032
rect 12268 23974 12499 23976
rect 12268 23972 12274 23974
rect 12433 23971 12499 23974
rect 13854 23972 13860 24036
rect 13924 24034 13930 24036
rect 17677 24034 17743 24037
rect 13924 24032 17743 24034
rect 13924 23976 17682 24032
rect 17738 23976 17743 24032
rect 13924 23974 17743 23976
rect 13924 23972 13930 23974
rect 17677 23971 17743 23974
rect 24710 23972 24716 24036
rect 24780 24034 24786 24036
rect 26200 24034 27000 24064
rect 24780 23974 27000 24034
rect 24780 23972 24786 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 26200 23944 27000 23974
rect 17946 23903 18262 23904
rect 5022 23836 5028 23900
rect 5092 23898 5098 23900
rect 7281 23898 7347 23901
rect 5092 23896 7347 23898
rect 5092 23840 7286 23896
rect 7342 23840 7347 23896
rect 5092 23838 7347 23840
rect 5092 23836 5098 23838
rect 7281 23835 7347 23838
rect 12390 23838 16314 23898
rect 0 23762 800 23792
rect 2773 23762 2839 23765
rect 0 23760 2839 23762
rect 0 23704 2778 23760
rect 2834 23704 2839 23760
rect 0 23702 2839 23704
rect 0 23672 800 23702
rect 2773 23699 2839 23702
rect 2957 23762 3023 23765
rect 12390 23762 12450 23838
rect 2957 23760 12450 23762
rect 2957 23704 2962 23760
rect 3018 23704 12450 23760
rect 2957 23702 12450 23704
rect 2957 23699 3023 23702
rect 12750 23700 12756 23764
rect 12820 23762 12826 23764
rect 16021 23762 16087 23765
rect 12820 23760 16087 23762
rect 12820 23704 16026 23760
rect 16082 23704 16087 23760
rect 12820 23702 16087 23704
rect 16254 23762 16314 23838
rect 18689 23762 18755 23765
rect 16254 23760 18755 23762
rect 16254 23704 18694 23760
rect 18750 23704 18755 23760
rect 16254 23702 18755 23704
rect 12820 23700 12826 23702
rect 16021 23699 16087 23702
rect 18689 23699 18755 23702
rect 2446 23564 2452 23628
rect 2516 23626 2522 23628
rect 6729 23626 6795 23629
rect 2516 23624 6795 23626
rect 2516 23568 6734 23624
rect 6790 23568 6795 23624
rect 2516 23566 6795 23568
rect 2516 23564 2522 23566
rect 6729 23563 6795 23566
rect 7598 23564 7604 23628
rect 7668 23626 7674 23628
rect 11697 23626 11763 23629
rect 7668 23624 11763 23626
rect 7668 23568 11702 23624
rect 11758 23568 11763 23624
rect 7668 23566 11763 23568
rect 7668 23564 7674 23566
rect 11697 23563 11763 23566
rect 11881 23626 11947 23629
rect 14089 23626 14155 23629
rect 11881 23624 14155 23626
rect 11881 23568 11886 23624
rect 11942 23568 14094 23624
rect 14150 23568 14155 23624
rect 11881 23566 14155 23568
rect 11881 23563 11947 23566
rect 14089 23563 14155 23566
rect 16430 23564 16436 23628
rect 16500 23626 16506 23628
rect 19333 23626 19399 23629
rect 16500 23624 19399 23626
rect 16500 23568 19338 23624
rect 19394 23568 19399 23624
rect 16500 23566 19399 23568
rect 16500 23564 16506 23566
rect 19333 23563 19399 23566
rect 25405 23628 25471 23629
rect 25405 23624 25452 23628
rect 25516 23626 25522 23628
rect 26049 23626 26115 23629
rect 26200 23626 27000 23656
rect 25405 23568 25410 23624
rect 25405 23564 25452 23568
rect 25516 23566 25562 23626
rect 26049 23624 27000 23626
rect 26049 23568 26054 23624
rect 26110 23568 27000 23624
rect 26049 23566 27000 23568
rect 25516 23564 25522 23566
rect 25405 23563 25471 23564
rect 26049 23563 26115 23566
rect 26200 23536 27000 23566
rect 5441 23490 5507 23493
rect 5942 23490 5948 23492
rect 5441 23488 5948 23490
rect 5441 23432 5446 23488
rect 5502 23432 5948 23488
rect 5441 23430 5948 23432
rect 5441 23427 5507 23430
rect 5942 23428 5948 23430
rect 6012 23428 6018 23492
rect 6729 23490 6795 23493
rect 9949 23490 10015 23493
rect 12617 23492 12683 23493
rect 12566 23490 12572 23492
rect 6729 23488 10015 23490
rect 6729 23432 6734 23488
rect 6790 23432 9954 23488
rect 10010 23432 10015 23488
rect 6729 23430 10015 23432
rect 12526 23430 12572 23490
rect 12636 23488 12683 23492
rect 12678 23432 12683 23488
rect 6729 23427 6795 23430
rect 9949 23427 10015 23430
rect 12566 23428 12572 23430
rect 12636 23428 12683 23432
rect 12617 23427 12683 23428
rect 13813 23490 13879 23493
rect 17125 23490 17191 23493
rect 20897 23492 20963 23493
rect 20846 23490 20852 23492
rect 13813 23488 17191 23490
rect 13813 23432 13818 23488
rect 13874 23432 17130 23488
rect 17186 23432 17191 23488
rect 13813 23430 17191 23432
rect 20806 23430 20852 23490
rect 20916 23488 20963 23492
rect 20958 23432 20963 23488
rect 13813 23427 13879 23430
rect 17125 23427 17191 23430
rect 20846 23428 20852 23430
rect 20916 23428 20963 23432
rect 20897 23427 20963 23428
rect 25221 23492 25287 23493
rect 25221 23488 25268 23492
rect 25332 23490 25338 23492
rect 25221 23432 25226 23488
rect 25221 23428 25268 23432
rect 25332 23430 25378 23490
rect 25332 23428 25338 23430
rect 25221 23427 25287 23428
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 4797 23354 4863 23357
rect 12750 23354 12756 23356
rect 4797 23352 12756 23354
rect 4797 23296 4802 23352
rect 4858 23296 12756 23352
rect 4797 23294 12756 23296
rect 4797 23291 4863 23294
rect 12750 23292 12756 23294
rect 12820 23292 12826 23356
rect 16246 23292 16252 23356
rect 16316 23354 16322 23356
rect 20805 23354 20871 23357
rect 16316 23352 20871 23354
rect 16316 23296 20810 23352
rect 20866 23296 20871 23352
rect 16316 23294 20871 23296
rect 16316 23292 16322 23294
rect 20805 23291 20871 23294
rect 2221 23218 2287 23221
rect 16021 23218 16087 23221
rect 2221 23216 16087 23218
rect 2221 23160 2226 23216
rect 2282 23160 16026 23216
rect 16082 23160 16087 23216
rect 2221 23158 16087 23160
rect 2221 23155 2287 23158
rect 16021 23155 16087 23158
rect 16205 23218 16271 23221
rect 18413 23218 18479 23221
rect 16205 23216 18479 23218
rect 16205 23160 16210 23216
rect 16266 23160 18418 23216
rect 18474 23160 18479 23216
rect 16205 23158 18479 23160
rect 16205 23155 16271 23158
rect 18413 23155 18479 23158
rect 25957 23218 26023 23221
rect 26200 23218 27000 23248
rect 25957 23216 27000 23218
rect 25957 23160 25962 23216
rect 26018 23160 27000 23216
rect 25957 23158 27000 23160
rect 25957 23155 26023 23158
rect 26200 23128 27000 23158
rect 1945 23082 2011 23085
rect 14549 23082 14615 23085
rect 1945 23080 14615 23082
rect 1945 23024 1950 23080
rect 2006 23024 14554 23080
rect 14610 23024 14615 23080
rect 1945 23022 14615 23024
rect 1945 23019 2011 23022
rect 14549 23019 14615 23022
rect 14825 23082 14891 23085
rect 19057 23082 19123 23085
rect 14825 23080 19123 23082
rect 14825 23024 14830 23080
rect 14886 23024 19062 23080
rect 19118 23024 19123 23080
rect 14825 23022 19123 23024
rect 14825 23019 14891 23022
rect 19057 23019 19123 23022
rect 23289 23082 23355 23085
rect 25998 23082 26004 23084
rect 23289 23080 26004 23082
rect 23289 23024 23294 23080
rect 23350 23024 26004 23080
rect 23289 23022 26004 23024
rect 23289 23019 23355 23022
rect 25998 23020 26004 23022
rect 26068 23020 26074 23084
rect 8661 22946 8727 22949
rect 14917 22946 14983 22949
rect 8661 22944 14983 22946
rect 8661 22888 8666 22944
rect 8722 22888 14922 22944
rect 14978 22888 14983 22944
rect 8661 22886 14983 22888
rect 8661 22883 8727 22886
rect 14917 22883 14983 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 9029 22810 9095 22813
rect 9806 22810 9812 22812
rect 9029 22808 9812 22810
rect 9029 22752 9034 22808
rect 9090 22752 9812 22808
rect 9029 22750 9812 22752
rect 9029 22747 9095 22750
rect 9806 22748 9812 22750
rect 9876 22748 9882 22812
rect 9949 22810 10015 22813
rect 13169 22810 13235 22813
rect 16849 22810 16915 22813
rect 17585 22810 17651 22813
rect 9949 22808 13235 22810
rect 9949 22752 9954 22808
rect 10010 22752 13174 22808
rect 13230 22752 13235 22808
rect 9949 22750 13235 22752
rect 9949 22747 10015 22750
rect 13169 22747 13235 22750
rect 13310 22750 14658 22810
rect 0 22674 800 22704
rect 3417 22674 3483 22677
rect 0 22672 3483 22674
rect 0 22616 3422 22672
rect 3478 22616 3483 22672
rect 0 22614 3483 22616
rect 0 22584 800 22614
rect 3417 22611 3483 22614
rect 9213 22674 9279 22677
rect 13310 22674 13370 22750
rect 9213 22672 13370 22674
rect 9213 22616 9218 22672
rect 9274 22616 13370 22672
rect 9213 22614 13370 22616
rect 9213 22611 9279 22614
rect 13486 22612 13492 22676
rect 13556 22674 13562 22676
rect 14365 22674 14431 22677
rect 13556 22672 14431 22674
rect 13556 22616 14370 22672
rect 14426 22616 14431 22672
rect 13556 22614 14431 22616
rect 14598 22674 14658 22750
rect 16849 22808 17651 22810
rect 16849 22752 16854 22808
rect 16910 22752 17590 22808
rect 17646 22752 17651 22808
rect 16849 22750 17651 22752
rect 16849 22747 16915 22750
rect 17585 22747 17651 22750
rect 18454 22748 18460 22812
rect 18524 22810 18530 22812
rect 18597 22810 18663 22813
rect 21449 22810 21515 22813
rect 18524 22808 21515 22810
rect 18524 22752 18602 22808
rect 18658 22752 21454 22808
rect 21510 22752 21515 22808
rect 18524 22750 21515 22752
rect 18524 22748 18530 22750
rect 18597 22747 18663 22750
rect 21449 22747 21515 22750
rect 26049 22810 26115 22813
rect 26200 22810 27000 22840
rect 26049 22808 27000 22810
rect 26049 22752 26054 22808
rect 26110 22752 27000 22808
rect 26049 22750 27000 22752
rect 26049 22747 26115 22750
rect 26200 22720 27000 22750
rect 19701 22674 19767 22677
rect 14598 22672 19767 22674
rect 14598 22616 19706 22672
rect 19762 22616 19767 22672
rect 14598 22614 19767 22616
rect 13556 22612 13562 22614
rect 14365 22611 14431 22614
rect 19701 22611 19767 22614
rect 20662 22612 20668 22676
rect 20732 22674 20738 22676
rect 20805 22674 20871 22677
rect 20732 22672 20871 22674
rect 20732 22616 20810 22672
rect 20866 22616 20871 22672
rect 20732 22614 20871 22616
rect 20732 22612 20738 22614
rect 20805 22611 20871 22614
rect 2681 22538 2747 22541
rect 15745 22538 15811 22541
rect 2681 22536 15811 22538
rect 2681 22480 2686 22536
rect 2742 22480 15750 22536
rect 15806 22480 15811 22536
rect 2681 22478 15811 22480
rect 2681 22475 2747 22478
rect 15745 22475 15811 22478
rect 15929 22538 15995 22541
rect 18873 22538 18939 22541
rect 15929 22536 18939 22538
rect 15929 22480 15934 22536
rect 15990 22480 18878 22536
rect 18934 22480 18939 22536
rect 15929 22478 18939 22480
rect 15929 22475 15995 22478
rect 18873 22475 18939 22478
rect 19609 22538 19675 22541
rect 24853 22538 24919 22541
rect 19609 22536 24919 22538
rect 19609 22480 19614 22536
rect 19670 22480 24858 22536
rect 24914 22480 24919 22536
rect 19609 22478 24919 22480
rect 19609 22475 19675 22478
rect 24853 22475 24919 22478
rect 9254 22340 9260 22404
rect 9324 22402 9330 22404
rect 9489 22402 9555 22405
rect 9324 22400 9555 22402
rect 9324 22344 9494 22400
rect 9550 22344 9555 22400
rect 9324 22342 9555 22344
rect 9324 22340 9330 22342
rect 9489 22339 9555 22342
rect 12390 22342 12818 22402
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 3693 22266 3759 22269
rect 3918 22266 3924 22268
rect 3693 22264 3924 22266
rect 3693 22208 3698 22264
rect 3754 22208 3924 22264
rect 3693 22206 3924 22208
rect 3693 22203 3759 22206
rect 3918 22204 3924 22206
rect 3988 22266 3994 22268
rect 12390 22266 12450 22342
rect 3988 22206 12450 22266
rect 3988 22204 3994 22206
rect 1853 22130 1919 22133
rect 3734 22130 3740 22132
rect 1853 22128 3740 22130
rect 1853 22072 1858 22128
rect 1914 22072 3740 22128
rect 1853 22070 3740 22072
rect 1853 22067 1919 22070
rect 3734 22068 3740 22070
rect 3804 22068 3810 22132
rect 4705 22130 4771 22133
rect 12566 22130 12572 22132
rect 4705 22128 12572 22130
rect 4705 22072 4710 22128
rect 4766 22072 12572 22128
rect 4705 22070 12572 22072
rect 4705 22067 4771 22070
rect 12566 22068 12572 22070
rect 12636 22068 12642 22132
rect 12758 22130 12818 22342
rect 14590 22340 14596 22404
rect 14660 22402 14666 22404
rect 22737 22402 22803 22405
rect 14660 22400 22803 22402
rect 14660 22344 22742 22400
rect 22798 22344 22803 22400
rect 14660 22342 22803 22344
rect 14660 22340 14666 22342
rect 22737 22339 22803 22342
rect 25773 22402 25839 22405
rect 26200 22402 27000 22432
rect 25773 22400 27000 22402
rect 25773 22344 25778 22400
rect 25834 22344 27000 22400
rect 25773 22342 27000 22344
rect 25773 22339 25839 22342
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 26200 22312 27000 22342
rect 22946 22271 23262 22272
rect 21909 22266 21975 22269
rect 13494 22264 21975 22266
rect 13494 22208 21914 22264
rect 21970 22208 21975 22264
rect 13494 22206 21975 22208
rect 13494 22130 13554 22206
rect 21909 22203 21975 22206
rect 12758 22070 13554 22130
rect 16021 22130 16087 22133
rect 18137 22130 18203 22133
rect 18873 22132 18939 22133
rect 19977 22132 20043 22133
rect 18454 22130 18460 22132
rect 16021 22128 18460 22130
rect 16021 22072 16026 22128
rect 16082 22072 18142 22128
rect 18198 22072 18460 22128
rect 16021 22070 18460 22072
rect 16021 22067 16087 22070
rect 18137 22067 18203 22070
rect 18454 22068 18460 22070
rect 18524 22068 18530 22132
rect 18822 22130 18828 22132
rect 18782 22070 18828 22130
rect 18892 22128 18939 22132
rect 19926 22130 19932 22132
rect 18934 22072 18939 22128
rect 18822 22068 18828 22070
rect 18892 22068 18939 22072
rect 19886 22070 19932 22130
rect 19996 22128 20043 22132
rect 20038 22072 20043 22128
rect 19926 22068 19932 22070
rect 19996 22068 20043 22072
rect 18873 22067 18939 22068
rect 19977 22067 20043 22068
rect 20345 22130 20411 22133
rect 22185 22130 22251 22133
rect 20345 22128 22251 22130
rect 20345 22072 20350 22128
rect 20406 22072 22190 22128
rect 22246 22072 22251 22128
rect 20345 22070 22251 22072
rect 20345 22067 20411 22070
rect 22185 22067 22251 22070
rect 4337 21994 4403 21997
rect 4613 21994 4679 21997
rect 4337 21992 6746 21994
rect 4337 21936 4342 21992
rect 4398 21936 4618 21992
rect 4674 21936 6746 21992
rect 4337 21934 6746 21936
rect 4337 21931 4403 21934
rect 4613 21931 4679 21934
rect 1894 21660 1900 21724
rect 1964 21722 1970 21724
rect 2129 21722 2195 21725
rect 1964 21720 2195 21722
rect 1964 21664 2134 21720
rect 2190 21664 2195 21720
rect 1964 21662 2195 21664
rect 1964 21660 1970 21662
rect 2129 21659 2195 21662
rect 3877 21722 3943 21725
rect 5165 21722 5231 21725
rect 3877 21720 5231 21722
rect 3877 21664 3882 21720
rect 3938 21664 5170 21720
rect 5226 21664 5231 21720
rect 3877 21662 5231 21664
rect 3877 21659 3943 21662
rect 5165 21659 5231 21662
rect 6494 21586 6500 21588
rect 2730 21526 6500 21586
rect 2497 21450 2563 21453
rect 2730 21450 2790 21526
rect 6494 21524 6500 21526
rect 6564 21524 6570 21588
rect 6686 21586 6746 21934
rect 7414 21932 7420 21996
rect 7484 21994 7490 21996
rect 9121 21994 9187 21997
rect 17401 21994 17467 21997
rect 7484 21934 8770 21994
rect 7484 21932 7490 21934
rect 8710 21858 8770 21934
rect 9121 21992 17467 21994
rect 9121 21936 9126 21992
rect 9182 21936 17406 21992
rect 17462 21936 17467 21992
rect 9121 21934 17467 21936
rect 9121 21931 9187 21934
rect 17401 21931 17467 21934
rect 18229 21994 18295 21997
rect 19190 21994 19196 21996
rect 18229 21992 19196 21994
rect 18229 21936 18234 21992
rect 18290 21936 19196 21992
rect 18229 21934 19196 21936
rect 18229 21931 18295 21934
rect 19190 21932 19196 21934
rect 19260 21932 19266 21996
rect 20529 21994 20595 21997
rect 26200 21994 27000 22024
rect 20529 21992 27000 21994
rect 20529 21936 20534 21992
rect 20590 21936 27000 21992
rect 20529 21934 27000 21936
rect 20529 21931 20595 21934
rect 26200 21904 27000 21934
rect 8710 21798 17786 21858
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 8385 21722 8451 21725
rect 15142 21722 15148 21724
rect 8385 21720 15148 21722
rect 8385 21664 8390 21720
rect 8446 21664 15148 21720
rect 8385 21662 15148 21664
rect 8385 21659 8451 21662
rect 15142 21660 15148 21662
rect 15212 21660 15218 21724
rect 9121 21586 9187 21589
rect 6686 21584 9187 21586
rect 6686 21528 9126 21584
rect 9182 21528 9187 21584
rect 6686 21526 9187 21528
rect 9121 21523 9187 21526
rect 11421 21586 11487 21589
rect 15285 21586 15351 21589
rect 11421 21584 15351 21586
rect 11421 21528 11426 21584
rect 11482 21528 15290 21584
rect 15346 21528 15351 21584
rect 11421 21526 15351 21528
rect 17726 21586 17786 21798
rect 18454 21796 18460 21860
rect 18524 21858 18530 21860
rect 19793 21858 19859 21861
rect 21357 21858 21423 21861
rect 18524 21856 21423 21858
rect 18524 21800 19798 21856
rect 19854 21800 21362 21856
rect 21418 21800 21423 21856
rect 18524 21798 21423 21800
rect 18524 21796 18530 21798
rect 19793 21795 19859 21798
rect 21357 21795 21423 21798
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 18597 21722 18663 21725
rect 22461 21722 22527 21725
rect 22829 21722 22895 21725
rect 18597 21720 22110 21722
rect 18597 21664 18602 21720
rect 18658 21664 22110 21720
rect 18597 21662 22110 21664
rect 18597 21659 18663 21662
rect 20069 21586 20135 21589
rect 20846 21586 20852 21588
rect 17726 21584 20852 21586
rect 17726 21528 20074 21584
rect 20130 21528 20852 21584
rect 17726 21526 20852 21528
rect 11421 21523 11487 21526
rect 15285 21523 15351 21526
rect 20069 21523 20135 21526
rect 20846 21524 20852 21526
rect 20916 21524 20922 21588
rect 2497 21448 2790 21450
rect 2497 21392 2502 21448
rect 2558 21392 2790 21448
rect 2497 21390 2790 21392
rect 6453 21450 6519 21453
rect 7414 21450 7420 21452
rect 6453 21448 7420 21450
rect 6453 21392 6458 21448
rect 6514 21392 7420 21448
rect 6453 21390 7420 21392
rect 2497 21387 2563 21390
rect 6453 21387 6519 21390
rect 7414 21388 7420 21390
rect 7484 21388 7490 21452
rect 16389 21450 16455 21453
rect 9216 21448 16455 21450
rect 9216 21392 16394 21448
rect 16450 21392 16455 21448
rect 9216 21390 16455 21392
rect 9216 21317 9276 21390
rect 16389 21387 16455 21390
rect 16665 21450 16731 21453
rect 21265 21450 21331 21453
rect 16665 21448 21331 21450
rect 16665 21392 16670 21448
rect 16726 21392 21270 21448
rect 21326 21392 21331 21448
rect 16665 21390 21331 21392
rect 22050 21450 22110 21662
rect 22461 21720 22895 21722
rect 22461 21664 22466 21720
rect 22522 21664 22834 21720
rect 22890 21664 22895 21720
rect 22461 21662 22895 21664
rect 22461 21659 22527 21662
rect 22829 21659 22895 21662
rect 22737 21586 22803 21589
rect 26200 21586 27000 21616
rect 22737 21584 27000 21586
rect 22737 21528 22742 21584
rect 22798 21528 27000 21584
rect 22737 21526 27000 21528
rect 22737 21523 22803 21526
rect 26200 21496 27000 21526
rect 25405 21450 25471 21453
rect 22050 21448 25471 21450
rect 22050 21392 25410 21448
rect 25466 21392 25471 21448
rect 22050 21390 25471 21392
rect 16665 21387 16731 21390
rect 21265 21387 21331 21390
rect 25405 21387 25471 21390
rect 6637 21314 6703 21317
rect 8569 21316 8635 21317
rect 8518 21314 8524 21316
rect 6637 21312 8524 21314
rect 8588 21314 8635 21316
rect 8588 21312 8680 21314
rect 6637 21256 6642 21312
rect 6698 21256 8524 21312
rect 8630 21256 8680 21312
rect 6637 21254 8524 21256
rect 6637 21251 6703 21254
rect 8518 21252 8524 21254
rect 8588 21254 8680 21256
rect 9213 21312 9279 21317
rect 9213 21256 9218 21312
rect 9274 21256 9279 21312
rect 8588 21252 8635 21254
rect 8569 21251 8635 21252
rect 9213 21251 9279 21256
rect 13353 21314 13419 21317
rect 13721 21314 13787 21317
rect 13353 21312 13787 21314
rect 13353 21256 13358 21312
rect 13414 21256 13726 21312
rect 13782 21256 13787 21312
rect 13353 21254 13787 21256
rect 13353 21251 13419 21254
rect 13721 21251 13787 21254
rect 16113 21314 16179 21317
rect 20621 21314 20687 21317
rect 16113 21312 20687 21314
rect 16113 21256 16118 21312
rect 16174 21256 20626 21312
rect 20682 21256 20687 21312
rect 16113 21254 20687 21256
rect 16113 21251 16179 21254
rect 20621 21251 20687 21254
rect 21214 21252 21220 21316
rect 21284 21314 21290 21316
rect 21449 21314 21515 21317
rect 21284 21312 21515 21314
rect 21284 21256 21454 21312
rect 21510 21256 21515 21312
rect 21284 21254 21515 21256
rect 21284 21252 21290 21254
rect 21449 21251 21515 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 7005 21178 7071 21181
rect 8569 21178 8635 21181
rect 7005 21176 8635 21178
rect 7005 21120 7010 21176
rect 7066 21120 8574 21176
rect 8630 21120 8635 21176
rect 7005 21118 8635 21120
rect 7005 21115 7071 21118
rect 8569 21115 8635 21118
rect 9397 21178 9463 21181
rect 11697 21178 11763 21181
rect 12198 21178 12204 21180
rect 9397 21176 12204 21178
rect 9397 21120 9402 21176
rect 9458 21120 11702 21176
rect 11758 21120 12204 21176
rect 9397 21118 12204 21120
rect 9397 21115 9463 21118
rect 11697 21115 11763 21118
rect 12198 21116 12204 21118
rect 12268 21116 12274 21180
rect 13629 21178 13695 21181
rect 14273 21178 14339 21181
rect 13629 21176 14339 21178
rect 13629 21120 13634 21176
rect 13690 21120 14278 21176
rect 14334 21120 14339 21176
rect 13629 21118 14339 21120
rect 13629 21115 13695 21118
rect 14273 21115 14339 21118
rect 14641 21178 14707 21181
rect 20897 21178 20963 21181
rect 14641 21176 20963 21178
rect 14641 21120 14646 21176
rect 14702 21120 20902 21176
rect 20958 21120 20963 21176
rect 14641 21118 20963 21120
rect 14641 21115 14707 21118
rect 20897 21115 20963 21118
rect 25681 21178 25747 21181
rect 26200 21178 27000 21208
rect 25681 21176 27000 21178
rect 25681 21120 25686 21176
rect 25742 21120 27000 21176
rect 25681 21118 27000 21120
rect 25681 21115 25747 21118
rect 26200 21088 27000 21118
rect 933 21042 999 21045
rect 9673 21042 9739 21045
rect 12065 21044 12131 21045
rect 12014 21042 12020 21044
rect 933 21040 9739 21042
rect 933 20984 938 21040
rect 994 20984 9678 21040
rect 9734 20984 9739 21040
rect 933 20982 9739 20984
rect 11974 20982 12020 21042
rect 12084 21040 12131 21044
rect 17493 21042 17559 21045
rect 22553 21042 22619 21045
rect 12126 20984 12131 21040
rect 933 20979 999 20982
rect 9673 20979 9739 20982
rect 12014 20980 12020 20982
rect 12084 20980 12131 20984
rect 12065 20979 12131 20980
rect 12390 21040 17559 21042
rect 12390 20984 17498 21040
rect 17554 20984 17559 21040
rect 12390 20982 17559 20984
rect 2221 20906 2287 20909
rect 7005 20906 7071 20909
rect 2221 20904 7071 20906
rect 2221 20848 2226 20904
rect 2282 20848 7010 20904
rect 7066 20848 7071 20904
rect 2221 20846 7071 20848
rect 2221 20843 2287 20846
rect 7005 20843 7071 20846
rect 7281 20906 7347 20909
rect 12390 20906 12450 20982
rect 17493 20979 17559 20982
rect 20440 21040 22619 21042
rect 20440 20984 22558 21040
rect 22614 20984 22619 21040
rect 20440 20982 22619 20984
rect 13813 20906 13879 20909
rect 7281 20904 12450 20906
rect 7281 20848 7286 20904
rect 7342 20848 12450 20904
rect 7281 20846 12450 20848
rect 13310 20904 13879 20906
rect 13310 20848 13818 20904
rect 13874 20848 13879 20904
rect 13310 20846 13879 20848
rect 7281 20843 7347 20846
rect 13310 20773 13370 20846
rect 13813 20843 13879 20846
rect 14365 20906 14431 20909
rect 15653 20906 15719 20909
rect 14365 20904 15719 20906
rect 14365 20848 14370 20904
rect 14426 20848 15658 20904
rect 15714 20848 15719 20904
rect 14365 20846 15719 20848
rect 14365 20843 14431 20846
rect 15653 20843 15719 20846
rect 15878 20844 15884 20908
rect 15948 20906 15954 20908
rect 19701 20906 19767 20909
rect 15948 20904 19767 20906
rect 15948 20848 19706 20904
rect 19762 20848 19767 20904
rect 15948 20846 19767 20848
rect 15948 20844 15954 20846
rect 19701 20843 19767 20846
rect 8753 20772 8819 20773
rect 8702 20708 8708 20772
rect 8772 20770 8819 20772
rect 8772 20768 8864 20770
rect 8814 20712 8864 20768
rect 8772 20710 8864 20712
rect 8772 20708 8819 20710
rect 9806 20708 9812 20772
rect 9876 20770 9882 20772
rect 9949 20770 10015 20773
rect 9876 20768 10015 20770
rect 9876 20712 9954 20768
rect 10010 20712 10015 20768
rect 9876 20710 10015 20712
rect 9876 20708 9882 20710
rect 8753 20707 8819 20708
rect 9949 20707 10015 20710
rect 12022 20710 13186 20770
rect 13310 20768 13419 20773
rect 13310 20712 13358 20768
rect 13414 20712 13419 20768
rect 13310 20710 13419 20712
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 4705 20634 4771 20637
rect 7649 20634 7715 20637
rect 4705 20632 7715 20634
rect 4705 20576 4710 20632
rect 4766 20576 7654 20632
rect 7710 20576 7715 20632
rect 4705 20574 7715 20576
rect 4705 20571 4771 20574
rect 7649 20571 7715 20574
rect 9581 20634 9647 20637
rect 12022 20634 12082 20710
rect 9581 20632 12082 20634
rect 9581 20576 9586 20632
rect 9642 20576 12082 20632
rect 9581 20574 12082 20576
rect 12157 20634 12223 20637
rect 12709 20634 12775 20637
rect 12157 20632 12775 20634
rect 12157 20576 12162 20632
rect 12218 20576 12714 20632
rect 12770 20576 12775 20632
rect 12157 20574 12775 20576
rect 13126 20634 13186 20710
rect 13353 20707 13419 20710
rect 13537 20770 13603 20773
rect 13670 20770 13676 20772
rect 13537 20768 13676 20770
rect 13537 20712 13542 20768
rect 13598 20712 13676 20768
rect 13537 20710 13676 20712
rect 13537 20707 13603 20710
rect 13670 20708 13676 20710
rect 13740 20708 13746 20772
rect 13813 20770 13879 20773
rect 15193 20770 15259 20773
rect 16849 20772 16915 20773
rect 16798 20770 16804 20772
rect 13813 20768 15259 20770
rect 13813 20712 13818 20768
rect 13874 20712 15198 20768
rect 15254 20712 15259 20768
rect 13813 20710 15259 20712
rect 16758 20710 16804 20770
rect 16868 20768 16915 20772
rect 16910 20712 16915 20768
rect 13813 20707 13879 20710
rect 15193 20707 15259 20710
rect 16798 20708 16804 20710
rect 16868 20708 16915 20712
rect 16849 20707 16915 20708
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 20440 20637 20500 20982
rect 22553 20979 22619 20982
rect 24526 20980 24532 21044
rect 24596 21042 24602 21044
rect 24669 21042 24735 21045
rect 24596 21040 24735 21042
rect 24596 20984 24674 21040
rect 24730 20984 24735 21040
rect 24596 20982 24735 20984
rect 24596 20980 24602 20982
rect 24669 20979 24735 20982
rect 21265 20906 21331 20909
rect 22185 20906 22251 20909
rect 21265 20904 22251 20906
rect 21265 20848 21270 20904
rect 21326 20848 22190 20904
rect 22246 20848 22251 20904
rect 21265 20846 22251 20848
rect 21265 20843 21331 20846
rect 22185 20843 22251 20846
rect 22502 20844 22508 20908
rect 22572 20906 22578 20908
rect 22645 20906 22711 20909
rect 22572 20904 22711 20906
rect 22572 20848 22650 20904
rect 22706 20848 22711 20904
rect 22572 20846 22711 20848
rect 22572 20844 22578 20846
rect 22645 20843 22711 20846
rect 22829 20906 22895 20909
rect 22829 20904 24778 20906
rect 22829 20848 22834 20904
rect 22890 20848 24778 20904
rect 22829 20846 24778 20848
rect 22829 20843 22895 20846
rect 21582 20708 21588 20772
rect 21652 20770 21658 20772
rect 22553 20770 22619 20773
rect 23565 20772 23631 20773
rect 23565 20770 23612 20772
rect 21652 20768 22619 20770
rect 21652 20712 22558 20768
rect 22614 20712 22619 20768
rect 21652 20710 22619 20712
rect 23520 20768 23612 20770
rect 23520 20712 23570 20768
rect 23520 20710 23612 20712
rect 21652 20708 21658 20710
rect 22553 20707 22619 20710
rect 23565 20708 23612 20710
rect 23676 20708 23682 20772
rect 24718 20770 24778 20846
rect 26200 20770 27000 20800
rect 24718 20710 27000 20770
rect 23565 20707 23631 20708
rect 26200 20680 27000 20710
rect 17493 20634 17559 20637
rect 19885 20634 19951 20637
rect 13126 20632 17559 20634
rect 13126 20576 17498 20632
rect 17554 20576 17559 20632
rect 13126 20574 17559 20576
rect 9581 20571 9647 20574
rect 12157 20571 12223 20574
rect 12709 20571 12775 20574
rect 17493 20571 17559 20574
rect 18462 20632 19951 20634
rect 18462 20576 19890 20632
rect 19946 20576 19951 20632
rect 18462 20574 19951 20576
rect 7833 20498 7899 20501
rect 14825 20498 14891 20501
rect 15377 20498 15443 20501
rect 7833 20496 12128 20498
rect 7833 20440 7838 20496
rect 7894 20440 12128 20496
rect 7833 20438 12128 20440
rect 7833 20435 7899 20438
rect 6637 20362 6703 20365
rect 9581 20362 9647 20365
rect 6637 20360 9647 20362
rect 6637 20304 6642 20360
rect 6698 20304 9586 20360
rect 9642 20304 9647 20360
rect 6637 20302 9647 20304
rect 6637 20299 6703 20302
rect 9581 20299 9647 20302
rect 10174 20300 10180 20364
rect 10244 20362 10250 20364
rect 11329 20362 11395 20365
rect 10244 20360 11395 20362
rect 10244 20304 11334 20360
rect 11390 20304 11395 20360
rect 10244 20302 11395 20304
rect 12068 20362 12128 20438
rect 12574 20496 15443 20498
rect 12574 20440 14830 20496
rect 14886 20440 15382 20496
rect 15438 20440 15443 20496
rect 12574 20438 15443 20440
rect 12574 20362 12634 20438
rect 14825 20435 14891 20438
rect 15377 20435 15443 20438
rect 17350 20436 17356 20500
rect 17420 20498 17426 20500
rect 18462 20498 18522 20574
rect 19885 20571 19951 20574
rect 20437 20632 20503 20637
rect 20437 20576 20442 20632
rect 20498 20576 20503 20632
rect 20437 20571 20503 20576
rect 21725 20634 21791 20637
rect 22185 20634 22251 20637
rect 23105 20634 23171 20637
rect 25589 20634 25655 20637
rect 21725 20632 25655 20634
rect 21725 20576 21730 20632
rect 21786 20576 22190 20632
rect 22246 20576 23110 20632
rect 23166 20576 25594 20632
rect 25650 20576 25655 20632
rect 21725 20574 25655 20576
rect 21725 20571 21791 20574
rect 22185 20571 22251 20574
rect 23105 20571 23171 20574
rect 25589 20571 25655 20574
rect 17420 20438 18522 20498
rect 19517 20498 19583 20501
rect 20662 20498 20668 20500
rect 19517 20496 20668 20498
rect 19517 20440 19522 20496
rect 19578 20440 20668 20496
rect 19517 20438 20668 20440
rect 17420 20436 17426 20438
rect 19517 20435 19583 20438
rect 20662 20436 20668 20438
rect 20732 20436 20738 20500
rect 12068 20302 12634 20362
rect 12709 20362 12775 20365
rect 15101 20362 15167 20365
rect 12709 20360 15167 20362
rect 12709 20304 12714 20360
rect 12770 20304 15106 20360
rect 15162 20304 15167 20360
rect 12709 20302 15167 20304
rect 10244 20300 10250 20302
rect 11329 20299 11395 20302
rect 12709 20299 12775 20302
rect 15101 20299 15167 20302
rect 16982 20300 16988 20364
rect 17052 20362 17058 20364
rect 19609 20362 19675 20365
rect 17052 20360 19675 20362
rect 17052 20304 19614 20360
rect 19670 20304 19675 20360
rect 17052 20302 19675 20304
rect 17052 20300 17058 20302
rect 19609 20299 19675 20302
rect 22318 20300 22324 20364
rect 22388 20362 22394 20364
rect 26200 20362 27000 20392
rect 22388 20302 27000 20362
rect 22388 20300 22394 20302
rect 26200 20272 27000 20302
rect 8845 20226 8911 20229
rect 11145 20226 11211 20229
rect 11697 20228 11763 20229
rect 8845 20224 11211 20226
rect 8845 20168 8850 20224
rect 8906 20168 11150 20224
rect 11206 20168 11211 20224
rect 8845 20166 11211 20168
rect 8845 20163 8911 20166
rect 11145 20163 11211 20166
rect 11646 20164 11652 20228
rect 11716 20226 11763 20228
rect 12157 20226 12223 20229
rect 12617 20226 12683 20229
rect 11716 20224 11808 20226
rect 11758 20168 11808 20224
rect 11716 20166 11808 20168
rect 12157 20224 12683 20226
rect 12157 20168 12162 20224
rect 12218 20168 12622 20224
rect 12678 20168 12683 20224
rect 12157 20166 12683 20168
rect 11716 20164 11763 20166
rect 11697 20163 11763 20164
rect 12157 20163 12223 20166
rect 12617 20163 12683 20166
rect 13721 20226 13787 20229
rect 15745 20226 15811 20229
rect 17769 20226 17835 20229
rect 19333 20228 19399 20229
rect 19333 20226 19380 20228
rect 13721 20224 17835 20226
rect 13721 20168 13726 20224
rect 13782 20168 15750 20224
rect 15806 20168 17774 20224
rect 17830 20168 17835 20224
rect 13721 20166 17835 20168
rect 19288 20224 19380 20226
rect 19288 20168 19338 20224
rect 19288 20166 19380 20168
rect 13721 20163 13787 20166
rect 15745 20163 15811 20166
rect 17769 20163 17835 20166
rect 19333 20164 19380 20166
rect 19444 20164 19450 20228
rect 19333 20163 19399 20164
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 8753 20090 8819 20093
rect 12433 20090 12499 20093
rect 12566 20090 12572 20092
rect 8753 20088 11162 20090
rect 8753 20032 8758 20088
rect 8814 20032 11162 20088
rect 8753 20030 11162 20032
rect 8753 20027 8819 20030
rect 6678 19892 6684 19956
rect 6748 19954 6754 19956
rect 10542 19954 10548 19956
rect 6748 19894 10548 19954
rect 6748 19892 6754 19894
rect 10542 19892 10548 19894
rect 10612 19892 10618 19956
rect 7373 19818 7439 19821
rect 9213 19818 9279 19821
rect 7373 19816 9279 19818
rect 7373 19760 7378 19816
rect 7434 19760 9218 19816
rect 9274 19760 9279 19816
rect 7373 19758 9279 19760
rect 7373 19755 7439 19758
rect 9213 19755 9279 19758
rect 10501 19818 10567 19821
rect 11102 19818 11162 20030
rect 12433 20088 12572 20090
rect 12433 20032 12438 20088
rect 12494 20032 12572 20088
rect 12433 20030 12572 20032
rect 12433 20027 12499 20030
rect 12566 20028 12572 20030
rect 12636 20028 12642 20092
rect 14549 20090 14615 20093
rect 15469 20090 15535 20093
rect 14549 20088 15535 20090
rect 14549 20032 14554 20088
rect 14610 20032 15474 20088
rect 15530 20032 15535 20088
rect 14549 20030 15535 20032
rect 14549 20027 14615 20030
rect 15469 20027 15535 20030
rect 17493 20090 17559 20093
rect 20805 20090 20871 20093
rect 17493 20088 20871 20090
rect 17493 20032 17498 20088
rect 17554 20032 20810 20088
rect 20866 20032 20871 20088
rect 17493 20030 20871 20032
rect 17493 20027 17559 20030
rect 20805 20027 20871 20030
rect 11237 19954 11303 19957
rect 18321 19954 18387 19957
rect 11237 19952 18387 19954
rect 11237 19896 11242 19952
rect 11298 19896 18326 19952
rect 18382 19896 18387 19952
rect 11237 19894 18387 19896
rect 11237 19891 11303 19894
rect 18321 19891 18387 19894
rect 23749 19956 23815 19957
rect 23749 19952 23796 19956
rect 23860 19954 23866 19956
rect 25957 19954 26023 19957
rect 26200 19954 27000 19984
rect 23749 19896 23754 19952
rect 23749 19892 23796 19896
rect 23860 19894 23906 19954
rect 25957 19952 27000 19954
rect 25957 19896 25962 19952
rect 26018 19896 27000 19952
rect 25957 19894 27000 19896
rect 23860 19892 23866 19894
rect 23749 19891 23815 19892
rect 25957 19891 26023 19894
rect 26200 19864 27000 19894
rect 13721 19818 13787 19821
rect 10501 19816 10978 19818
rect 10501 19760 10506 19816
rect 10562 19760 10978 19816
rect 10501 19758 10978 19760
rect 11102 19816 13787 19818
rect 11102 19760 13726 19816
rect 13782 19760 13787 19816
rect 11102 19758 13787 19760
rect 10501 19755 10567 19758
rect 9397 19682 9463 19685
rect 10409 19682 10475 19685
rect 9397 19680 10475 19682
rect 9397 19624 9402 19680
rect 9458 19624 10414 19680
rect 10470 19624 10475 19680
rect 9397 19622 10475 19624
rect 9397 19619 9463 19622
rect 10409 19619 10475 19622
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 10317 19548 10383 19549
rect 10317 19544 10364 19548
rect 10428 19546 10434 19548
rect 10918 19546 10978 19758
rect 13721 19755 13787 19758
rect 15469 19818 15535 19821
rect 24577 19818 24643 19821
rect 15469 19816 24643 19818
rect 15469 19760 15474 19816
rect 15530 19760 24582 19816
rect 24638 19760 24643 19816
rect 15469 19758 24643 19760
rect 15469 19755 15535 19758
rect 24577 19755 24643 19758
rect 13813 19682 13879 19685
rect 17585 19682 17651 19685
rect 13813 19680 17651 19682
rect 13813 19624 13818 19680
rect 13874 19624 17590 19680
rect 17646 19624 17651 19680
rect 13813 19622 17651 19624
rect 13813 19619 13879 19622
rect 17585 19619 17651 19622
rect 21214 19620 21220 19684
rect 21284 19682 21290 19684
rect 23013 19682 23079 19685
rect 21284 19680 23079 19682
rect 21284 19624 23018 19680
rect 23074 19624 23079 19680
rect 21284 19622 23079 19624
rect 21284 19620 21290 19622
rect 23013 19619 23079 19622
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 15561 19546 15627 19549
rect 10317 19488 10322 19544
rect 10317 19484 10364 19488
rect 10428 19486 10474 19546
rect 10918 19544 15627 19546
rect 10918 19488 15566 19544
rect 15622 19488 15627 19544
rect 10918 19486 15627 19488
rect 10428 19484 10434 19486
rect 10317 19483 10383 19484
rect 15561 19483 15627 19486
rect 15694 19484 15700 19548
rect 15764 19546 15770 19548
rect 22461 19546 22527 19549
rect 26200 19546 27000 19576
rect 15764 19486 16682 19546
rect 15764 19484 15770 19486
rect 4061 19410 4127 19413
rect 11053 19410 11119 19413
rect 4061 19408 11119 19410
rect 4061 19352 4066 19408
rect 4122 19352 11058 19408
rect 11114 19352 11119 19408
rect 4061 19350 11119 19352
rect 4061 19347 4127 19350
rect 11053 19347 11119 19350
rect 12065 19410 12131 19413
rect 12198 19410 12204 19412
rect 12065 19408 12204 19410
rect 12065 19352 12070 19408
rect 12126 19352 12204 19408
rect 12065 19350 12204 19352
rect 12065 19347 12131 19350
rect 12198 19348 12204 19350
rect 12268 19348 12274 19412
rect 14038 19348 14044 19412
rect 14108 19410 14114 19412
rect 14917 19410 14983 19413
rect 14108 19408 14983 19410
rect 14108 19352 14922 19408
rect 14978 19352 14983 19408
rect 14108 19350 14983 19352
rect 14108 19348 14114 19350
rect 14917 19347 14983 19350
rect 15142 19348 15148 19412
rect 15212 19410 15218 19412
rect 16481 19410 16547 19413
rect 15212 19408 16547 19410
rect 15212 19352 16486 19408
rect 16542 19352 16547 19408
rect 15212 19350 16547 19352
rect 16622 19410 16682 19486
rect 18462 19544 22527 19546
rect 18462 19488 22466 19544
rect 22522 19488 22527 19544
rect 18462 19486 22527 19488
rect 18462 19410 18522 19486
rect 22461 19483 22527 19486
rect 22694 19486 27000 19546
rect 16622 19350 18522 19410
rect 21081 19410 21147 19413
rect 22185 19410 22251 19413
rect 22694 19410 22754 19486
rect 26200 19456 27000 19486
rect 21081 19408 22251 19410
rect 21081 19352 21086 19408
rect 21142 19352 22190 19408
rect 22246 19352 22251 19408
rect 21081 19350 22251 19352
rect 15212 19348 15218 19350
rect 16481 19347 16547 19350
rect 21081 19347 21147 19350
rect 22185 19347 22251 19350
rect 22326 19350 22754 19410
rect 5574 19212 5580 19276
rect 5644 19274 5650 19276
rect 5809 19274 5875 19277
rect 5644 19272 5875 19274
rect 5644 19216 5814 19272
rect 5870 19216 5875 19272
rect 5644 19214 5875 19216
rect 5644 19212 5650 19214
rect 5809 19211 5875 19214
rect 6310 19212 6316 19276
rect 6380 19274 6386 19276
rect 11421 19274 11487 19277
rect 11881 19276 11947 19277
rect 6380 19272 11487 19274
rect 6380 19216 11426 19272
rect 11482 19216 11487 19272
rect 6380 19214 11487 19216
rect 6380 19212 6386 19214
rect 11421 19211 11487 19214
rect 11830 19212 11836 19276
rect 11900 19274 11947 19276
rect 16205 19274 16271 19277
rect 11900 19272 11992 19274
rect 11942 19216 11992 19272
rect 11900 19214 11992 19216
rect 12390 19272 16271 19274
rect 12390 19216 16210 19272
rect 16266 19216 16271 19272
rect 12390 19214 16271 19216
rect 11900 19212 11947 19214
rect 11881 19211 11947 19212
rect 8569 19138 8635 19141
rect 12390 19138 12450 19214
rect 16205 19211 16271 19214
rect 16389 19274 16455 19277
rect 20437 19274 20503 19277
rect 16389 19272 20503 19274
rect 16389 19216 16394 19272
rect 16450 19216 20442 19272
rect 20498 19216 20503 19272
rect 16389 19214 20503 19216
rect 16389 19211 16455 19214
rect 20437 19211 20503 19214
rect 22134 19212 22140 19276
rect 22204 19274 22210 19276
rect 22326 19274 22386 19350
rect 23422 19348 23428 19412
rect 23492 19410 23498 19412
rect 23749 19410 23815 19413
rect 23492 19408 23815 19410
rect 23492 19352 23754 19408
rect 23810 19352 23815 19408
rect 23492 19350 23815 19352
rect 23492 19348 23498 19350
rect 23749 19347 23815 19350
rect 24301 19410 24367 19413
rect 25313 19410 25379 19413
rect 25630 19410 25636 19412
rect 24301 19408 24410 19410
rect 24301 19352 24306 19408
rect 24362 19352 24410 19408
rect 24301 19347 24410 19352
rect 25313 19408 25636 19410
rect 25313 19352 25318 19408
rect 25374 19352 25636 19408
rect 25313 19350 25636 19352
rect 25313 19347 25379 19350
rect 25630 19348 25636 19350
rect 25700 19348 25706 19412
rect 22204 19214 22386 19274
rect 22204 19212 22210 19214
rect 18689 19138 18755 19141
rect 19977 19140 20043 19141
rect 8569 19136 12450 19138
rect 8569 19080 8574 19136
rect 8630 19080 12450 19136
rect 8569 19078 12450 19080
rect 15334 19136 18755 19138
rect 15334 19080 18694 19136
rect 18750 19080 18755 19136
rect 15334 19078 18755 19080
rect 8569 19075 8635 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 4061 19002 4127 19005
rect 10910 19002 10916 19004
rect 4061 19000 10916 19002
rect 4061 18944 4066 19000
rect 4122 18944 10916 19000
rect 4061 18942 10916 18944
rect 4061 18939 4127 18942
rect 10910 18940 10916 18942
rect 10980 18940 10986 19004
rect 14457 19002 14523 19005
rect 15334 19002 15394 19078
rect 18689 19075 18755 19078
rect 19926 19076 19932 19140
rect 19996 19138 20043 19140
rect 19996 19136 20088 19138
rect 20038 19080 20088 19136
rect 19996 19078 20088 19080
rect 19996 19076 20043 19078
rect 21398 19076 21404 19140
rect 21468 19138 21474 19140
rect 22737 19138 22803 19141
rect 21468 19136 22803 19138
rect 21468 19080 22742 19136
rect 22798 19080 22803 19136
rect 21468 19078 22803 19080
rect 24350 19138 24410 19347
rect 26200 19138 27000 19168
rect 24350 19078 27000 19138
rect 21468 19076 21474 19078
rect 19977 19075 20043 19076
rect 22737 19075 22803 19078
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 26200 19048 27000 19078
rect 22946 19007 23262 19008
rect 14457 19000 15394 19002
rect 14457 18944 14462 19000
rect 14518 18944 15394 19000
rect 14457 18942 15394 18944
rect 15561 19002 15627 19005
rect 16430 19002 16436 19004
rect 15561 19000 16436 19002
rect 15561 18944 15566 19000
rect 15622 18944 16436 19000
rect 15561 18942 16436 18944
rect 14457 18939 14523 18942
rect 15561 18939 15627 18942
rect 16430 18940 16436 18942
rect 16500 18940 16506 19004
rect 17033 19002 17099 19005
rect 17309 19002 17375 19005
rect 17033 19000 17375 19002
rect 17033 18944 17038 19000
rect 17094 18944 17314 19000
rect 17370 18944 17375 19000
rect 17033 18942 17375 18944
rect 17033 18939 17099 18942
rect 17309 18939 17375 18942
rect 17718 18940 17724 19004
rect 17788 19002 17794 19004
rect 18413 19002 18479 19005
rect 17788 19000 18479 19002
rect 17788 18944 18418 19000
rect 18474 18944 18479 19000
rect 17788 18942 18479 18944
rect 17788 18940 17794 18942
rect 18413 18939 18479 18942
rect 21173 19002 21239 19005
rect 22686 19002 22692 19004
rect 21173 19000 22692 19002
rect 21173 18944 21178 19000
rect 21234 18944 22692 19000
rect 21173 18942 22692 18944
rect 21173 18939 21239 18942
rect 22686 18940 22692 18942
rect 22756 18940 22762 19004
rect 4153 18866 4219 18869
rect 15101 18866 15167 18869
rect 4153 18864 15167 18866
rect 4153 18808 4158 18864
rect 4214 18808 15106 18864
rect 15162 18808 15167 18864
rect 4153 18806 15167 18808
rect 4153 18803 4219 18806
rect 15101 18803 15167 18806
rect 16430 18804 16436 18868
rect 16500 18866 16506 18868
rect 18965 18866 19031 18869
rect 19609 18866 19675 18869
rect 16500 18864 19675 18866
rect 16500 18808 18970 18864
rect 19026 18808 19614 18864
rect 19670 18808 19675 18864
rect 16500 18806 19675 18808
rect 16500 18804 16506 18806
rect 18965 18803 19031 18806
rect 19609 18803 19675 18806
rect 24025 18866 24091 18869
rect 24025 18864 25330 18866
rect 24025 18808 24030 18864
rect 24086 18808 25330 18864
rect 24025 18806 25330 18808
rect 24025 18803 24091 18806
rect 4981 18730 5047 18733
rect 9949 18730 10015 18733
rect 4981 18728 10015 18730
rect 4981 18672 4986 18728
rect 5042 18672 9954 18728
rect 10010 18672 10015 18728
rect 4981 18670 10015 18672
rect 4981 18667 5047 18670
rect 9949 18667 10015 18670
rect 11513 18730 11579 18733
rect 25129 18730 25195 18733
rect 11513 18728 25195 18730
rect 11513 18672 11518 18728
rect 11574 18672 25134 18728
rect 25190 18672 25195 18728
rect 11513 18670 25195 18672
rect 25270 18730 25330 18806
rect 26200 18730 27000 18760
rect 25270 18670 27000 18730
rect 11513 18667 11579 18670
rect 25129 18667 25195 18670
rect 26200 18640 27000 18670
rect 9029 18594 9095 18597
rect 9581 18594 9647 18597
rect 9029 18592 9647 18594
rect 9029 18536 9034 18592
rect 9090 18536 9586 18592
rect 9642 18536 9647 18592
rect 9029 18534 9647 18536
rect 9029 18531 9095 18534
rect 9581 18531 9647 18534
rect 11421 18594 11487 18597
rect 14181 18594 14247 18597
rect 11421 18592 14247 18594
rect 11421 18536 11426 18592
rect 11482 18536 14186 18592
rect 14242 18536 14247 18592
rect 11421 18534 14247 18536
rect 11421 18531 11487 18534
rect 14181 18531 14247 18534
rect 16062 18532 16068 18596
rect 16132 18594 16138 18596
rect 16757 18594 16823 18597
rect 16132 18592 16823 18594
rect 16132 18536 16762 18592
rect 16818 18536 16823 18592
rect 16132 18534 16823 18536
rect 16132 18532 16138 18534
rect 16757 18531 16823 18534
rect 19558 18532 19564 18596
rect 19628 18594 19634 18596
rect 25497 18594 25563 18597
rect 19628 18592 25563 18594
rect 19628 18536 25502 18592
rect 25558 18536 25563 18592
rect 19628 18534 25563 18536
rect 19628 18532 19634 18534
rect 25497 18531 25563 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 5942 18396 5948 18460
rect 6012 18458 6018 18460
rect 6177 18458 6243 18461
rect 6012 18456 6243 18458
rect 6012 18400 6182 18456
rect 6238 18400 6243 18456
rect 6012 18398 6243 18400
rect 6012 18396 6018 18398
rect 6177 18395 6243 18398
rect 9070 18396 9076 18460
rect 9140 18458 9146 18460
rect 9305 18458 9371 18461
rect 17401 18458 17467 18461
rect 9140 18456 9371 18458
rect 9140 18400 9310 18456
rect 9366 18400 9371 18456
rect 9140 18398 9371 18400
rect 9140 18396 9146 18398
rect 9305 18395 9371 18398
rect 9446 18456 17467 18458
rect 9446 18400 17406 18456
rect 17462 18400 17467 18456
rect 9446 18398 17467 18400
rect 6361 18322 6427 18325
rect 9446 18322 9506 18398
rect 17401 18395 17467 18398
rect 20478 18396 20484 18460
rect 20548 18458 20554 18460
rect 24393 18458 24459 18461
rect 20548 18456 24459 18458
rect 20548 18400 24398 18456
rect 24454 18400 24459 18456
rect 20548 18398 24459 18400
rect 20548 18396 20554 18398
rect 24393 18395 24459 18398
rect 6361 18320 9506 18322
rect 6361 18264 6366 18320
rect 6422 18264 9506 18320
rect 6361 18262 9506 18264
rect 9949 18322 10015 18325
rect 22737 18322 22803 18325
rect 26200 18322 27000 18352
rect 9949 18320 22110 18322
rect 9949 18264 9954 18320
rect 10010 18264 22110 18320
rect 9949 18262 22110 18264
rect 6361 18259 6427 18262
rect 9949 18259 10015 18262
rect 2262 18124 2268 18188
rect 2332 18186 2338 18188
rect 9121 18186 9187 18189
rect 9254 18186 9260 18188
rect 2332 18126 7666 18186
rect 2332 18124 2338 18126
rect 7606 18050 7666 18126
rect 9121 18184 9260 18186
rect 9121 18128 9126 18184
rect 9182 18128 9260 18184
rect 9121 18126 9260 18128
rect 9121 18123 9187 18126
rect 9254 18124 9260 18126
rect 9324 18124 9330 18188
rect 11278 18124 11284 18188
rect 11348 18186 11354 18188
rect 12985 18186 13051 18189
rect 11348 18184 13051 18186
rect 11348 18128 12990 18184
rect 13046 18128 13051 18184
rect 11348 18126 13051 18128
rect 11348 18124 11354 18126
rect 12985 18123 13051 18126
rect 13721 18186 13787 18189
rect 16481 18186 16547 18189
rect 21081 18186 21147 18189
rect 13721 18184 16547 18186
rect 13721 18128 13726 18184
rect 13782 18128 16486 18184
rect 16542 18128 16547 18184
rect 13721 18126 16547 18128
rect 13721 18123 13787 18126
rect 16481 18123 16547 18126
rect 18278 18184 21147 18186
rect 18278 18128 21086 18184
rect 21142 18128 21147 18184
rect 18278 18126 21147 18128
rect 22050 18186 22110 18262
rect 22737 18320 27000 18322
rect 22737 18264 22742 18320
rect 22798 18264 27000 18320
rect 22737 18262 27000 18264
rect 22737 18259 22803 18262
rect 26200 18232 27000 18262
rect 24761 18186 24827 18189
rect 22050 18184 24827 18186
rect 22050 18128 24766 18184
rect 24822 18128 24827 18184
rect 22050 18126 24827 18128
rect 12433 18050 12499 18053
rect 7606 18048 12499 18050
rect 7606 17992 12438 18048
rect 12494 17992 12499 18048
rect 7606 17990 12499 17992
rect 12433 17987 12499 17990
rect 15694 17988 15700 18052
rect 15764 18050 15770 18052
rect 18278 18050 18338 18126
rect 21081 18123 21147 18126
rect 24761 18123 24827 18126
rect 18505 18052 18571 18053
rect 18454 18050 18460 18052
rect 15764 17990 18338 18050
rect 18414 17990 18460 18050
rect 18524 18048 18571 18052
rect 18566 17992 18571 18048
rect 15764 17988 15770 17990
rect 18454 17988 18460 17990
rect 18524 17988 18571 17992
rect 18505 17987 18571 17988
rect 19701 18052 19767 18053
rect 19701 18048 19748 18052
rect 19812 18050 19818 18052
rect 24577 18050 24643 18053
rect 24945 18052 25011 18053
rect 24710 18050 24716 18052
rect 19701 17992 19706 18048
rect 19701 17988 19748 17992
rect 19812 17990 19858 18050
rect 24577 18048 24716 18050
rect 24577 17992 24582 18048
rect 24638 17992 24716 18048
rect 24577 17990 24716 17992
rect 19812 17988 19818 17990
rect 19701 17987 19767 17988
rect 24577 17987 24643 17990
rect 24710 17988 24716 17990
rect 24780 17988 24786 18052
rect 24894 18050 24900 18052
rect 24854 17990 24900 18050
rect 24964 18048 25011 18052
rect 25006 17992 25011 18048
rect 24894 17988 24900 17990
rect 24964 17988 25011 17992
rect 24945 17987 25011 17988
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 7782 17852 7788 17916
rect 7852 17914 7858 17916
rect 8569 17914 8635 17917
rect 7852 17912 8635 17914
rect 7852 17856 8574 17912
rect 8630 17856 8635 17912
rect 7852 17854 8635 17856
rect 7852 17852 7858 17854
rect 8569 17851 8635 17854
rect 8886 17852 8892 17916
rect 8956 17914 8962 17916
rect 9397 17914 9463 17917
rect 8956 17912 9463 17914
rect 8956 17856 9402 17912
rect 9458 17856 9463 17912
rect 8956 17854 9463 17856
rect 8956 17852 8962 17854
rect 9397 17851 9463 17854
rect 9673 17914 9739 17917
rect 12157 17914 12223 17917
rect 9673 17912 12223 17914
rect 9673 17856 9678 17912
rect 9734 17856 12162 17912
rect 12218 17856 12223 17912
rect 9673 17854 12223 17856
rect 9673 17851 9739 17854
rect 12157 17851 12223 17854
rect 17166 17852 17172 17916
rect 17236 17914 17242 17916
rect 20529 17914 20595 17917
rect 26200 17914 27000 17944
rect 17236 17912 20595 17914
rect 17236 17856 20534 17912
rect 20590 17856 20595 17912
rect 17236 17854 20595 17856
rect 17236 17852 17242 17854
rect 20529 17851 20595 17854
rect 20670 17854 22800 17914
rect 3969 17778 4035 17781
rect 17217 17778 17283 17781
rect 3969 17776 17283 17778
rect 3969 17720 3974 17776
rect 4030 17720 17222 17776
rect 17278 17720 17283 17776
rect 3969 17718 17283 17720
rect 3969 17715 4035 17718
rect 17217 17715 17283 17718
rect 17677 17778 17743 17781
rect 20670 17778 20730 17854
rect 17677 17776 20730 17778
rect 17677 17720 17682 17776
rect 17738 17720 20730 17776
rect 17677 17718 20730 17720
rect 17677 17715 17743 17718
rect 21950 17716 21956 17780
rect 22020 17778 22026 17780
rect 22134 17778 22140 17780
rect 22020 17718 22140 17778
rect 22020 17716 22026 17718
rect 22134 17716 22140 17718
rect 22204 17716 22210 17780
rect 22740 17778 22800 17854
rect 23430 17854 27000 17914
rect 23430 17778 23490 17854
rect 26200 17824 27000 17854
rect 22740 17718 23490 17778
rect 3417 17642 3483 17645
rect 20989 17642 21055 17645
rect 22829 17642 22895 17645
rect 3417 17640 21055 17642
rect 3417 17584 3422 17640
rect 3478 17584 20994 17640
rect 21050 17584 21055 17640
rect 3417 17582 21055 17584
rect 3417 17579 3483 17582
rect 20989 17579 21055 17582
rect 21222 17640 22895 17642
rect 21222 17584 22834 17640
rect 22890 17584 22895 17640
rect 21222 17582 22895 17584
rect 9121 17506 9187 17509
rect 9438 17506 9444 17508
rect 9121 17504 9444 17506
rect 9121 17448 9126 17504
rect 9182 17448 9444 17504
rect 9121 17446 9444 17448
rect 9121 17443 9187 17446
rect 9438 17444 9444 17446
rect 9508 17444 9514 17508
rect 9857 17506 9923 17509
rect 9990 17506 9996 17508
rect 9857 17504 9996 17506
rect 9857 17448 9862 17504
rect 9918 17448 9996 17504
rect 9857 17446 9996 17448
rect 9857 17443 9923 17446
rect 9990 17444 9996 17446
rect 10060 17444 10066 17508
rect 10777 17506 10843 17509
rect 13721 17506 13787 17509
rect 10777 17504 13787 17506
rect 10777 17448 10782 17504
rect 10838 17448 13726 17504
rect 13782 17448 13787 17504
rect 10777 17446 13787 17448
rect 10777 17443 10843 17446
rect 13721 17443 13787 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 8661 17370 8727 17373
rect 9581 17370 9647 17373
rect 8661 17368 9647 17370
rect 8661 17312 8666 17368
rect 8722 17312 9586 17368
rect 9642 17312 9647 17368
rect 8661 17310 9647 17312
rect 8661 17307 8727 17310
rect 9581 17307 9647 17310
rect 9765 17370 9831 17373
rect 10542 17370 10548 17372
rect 9765 17368 10548 17370
rect 9765 17312 9770 17368
rect 9826 17312 10548 17368
rect 9765 17310 10548 17312
rect 9765 17307 9831 17310
rect 10542 17308 10548 17310
rect 10612 17308 10618 17372
rect 15009 17370 15075 17373
rect 12390 17368 15075 17370
rect 12390 17312 15014 17368
rect 15070 17312 15075 17368
rect 12390 17310 15075 17312
rect 5349 17234 5415 17237
rect 12390 17234 12450 17310
rect 15009 17307 15075 17310
rect 5349 17232 12450 17234
rect 5349 17176 5354 17232
rect 5410 17176 12450 17232
rect 5349 17174 12450 17176
rect 14365 17234 14431 17237
rect 21222 17234 21282 17582
rect 22829 17579 22895 17582
rect 26200 17506 27000 17536
rect 14365 17232 21282 17234
rect 14365 17176 14370 17232
rect 14426 17176 21282 17232
rect 14365 17174 21282 17176
rect 22050 17446 27000 17506
rect 5349 17171 5415 17174
rect 14365 17171 14431 17174
rect 7281 17098 7347 17101
rect 8334 17098 8340 17100
rect 7281 17096 8340 17098
rect 7281 17040 7286 17096
rect 7342 17040 8340 17096
rect 7281 17038 8340 17040
rect 7281 17035 7347 17038
rect 8334 17036 8340 17038
rect 8404 17036 8410 17100
rect 8477 17098 8543 17101
rect 22050 17098 22110 17446
rect 26200 17416 27000 17446
rect 8477 17096 22110 17098
rect 8477 17040 8482 17096
rect 8538 17040 22110 17096
rect 8477 17038 22110 17040
rect 25221 17098 25287 17101
rect 26200 17098 27000 17128
rect 25221 17096 27000 17098
rect 25221 17040 25226 17096
rect 25282 17040 27000 17096
rect 25221 17038 27000 17040
rect 8477 17035 8543 17038
rect 25221 17035 25287 17038
rect 26200 17008 27000 17038
rect 8334 16900 8340 16964
rect 8404 16962 8410 16964
rect 11145 16962 11211 16965
rect 8404 16960 11211 16962
rect 8404 16904 11150 16960
rect 11206 16904 11211 16960
rect 8404 16902 11211 16904
rect 8404 16900 8410 16902
rect 11145 16899 11211 16902
rect 13997 16962 14063 16965
rect 16113 16962 16179 16965
rect 13997 16960 16179 16962
rect 13997 16904 14002 16960
rect 14058 16904 16118 16960
rect 16174 16904 16179 16960
rect 13997 16902 16179 16904
rect 13997 16899 14063 16902
rect 16113 16899 16179 16902
rect 17217 16962 17283 16965
rect 22185 16962 22251 16965
rect 17217 16960 22251 16962
rect 17217 16904 17222 16960
rect 17278 16904 22190 16960
rect 22246 16904 22251 16960
rect 17217 16902 22251 16904
rect 17217 16899 17283 16902
rect 22185 16899 22251 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 8477 16826 8543 16829
rect 10869 16826 10935 16829
rect 12525 16826 12591 16829
rect 15929 16826 15995 16829
rect 3374 16824 8543 16826
rect 3374 16768 8482 16824
rect 8538 16768 8543 16824
rect 3374 16766 8543 16768
rect 2865 16690 2931 16693
rect 3374 16690 3434 16766
rect 8477 16763 8543 16766
rect 8664 16766 9506 16826
rect 2865 16688 3434 16690
rect 2865 16632 2870 16688
rect 2926 16632 3434 16688
rect 2865 16630 3434 16632
rect 7649 16690 7715 16693
rect 8664 16690 8724 16766
rect 9446 16690 9506 16766
rect 10869 16824 12591 16826
rect 10869 16768 10874 16824
rect 10930 16768 12530 16824
rect 12586 16768 12591 16824
rect 10869 16766 12591 16768
rect 10869 16763 10935 16766
rect 12525 16763 12591 16766
rect 13494 16824 15995 16826
rect 13494 16768 15934 16824
rect 15990 16768 15995 16824
rect 13494 16766 15995 16768
rect 10225 16690 10291 16693
rect 7649 16688 8724 16690
rect 7649 16632 7654 16688
rect 7710 16632 8724 16688
rect 7649 16630 8724 16632
rect 8894 16630 9322 16690
rect 9446 16688 10291 16690
rect 9446 16632 10230 16688
rect 10286 16632 10291 16688
rect 9446 16630 10291 16632
rect 2865 16627 2931 16630
rect 7649 16627 7715 16630
rect 4613 16554 4679 16557
rect 8894 16554 8954 16630
rect 4613 16552 8954 16554
rect 4613 16496 4618 16552
rect 4674 16496 8954 16552
rect 4613 16494 8954 16496
rect 9262 16554 9322 16630
rect 10225 16627 10291 16630
rect 10726 16628 10732 16692
rect 10796 16690 10802 16692
rect 11881 16690 11947 16693
rect 10796 16688 11947 16690
rect 10796 16632 11886 16688
rect 11942 16632 11947 16688
rect 10796 16630 11947 16632
rect 10796 16628 10802 16630
rect 11881 16627 11947 16630
rect 12525 16690 12591 16693
rect 13494 16690 13554 16766
rect 15929 16763 15995 16766
rect 16481 16826 16547 16829
rect 17953 16826 18019 16829
rect 16481 16824 18019 16826
rect 16481 16768 16486 16824
rect 16542 16768 17958 16824
rect 18014 16768 18019 16824
rect 16481 16766 18019 16768
rect 16481 16763 16547 16766
rect 17953 16763 18019 16766
rect 20713 16826 20779 16829
rect 22318 16826 22324 16828
rect 20713 16824 22324 16826
rect 20713 16768 20718 16824
rect 20774 16768 22324 16824
rect 20713 16766 22324 16768
rect 20713 16763 20779 16766
rect 22318 16764 22324 16766
rect 22388 16764 22394 16828
rect 23657 16826 23723 16829
rect 25589 16826 25655 16829
rect 23657 16824 25655 16826
rect 23657 16768 23662 16824
rect 23718 16768 25594 16824
rect 25650 16768 25655 16824
rect 23657 16766 25655 16768
rect 23657 16763 23723 16766
rect 25589 16763 25655 16766
rect 15510 16690 15516 16692
rect 12525 16688 13554 16690
rect 12525 16632 12530 16688
rect 12586 16632 13554 16688
rect 12525 16630 13554 16632
rect 13678 16630 15516 16690
rect 12525 16627 12591 16630
rect 10174 16554 10180 16556
rect 9262 16494 10180 16554
rect 4613 16491 4679 16494
rect 10174 16492 10180 16494
rect 10244 16492 10250 16556
rect 12433 16554 12499 16557
rect 13678 16554 13738 16630
rect 15510 16628 15516 16630
rect 15580 16628 15586 16692
rect 15653 16690 15719 16693
rect 16941 16690 17007 16693
rect 15653 16688 17007 16690
rect 15653 16632 15658 16688
rect 15714 16632 16946 16688
rect 17002 16632 17007 16688
rect 15653 16630 17007 16632
rect 15653 16627 15719 16630
rect 16941 16627 17007 16630
rect 17585 16690 17651 16693
rect 17718 16690 17724 16692
rect 17585 16688 17724 16690
rect 17585 16632 17590 16688
rect 17646 16632 17724 16688
rect 17585 16630 17724 16632
rect 17585 16627 17651 16630
rect 17718 16628 17724 16630
rect 17788 16628 17794 16692
rect 23197 16690 23263 16693
rect 26200 16690 27000 16720
rect 23197 16688 27000 16690
rect 23197 16632 23202 16688
rect 23258 16632 27000 16688
rect 23197 16630 27000 16632
rect 23197 16627 23263 16630
rect 26200 16600 27000 16630
rect 12433 16552 13738 16554
rect 12433 16496 12438 16552
rect 12494 16496 13738 16552
rect 12433 16494 13738 16496
rect 12433 16491 12499 16494
rect 14590 16492 14596 16556
rect 14660 16554 14666 16556
rect 16389 16554 16455 16557
rect 14660 16552 16455 16554
rect 14660 16496 16394 16552
rect 16450 16496 16455 16552
rect 14660 16494 16455 16496
rect 14660 16492 14666 16494
rect 16389 16491 16455 16494
rect 19190 16492 19196 16556
rect 19260 16554 19266 16556
rect 20294 16554 20300 16556
rect 19260 16494 20300 16554
rect 19260 16492 19266 16494
rect 20294 16492 20300 16494
rect 20364 16492 20370 16556
rect 9397 16418 9463 16421
rect 13445 16418 13511 16421
rect 9397 16416 13511 16418
rect 9397 16360 9402 16416
rect 9458 16360 13450 16416
rect 13506 16360 13511 16416
rect 9397 16358 13511 16360
rect 9397 16355 9463 16358
rect 13445 16355 13511 16358
rect 18822 16356 18828 16420
rect 18892 16418 18898 16420
rect 22093 16418 22159 16421
rect 18892 16416 22159 16418
rect 18892 16360 22098 16416
rect 22154 16360 22159 16416
rect 18892 16358 22159 16360
rect 18892 16356 18898 16358
rect 22093 16355 22159 16358
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 8661 16282 8727 16285
rect 11145 16282 11211 16285
rect 8661 16280 11211 16282
rect 8661 16224 8666 16280
rect 8722 16224 11150 16280
rect 11206 16224 11211 16280
rect 8661 16222 11211 16224
rect 8661 16219 8727 16222
rect 11145 16219 11211 16222
rect 14089 16282 14155 16285
rect 17033 16282 17099 16285
rect 14089 16280 17099 16282
rect 14089 16224 14094 16280
rect 14150 16224 17038 16280
rect 17094 16224 17099 16280
rect 14089 16222 17099 16224
rect 14089 16219 14155 16222
rect 17033 16219 17099 16222
rect 22001 16282 22067 16285
rect 26200 16282 27000 16312
rect 22001 16280 27000 16282
rect 22001 16224 22006 16280
rect 22062 16224 27000 16280
rect 22001 16222 27000 16224
rect 22001 16219 22067 16222
rect 26200 16192 27000 16222
rect 6545 16146 6611 16149
rect 6545 16144 8908 16146
rect 6545 16088 6550 16144
rect 6606 16112 8908 16144
rect 6606 16088 9322 16112
rect 6545 16086 9322 16088
rect 6545 16083 6611 16086
rect 8848 16052 9322 16086
rect 9438 16084 9444 16148
rect 9508 16146 9514 16148
rect 9508 16086 24226 16146
rect 9508 16084 9514 16086
rect 9262 16010 9322 16052
rect 12525 16010 12591 16013
rect 9262 16008 12591 16010
rect 9262 15952 12530 16008
rect 12586 15952 12591 16008
rect 9262 15950 12591 15952
rect 12525 15947 12591 15950
rect 12750 15948 12756 16012
rect 12820 16010 12826 16012
rect 14038 16010 14044 16012
rect 12820 15950 14044 16010
rect 12820 15948 12826 15950
rect 14038 15948 14044 15950
rect 14108 15948 14114 16012
rect 14222 15948 14228 16012
rect 14292 16010 14298 16012
rect 16246 16010 16252 16012
rect 14292 15950 16252 16010
rect 14292 15948 14298 15950
rect 16246 15948 16252 15950
rect 16316 15948 16322 16012
rect 18413 16010 18479 16013
rect 16392 16008 18479 16010
rect 16392 15952 18418 16008
rect 18474 15952 18479 16008
rect 16392 15950 18479 15952
rect 3969 15874 4035 15877
rect 9806 15874 9812 15876
rect 3969 15872 9812 15874
rect 3969 15816 3974 15872
rect 4030 15816 9812 15872
rect 3969 15814 9812 15816
rect 3969 15811 4035 15814
rect 9806 15812 9812 15814
rect 9876 15812 9882 15876
rect 9949 15874 10015 15877
rect 12249 15874 12315 15877
rect 9949 15872 12315 15874
rect 9949 15816 9954 15872
rect 10010 15816 12254 15872
rect 12310 15816 12315 15872
rect 9949 15814 12315 15816
rect 9949 15811 10015 15814
rect 12249 15811 12315 15814
rect 14089 15874 14155 15877
rect 16392 15874 16452 15950
rect 18413 15947 18479 15950
rect 22093 16010 22159 16013
rect 23422 16010 23428 16012
rect 22093 16008 23428 16010
rect 22093 15952 22098 16008
rect 22154 15952 23428 16008
rect 22093 15950 23428 15952
rect 22093 15947 22159 15950
rect 23422 15948 23428 15950
rect 23492 15948 23498 16012
rect 14089 15872 16452 15874
rect 14089 15816 14094 15872
rect 14150 15816 16452 15872
rect 14089 15814 16452 15816
rect 16941 15874 17007 15877
rect 21909 15874 21975 15877
rect 16941 15872 21975 15874
rect 16941 15816 16946 15872
rect 17002 15816 21914 15872
rect 21970 15816 21975 15872
rect 16941 15814 21975 15816
rect 24166 15874 24226 16086
rect 26200 15874 27000 15904
rect 24166 15814 27000 15874
rect 14089 15811 14155 15814
rect 16941 15811 17007 15814
rect 21909 15811 21975 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 26200 15784 27000 15814
rect 22946 15743 23262 15744
rect 8845 15738 8911 15741
rect 12341 15738 12407 15741
rect 13813 15740 13879 15741
rect 16573 15740 16639 15741
rect 13813 15738 13860 15740
rect 8845 15736 12407 15738
rect 8845 15680 8850 15736
rect 8906 15680 12346 15736
rect 12402 15680 12407 15736
rect 8845 15678 12407 15680
rect 13768 15736 13860 15738
rect 13768 15680 13818 15736
rect 13768 15678 13860 15680
rect 8845 15675 8911 15678
rect 12341 15675 12407 15678
rect 13813 15676 13860 15678
rect 13924 15676 13930 15740
rect 16246 15676 16252 15740
rect 16316 15738 16322 15740
rect 16573 15738 16620 15740
rect 16316 15736 16620 15738
rect 16316 15680 16578 15736
rect 16316 15678 16620 15680
rect 16316 15676 16322 15678
rect 16573 15676 16620 15678
rect 16684 15676 16690 15740
rect 19006 15738 19012 15740
rect 16760 15678 19012 15738
rect 13813 15675 13879 15676
rect 16573 15675 16639 15676
rect 5758 15540 5764 15604
rect 5828 15602 5834 15604
rect 12433 15602 12499 15605
rect 5828 15600 12499 15602
rect 5828 15544 12438 15600
rect 12494 15544 12499 15600
rect 5828 15542 12499 15544
rect 5828 15540 5834 15542
rect 12433 15539 12499 15542
rect 15837 15602 15903 15605
rect 16760 15602 16820 15678
rect 19006 15676 19012 15678
rect 19076 15676 19082 15740
rect 20846 15676 20852 15740
rect 20916 15738 20922 15740
rect 22001 15738 22067 15741
rect 20916 15736 22067 15738
rect 20916 15680 22006 15736
rect 22062 15680 22067 15736
rect 20916 15678 22067 15680
rect 20916 15676 20922 15678
rect 22001 15675 22067 15678
rect 23974 15676 23980 15740
rect 24044 15738 24050 15740
rect 25773 15738 25839 15741
rect 24044 15736 25839 15738
rect 24044 15680 25778 15736
rect 25834 15680 25839 15736
rect 24044 15678 25839 15680
rect 24044 15676 24050 15678
rect 25773 15675 25839 15678
rect 15837 15600 16820 15602
rect 15837 15544 15842 15600
rect 15898 15544 16820 15600
rect 15837 15542 16820 15544
rect 17217 15602 17283 15605
rect 25221 15602 25287 15605
rect 17217 15600 25287 15602
rect 17217 15544 17222 15600
rect 17278 15544 25226 15600
rect 25282 15544 25287 15600
rect 17217 15542 25287 15544
rect 15837 15539 15903 15542
rect 17217 15539 17283 15542
rect 25221 15539 25287 15542
rect 1209 15466 1275 15469
rect 7833 15466 7899 15469
rect 9121 15468 9187 15469
rect 9489 15468 9555 15469
rect 1209 15464 7899 15466
rect 1209 15408 1214 15464
rect 1270 15408 7838 15464
rect 7894 15408 7899 15464
rect 1209 15406 7899 15408
rect 1209 15403 1275 15406
rect 7833 15403 7899 15406
rect 9070 15404 9076 15468
rect 9140 15466 9187 15468
rect 9140 15464 9232 15466
rect 9182 15408 9232 15464
rect 9140 15406 9232 15408
rect 9140 15404 9187 15406
rect 9438 15404 9444 15468
rect 9508 15466 9555 15468
rect 9673 15466 9739 15469
rect 19425 15466 19491 15469
rect 9508 15464 9600 15466
rect 9550 15408 9600 15464
rect 9508 15406 9600 15408
rect 9673 15464 19491 15466
rect 9673 15408 9678 15464
rect 9734 15408 19430 15464
rect 19486 15408 19491 15464
rect 9673 15406 19491 15408
rect 9508 15404 9555 15406
rect 9121 15403 9187 15404
rect 9489 15403 9555 15404
rect 9673 15403 9739 15406
rect 19425 15403 19491 15406
rect 20662 15404 20668 15468
rect 20732 15466 20738 15468
rect 23422 15466 23428 15468
rect 20732 15406 23428 15466
rect 20732 15404 20738 15406
rect 23422 15404 23428 15406
rect 23492 15404 23498 15468
rect 25773 15466 25839 15469
rect 26200 15466 27000 15496
rect 25773 15464 27000 15466
rect 25773 15408 25778 15464
rect 25834 15408 27000 15464
rect 25773 15406 27000 15408
rect 25773 15403 25839 15406
rect 26200 15376 27000 15406
rect 473 15330 539 15333
rect 1393 15330 1459 15333
rect 473 15328 1459 15330
rect 473 15272 478 15328
rect 534 15272 1398 15328
rect 1454 15272 1459 15328
rect 473 15270 1459 15272
rect 473 15267 539 15270
rect 1393 15267 1459 15270
rect 9806 15268 9812 15332
rect 9876 15330 9882 15332
rect 10777 15330 10843 15333
rect 11237 15332 11303 15333
rect 11237 15330 11284 15332
rect 9876 15328 10843 15330
rect 9876 15272 10782 15328
rect 10838 15272 10843 15328
rect 9876 15270 10843 15272
rect 11192 15328 11284 15330
rect 11192 15272 11242 15328
rect 11192 15270 11284 15272
rect 9876 15268 9882 15270
rect 10777 15267 10843 15270
rect 11237 15268 11284 15270
rect 11348 15268 11354 15332
rect 11697 15330 11763 15333
rect 12014 15330 12020 15332
rect 11697 15328 12020 15330
rect 11697 15272 11702 15328
rect 11758 15272 12020 15328
rect 11697 15270 12020 15272
rect 11237 15267 11303 15268
rect 11697 15267 11763 15270
rect 12014 15268 12020 15270
rect 12084 15268 12090 15332
rect 12341 15330 12407 15333
rect 15929 15330 15995 15333
rect 12341 15328 15995 15330
rect 12341 15272 12346 15328
rect 12402 15272 15934 15328
rect 15990 15272 15995 15328
rect 12341 15270 15995 15272
rect 12341 15267 12407 15270
rect 15929 15267 15995 15270
rect 19609 15330 19675 15333
rect 20662 15330 20668 15332
rect 19609 15328 20668 15330
rect 19609 15272 19614 15328
rect 19670 15272 20668 15328
rect 19609 15270 20668 15272
rect 19609 15267 19675 15270
rect 20662 15268 20668 15270
rect 20732 15268 20738 15332
rect 22134 15268 22140 15332
rect 22204 15330 22210 15332
rect 23381 15330 23447 15333
rect 22204 15328 23447 15330
rect 22204 15272 23386 15328
rect 23442 15272 23447 15328
rect 22204 15270 23447 15272
rect 22204 15268 22210 15270
rect 23381 15267 23447 15270
rect 25078 15268 25084 15332
rect 25148 15330 25154 15332
rect 25221 15330 25287 15333
rect 25148 15328 25287 15330
rect 25148 15272 25226 15328
rect 25282 15272 25287 15328
rect 25148 15270 25287 15272
rect 25148 15268 25154 15270
rect 25221 15267 25287 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 4429 15194 4495 15197
rect 5022 15194 5028 15196
rect 4429 15192 5028 15194
rect 4429 15136 4434 15192
rect 4490 15136 5028 15192
rect 4429 15134 5028 15136
rect 4429 15131 4495 15134
rect 5022 15132 5028 15134
rect 5092 15132 5098 15196
rect 10910 15132 10916 15196
rect 10980 15194 10986 15196
rect 16113 15194 16179 15197
rect 10980 15192 16179 15194
rect 10980 15136 16118 15192
rect 16174 15136 16179 15192
rect 10980 15134 16179 15136
rect 10980 15132 10986 15134
rect 16113 15131 16179 15134
rect 18638 15132 18644 15196
rect 18708 15194 18714 15196
rect 19241 15194 19307 15197
rect 18708 15192 19307 15194
rect 18708 15136 19246 15192
rect 19302 15136 19307 15192
rect 18708 15134 19307 15136
rect 18708 15132 18714 15134
rect 19241 15131 19307 15134
rect 21449 15194 21515 15197
rect 23565 15194 23631 15197
rect 21449 15192 23631 15194
rect 21449 15136 21454 15192
rect 21510 15136 23570 15192
rect 23626 15136 23631 15192
rect 21449 15134 23631 15136
rect 21449 15131 21515 15134
rect 23565 15131 23631 15134
rect 24117 15194 24183 15197
rect 25998 15194 26004 15196
rect 24117 15192 26004 15194
rect 24117 15136 24122 15192
rect 24178 15136 26004 15192
rect 24117 15134 26004 15136
rect 24117 15131 24183 15134
rect 25998 15132 26004 15134
rect 26068 15132 26074 15196
rect 2589 15058 2655 15061
rect 8334 15058 8340 15060
rect 2589 15056 8340 15058
rect 2589 15000 2594 15056
rect 2650 15000 8340 15056
rect 2589 14998 8340 15000
rect 2589 14995 2655 14998
rect 8334 14996 8340 14998
rect 8404 14996 8410 15060
rect 10133 15058 10199 15061
rect 14641 15058 14707 15061
rect 10133 15056 14707 15058
rect 10133 15000 10138 15056
rect 10194 15000 14646 15056
rect 14702 15000 14707 15056
rect 10133 14998 14707 15000
rect 10133 14995 10199 14998
rect 14641 14995 14707 14998
rect 15510 14996 15516 15060
rect 15580 15058 15586 15060
rect 16798 15058 16804 15060
rect 15580 14998 16804 15058
rect 15580 14996 15586 14998
rect 16798 14996 16804 14998
rect 16868 14996 16874 15060
rect 17953 15058 18019 15061
rect 18822 15058 18828 15060
rect 17953 15056 18828 15058
rect 17953 15000 17958 15056
rect 18014 15000 18828 15056
rect 17953 14998 18828 15000
rect 17953 14995 18019 14998
rect 18822 14996 18828 14998
rect 18892 14996 18898 15060
rect 22645 15058 22711 15061
rect 26200 15058 27000 15088
rect 22645 15056 27000 15058
rect 22645 15000 22650 15056
rect 22706 15000 27000 15056
rect 22645 14998 27000 15000
rect 22645 14995 22711 14998
rect 26200 14968 27000 14998
rect 4705 14922 4771 14925
rect 15142 14922 15148 14924
rect 4705 14920 15148 14922
rect 4705 14864 4710 14920
rect 4766 14864 15148 14920
rect 4705 14862 15148 14864
rect 4705 14859 4771 14862
rect 15142 14860 15148 14862
rect 15212 14860 15218 14924
rect 20713 14922 20779 14925
rect 15288 14920 20779 14922
rect 15288 14864 20718 14920
rect 20774 14864 20779 14920
rect 15288 14862 20779 14864
rect 3785 14786 3851 14789
rect 12249 14786 12315 14789
rect 3785 14784 12315 14786
rect 3785 14728 3790 14784
rect 3846 14728 12254 14784
rect 12310 14728 12315 14784
rect 3785 14726 12315 14728
rect 3785 14723 3851 14726
rect 12249 14723 12315 14726
rect 14365 14786 14431 14789
rect 15288 14786 15348 14862
rect 20713 14859 20779 14862
rect 21909 14922 21975 14925
rect 24761 14922 24827 14925
rect 25078 14922 25084 14924
rect 21909 14920 24226 14922
rect 21909 14864 21914 14920
rect 21970 14864 24226 14920
rect 21909 14862 24226 14864
rect 21909 14859 21975 14862
rect 14365 14784 15348 14786
rect 14365 14728 14370 14784
rect 14426 14728 15348 14784
rect 14365 14726 15348 14728
rect 14365 14723 14431 14726
rect 17534 14724 17540 14788
rect 17604 14786 17610 14788
rect 21541 14786 21607 14789
rect 17604 14784 21607 14786
rect 17604 14728 21546 14784
rect 21602 14728 21607 14784
rect 17604 14726 21607 14728
rect 17604 14724 17610 14726
rect 21541 14723 21607 14726
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 9029 14650 9095 14653
rect 9029 14648 12450 14650
rect 9029 14592 9034 14648
rect 9090 14592 12450 14648
rect 9029 14590 12450 14592
rect 9029 14587 9095 14590
rect 6361 14514 6427 14517
rect 10961 14514 11027 14517
rect 11513 14516 11579 14517
rect 11462 14514 11468 14516
rect 6361 14512 11027 14514
rect 6361 14456 6366 14512
rect 6422 14456 10966 14512
rect 11022 14456 11027 14512
rect 6361 14454 11027 14456
rect 11422 14454 11468 14514
rect 11532 14512 11579 14516
rect 11574 14456 11579 14512
rect 6361 14451 6427 14454
rect 10961 14451 11027 14454
rect 11462 14452 11468 14454
rect 11532 14452 11579 14456
rect 12390 14514 12450 14590
rect 14406 14588 14412 14652
rect 14476 14650 14482 14652
rect 16430 14650 16436 14652
rect 14476 14590 16436 14650
rect 14476 14588 14482 14590
rect 16430 14588 16436 14590
rect 16500 14588 16506 14652
rect 16665 14650 16731 14653
rect 20345 14650 20411 14653
rect 21817 14652 21883 14653
rect 21766 14650 21772 14652
rect 16665 14648 20411 14650
rect 16665 14592 16670 14648
rect 16726 14592 20350 14648
rect 20406 14592 20411 14648
rect 16665 14590 20411 14592
rect 21726 14590 21772 14650
rect 21836 14648 21883 14652
rect 21878 14592 21883 14648
rect 16665 14587 16731 14590
rect 20345 14587 20411 14590
rect 21766 14588 21772 14590
rect 21836 14588 21883 14592
rect 24166 14650 24226 14862
rect 24761 14920 25084 14922
rect 24761 14864 24766 14920
rect 24822 14864 25084 14920
rect 24761 14862 25084 14864
rect 24761 14859 24827 14862
rect 25078 14860 25084 14862
rect 25148 14860 25154 14924
rect 26200 14650 27000 14680
rect 24166 14590 27000 14650
rect 21817 14587 21883 14588
rect 26200 14560 27000 14590
rect 17166 14514 17172 14516
rect 12390 14454 17172 14514
rect 17166 14452 17172 14454
rect 17236 14452 17242 14516
rect 17585 14514 17651 14517
rect 17769 14514 17835 14517
rect 17585 14512 17835 14514
rect 17585 14456 17590 14512
rect 17646 14456 17774 14512
rect 17830 14456 17835 14512
rect 17585 14454 17835 14456
rect 11513 14451 11579 14452
rect 17585 14451 17651 14454
rect 17769 14451 17835 14454
rect 19374 14452 19380 14516
rect 19444 14514 19450 14516
rect 23657 14514 23723 14517
rect 24342 14514 24348 14516
rect 19444 14454 22156 14514
rect 19444 14452 19450 14454
rect 3969 14378 4035 14381
rect 14457 14378 14523 14381
rect 3969 14376 14523 14378
rect 3969 14320 3974 14376
rect 4030 14320 14462 14376
rect 14518 14320 14523 14376
rect 3969 14318 14523 14320
rect 3969 14315 4035 14318
rect 14457 14315 14523 14318
rect 17585 14378 17651 14381
rect 21950 14378 21956 14380
rect 17585 14376 21956 14378
rect 17585 14320 17590 14376
rect 17646 14320 21956 14376
rect 17585 14318 21956 14320
rect 17585 14315 17651 14318
rect 21950 14316 21956 14318
rect 22020 14316 22026 14380
rect 22096 14378 22156 14454
rect 23657 14512 24348 14514
rect 23657 14456 23662 14512
rect 23718 14456 24348 14512
rect 23657 14454 24348 14456
rect 23657 14451 23723 14454
rect 24342 14452 24348 14454
rect 24412 14452 24418 14516
rect 26049 14378 26115 14381
rect 22096 14376 26115 14378
rect 22096 14320 26054 14376
rect 26110 14320 26115 14376
rect 22096 14318 26115 14320
rect 26049 14315 26115 14318
rect 11329 14242 11395 14245
rect 13486 14242 13492 14244
rect 11329 14240 13492 14242
rect 11329 14184 11334 14240
rect 11390 14184 13492 14240
rect 11329 14182 13492 14184
rect 11329 14179 11395 14182
rect 13486 14180 13492 14182
rect 13556 14180 13562 14244
rect 19006 14180 19012 14244
rect 19076 14242 19082 14244
rect 20437 14242 20503 14245
rect 19076 14240 20503 14242
rect 19076 14184 20442 14240
rect 20498 14184 20503 14240
rect 19076 14182 20503 14184
rect 19076 14180 19082 14182
rect 20437 14179 20503 14182
rect 26049 14242 26115 14245
rect 26200 14242 27000 14272
rect 26049 14240 27000 14242
rect 26049 14184 26054 14240
rect 26110 14184 27000 14240
rect 26049 14182 27000 14184
rect 26049 14179 26115 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 26200 14152 27000 14182
rect 17946 14111 18262 14112
rect 11697 14106 11763 14109
rect 8342 14104 11763 14106
rect 8342 14048 11702 14104
rect 11758 14048 11763 14104
rect 8342 14046 11763 14048
rect 4102 13908 4108 13972
rect 4172 13970 4178 13972
rect 8342 13970 8402 14046
rect 11697 14043 11763 14046
rect 11881 14106 11947 14109
rect 16665 14106 16731 14109
rect 19558 14106 19564 14108
rect 11881 14104 16731 14106
rect 11881 14048 11886 14104
rect 11942 14048 16670 14104
rect 16726 14048 16731 14104
rect 11881 14046 16731 14048
rect 11881 14043 11947 14046
rect 16665 14043 16731 14046
rect 18462 14046 19564 14106
rect 4172 13910 8402 13970
rect 11237 13970 11303 13973
rect 11646 13970 11652 13972
rect 11237 13968 11652 13970
rect 11237 13912 11242 13968
rect 11298 13912 11652 13968
rect 11237 13910 11652 13912
rect 4172 13908 4178 13910
rect 11237 13907 11303 13910
rect 11646 13908 11652 13910
rect 11716 13908 11722 13972
rect 18462 13970 18522 14046
rect 19558 14044 19564 14046
rect 19628 14044 19634 14108
rect 20437 14106 20503 14109
rect 23013 14106 23079 14109
rect 20437 14104 23079 14106
rect 20437 14048 20442 14104
rect 20498 14048 23018 14104
rect 23074 14048 23079 14104
rect 20437 14046 23079 14048
rect 20437 14043 20503 14046
rect 23013 14043 23079 14046
rect 15702 13910 18522 13970
rect 22737 13970 22803 13973
rect 22737 13968 26066 13970
rect 22737 13912 22742 13968
rect 22798 13912 26066 13968
rect 22737 13910 26066 13912
rect 8293 13834 8359 13837
rect 12801 13834 12867 13837
rect 15702 13834 15762 13910
rect 22737 13907 22803 13910
rect 8293 13832 15762 13834
rect 8293 13776 8298 13832
rect 8354 13776 12806 13832
rect 12862 13776 15762 13832
rect 8293 13774 15762 13776
rect 8293 13771 8359 13774
rect 12801 13771 12867 13774
rect 16614 13772 16620 13836
rect 16684 13834 16690 13836
rect 21725 13834 21791 13837
rect 22369 13836 22435 13837
rect 22318 13834 22324 13836
rect 16684 13832 21791 13834
rect 16684 13776 21730 13832
rect 21786 13776 21791 13832
rect 16684 13774 21791 13776
rect 22278 13774 22324 13834
rect 22388 13832 22435 13836
rect 22430 13776 22435 13832
rect 16684 13772 16690 13774
rect 21725 13771 21791 13774
rect 22318 13772 22324 13774
rect 22388 13772 22435 13776
rect 22369 13771 22435 13772
rect 25589 13834 25655 13837
rect 25814 13834 25820 13836
rect 25589 13832 25820 13834
rect 25589 13776 25594 13832
rect 25650 13776 25820 13832
rect 25589 13774 25820 13776
rect 25589 13771 25655 13774
rect 25814 13772 25820 13774
rect 25884 13772 25890 13836
rect 26006 13834 26066 13910
rect 26200 13834 27000 13864
rect 26006 13774 27000 13834
rect 26200 13744 27000 13774
rect 10409 13698 10475 13701
rect 12249 13698 12315 13701
rect 10409 13696 12315 13698
rect 10409 13640 10414 13696
rect 10470 13640 12254 13696
rect 12310 13640 12315 13696
rect 10409 13638 12315 13640
rect 10409 13635 10475 13638
rect 12249 13635 12315 13638
rect 17217 13698 17283 13701
rect 19926 13698 19932 13700
rect 17217 13696 19932 13698
rect 17217 13640 17222 13696
rect 17278 13640 19932 13696
rect 17217 13638 19932 13640
rect 17217 13635 17283 13638
rect 19926 13636 19932 13638
rect 19996 13636 20002 13700
rect 20110 13636 20116 13700
rect 20180 13698 20186 13700
rect 20805 13698 20871 13701
rect 20180 13696 20871 13698
rect 20180 13640 20810 13696
rect 20866 13640 20871 13696
rect 20180 13638 20871 13640
rect 20180 13636 20186 13638
rect 20805 13635 20871 13638
rect 21214 13636 21220 13700
rect 21284 13698 21290 13700
rect 21357 13698 21423 13701
rect 21284 13696 21423 13698
rect 21284 13640 21362 13696
rect 21418 13640 21423 13696
rect 21284 13638 21423 13640
rect 21284 13636 21290 13638
rect 21357 13635 21423 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 5809 13562 5875 13565
rect 8886 13562 8892 13564
rect 5809 13560 8892 13562
rect 5809 13504 5814 13560
rect 5870 13504 8892 13560
rect 5809 13502 8892 13504
rect 5809 13499 5875 13502
rect 8886 13500 8892 13502
rect 8956 13500 8962 13564
rect 9213 13562 9279 13565
rect 9622 13562 9628 13564
rect 9213 13560 9628 13562
rect 9213 13504 9218 13560
rect 9274 13504 9628 13560
rect 9213 13502 9628 13504
rect 9213 13499 9279 13502
rect 9622 13500 9628 13502
rect 9692 13500 9698 13564
rect 13353 13562 13419 13565
rect 16113 13562 16179 13565
rect 20253 13562 20319 13565
rect 13353 13560 15992 13562
rect 13353 13504 13358 13560
rect 13414 13504 15992 13560
rect 13353 13502 15992 13504
rect 13353 13499 13419 13502
rect 7281 13426 7347 13429
rect 9489 13426 9555 13429
rect 7281 13424 9555 13426
rect 7281 13368 7286 13424
rect 7342 13368 9494 13424
rect 9550 13368 9555 13424
rect 7281 13366 9555 13368
rect 7281 13363 7347 13366
rect 9489 13363 9555 13366
rect 10133 13426 10199 13429
rect 15932 13426 15992 13502
rect 16113 13560 20319 13562
rect 16113 13504 16118 13560
rect 16174 13504 20258 13560
rect 20314 13504 20319 13560
rect 16113 13502 20319 13504
rect 16113 13499 16179 13502
rect 20253 13499 20319 13502
rect 21582 13426 21588 13428
rect 10133 13424 15762 13426
rect 10133 13368 10138 13424
rect 10194 13368 15762 13424
rect 10133 13366 15762 13368
rect 15932 13366 21588 13426
rect 10133 13363 10199 13366
rect 3233 13290 3299 13293
rect 15469 13290 15535 13293
rect 3233 13288 15535 13290
rect 3233 13232 3238 13288
rect 3294 13232 15474 13288
rect 15530 13232 15535 13288
rect 3233 13230 15535 13232
rect 15702 13290 15762 13366
rect 21582 13364 21588 13366
rect 21652 13426 21658 13428
rect 21725 13426 21791 13429
rect 21652 13424 21791 13426
rect 21652 13368 21730 13424
rect 21786 13368 21791 13424
rect 21652 13366 21791 13368
rect 21652 13364 21658 13366
rect 21725 13363 21791 13366
rect 22921 13426 22987 13429
rect 26200 13426 27000 13456
rect 22921 13424 27000 13426
rect 22921 13368 22926 13424
rect 22982 13368 27000 13424
rect 22921 13366 27000 13368
rect 22921 13363 22987 13366
rect 26200 13336 27000 13366
rect 16614 13290 16620 13292
rect 15702 13230 16620 13290
rect 3233 13227 3299 13230
rect 15469 13227 15535 13230
rect 16614 13228 16620 13230
rect 16684 13228 16690 13292
rect 19517 13290 19583 13293
rect 20478 13290 20484 13292
rect 19517 13288 20484 13290
rect 19517 13232 19522 13288
rect 19578 13232 20484 13288
rect 19517 13230 20484 13232
rect 19517 13227 19583 13230
rect 20478 13228 20484 13230
rect 20548 13228 20554 13292
rect 23013 13290 23079 13293
rect 23606 13290 23612 13292
rect 23013 13288 23612 13290
rect 23013 13232 23018 13288
rect 23074 13232 23612 13288
rect 23013 13230 23612 13232
rect 23013 13227 23079 13230
rect 23606 13228 23612 13230
rect 23676 13228 23682 13292
rect 10593 13154 10659 13157
rect 14273 13154 14339 13157
rect 10593 13152 14339 13154
rect 10593 13096 10598 13152
rect 10654 13096 14278 13152
rect 14334 13096 14339 13152
rect 10593 13094 14339 13096
rect 10593 13091 10659 13094
rect 14273 13091 14339 13094
rect 15193 13154 15259 13157
rect 16113 13154 16179 13157
rect 16389 13154 16455 13157
rect 15193 13152 16179 13154
rect 15193 13096 15198 13152
rect 15254 13096 16118 13152
rect 16174 13096 16179 13152
rect 15193 13094 16179 13096
rect 15193 13091 15259 13094
rect 16113 13091 16179 13094
rect 16254 13152 16455 13154
rect 16254 13096 16394 13152
rect 16450 13096 16455 13152
rect 16254 13094 16455 13096
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 6913 13020 6979 13021
rect 6862 13018 6868 13020
rect 6822 12958 6868 13018
rect 6932 13016 6979 13020
rect 6974 12960 6979 13016
rect 6862 12956 6868 12958
rect 6932 12956 6979 12960
rect 6913 12955 6979 12956
rect 8569 13018 8635 13021
rect 13077 13018 13143 13021
rect 16254 13018 16314 13094
rect 16389 13091 16455 13094
rect 19425 13154 19491 13157
rect 20253 13154 20319 13157
rect 19425 13152 20319 13154
rect 19425 13096 19430 13152
rect 19486 13096 20258 13152
rect 20314 13096 20319 13152
rect 19425 13094 20319 13096
rect 19425 13091 19491 13094
rect 20253 13091 20319 13094
rect 21265 13154 21331 13157
rect 21449 13154 21515 13157
rect 21265 13152 21515 13154
rect 21265 13096 21270 13152
rect 21326 13096 21454 13152
rect 21510 13096 21515 13152
rect 21265 13094 21515 13096
rect 21265 13091 21331 13094
rect 21449 13091 21515 13094
rect 22001 13154 22067 13157
rect 23790 13154 23796 13156
rect 22001 13152 23796 13154
rect 22001 13096 22006 13152
rect 22062 13096 23796 13152
rect 22001 13094 23796 13096
rect 22001 13091 22067 13094
rect 23790 13092 23796 13094
rect 23860 13092 23866 13156
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 8569 13016 12772 13018
rect 8569 12960 8574 13016
rect 8630 12960 12772 13016
rect 8569 12958 12772 12960
rect 8569 12955 8635 12958
rect 2446 12820 2452 12884
rect 2516 12882 2522 12884
rect 2865 12882 2931 12885
rect 2516 12880 2931 12882
rect 2516 12824 2870 12880
rect 2926 12824 2931 12880
rect 2516 12822 2931 12824
rect 2516 12820 2522 12822
rect 2865 12819 2931 12822
rect 6821 12882 6887 12885
rect 10593 12882 10659 12885
rect 6821 12880 10659 12882
rect 6821 12824 6826 12880
rect 6882 12824 10598 12880
rect 10654 12824 10659 12880
rect 6821 12822 10659 12824
rect 12712 12882 12772 12958
rect 13077 13016 16314 13018
rect 13077 12960 13082 13016
rect 13138 12960 16314 13016
rect 13077 12958 16314 12960
rect 13077 12955 13143 12958
rect 16614 12956 16620 13020
rect 16684 13018 16690 13020
rect 17585 13018 17651 13021
rect 16684 13016 17651 13018
rect 16684 12960 17590 13016
rect 17646 12960 17651 13016
rect 16684 12958 17651 12960
rect 16684 12956 16690 12958
rect 17585 12955 17651 12958
rect 18597 13018 18663 13021
rect 18597 13016 20362 13018
rect 18597 12960 18602 13016
rect 18658 12960 20362 13016
rect 18597 12958 20362 12960
rect 18597 12955 18663 12958
rect 14222 12882 14228 12884
rect 12712 12822 14228 12882
rect 6821 12819 6887 12822
rect 10593 12819 10659 12822
rect 14222 12820 14228 12822
rect 14292 12820 14298 12884
rect 14733 12882 14799 12885
rect 17534 12882 17540 12884
rect 14733 12880 17540 12882
rect 14733 12824 14738 12880
rect 14794 12824 17540 12880
rect 14733 12822 17540 12824
rect 14733 12819 14799 12822
rect 17534 12820 17540 12822
rect 17604 12820 17610 12884
rect 17718 12820 17724 12884
rect 17788 12882 17794 12884
rect 20161 12882 20227 12885
rect 17788 12880 20227 12882
rect 17788 12824 20166 12880
rect 20222 12824 20227 12880
rect 17788 12822 20227 12824
rect 20302 12882 20362 12958
rect 21030 12956 21036 13020
rect 21100 13018 21106 13020
rect 23381 13018 23447 13021
rect 21100 13016 23447 13018
rect 21100 12960 23386 13016
rect 23442 12960 23447 13016
rect 21100 12958 23447 12960
rect 21100 12956 21106 12958
rect 23381 12955 23447 12958
rect 25221 13018 25287 13021
rect 26200 13018 27000 13048
rect 25221 13016 27000 13018
rect 25221 12960 25226 13016
rect 25282 12960 27000 13016
rect 25221 12958 27000 12960
rect 25221 12955 25287 12958
rect 26200 12928 27000 12958
rect 21357 12882 21423 12885
rect 20302 12880 21423 12882
rect 20302 12824 21362 12880
rect 21418 12824 21423 12880
rect 20302 12822 21423 12824
rect 17788 12820 17794 12822
rect 20161 12819 20227 12822
rect 21357 12819 21423 12822
rect 21725 12882 21791 12885
rect 22001 12882 22067 12885
rect 21725 12880 22067 12882
rect 21725 12824 21730 12880
rect 21786 12824 22006 12880
rect 22062 12824 22067 12880
rect 21725 12822 22067 12824
rect 21725 12819 21791 12822
rect 22001 12819 22067 12822
rect 4705 12746 4771 12749
rect 6821 12746 6887 12749
rect 4705 12744 6887 12746
rect 4705 12688 4710 12744
rect 4766 12688 6826 12744
rect 6882 12688 6887 12744
rect 4705 12686 6887 12688
rect 4705 12683 4771 12686
rect 6821 12683 6887 12686
rect 7005 12746 7071 12749
rect 8569 12746 8635 12749
rect 12617 12746 12683 12749
rect 13077 12746 13143 12749
rect 7005 12744 8635 12746
rect 7005 12688 7010 12744
rect 7066 12688 8574 12744
rect 8630 12688 8635 12744
rect 7005 12686 8635 12688
rect 7005 12683 7071 12686
rect 8569 12683 8635 12686
rect 8710 12744 12683 12746
rect 8710 12688 12622 12744
rect 12678 12688 12683 12744
rect 8710 12686 12683 12688
rect 5809 12610 5875 12613
rect 8710 12610 8770 12686
rect 12617 12683 12683 12686
rect 12804 12744 13143 12746
rect 12804 12688 13082 12744
rect 13138 12688 13143 12744
rect 12804 12686 13143 12688
rect 11697 12610 11763 12613
rect 5809 12608 8770 12610
rect 5809 12552 5814 12608
rect 5870 12552 8770 12608
rect 5809 12550 8770 12552
rect 8894 12608 11763 12610
rect 8894 12552 11702 12608
rect 11758 12552 11763 12608
rect 8894 12550 11763 12552
rect 5809 12547 5875 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 5257 12474 5323 12477
rect 6126 12474 6132 12476
rect 5257 12472 6132 12474
rect 5257 12416 5262 12472
rect 5318 12416 6132 12472
rect 5257 12414 6132 12416
rect 5257 12411 5323 12414
rect 6126 12412 6132 12414
rect 6196 12412 6202 12476
rect 6913 12474 6979 12477
rect 8894 12474 8954 12550
rect 11697 12547 11763 12550
rect 12433 12610 12499 12613
rect 12804 12610 12864 12686
rect 13077 12683 13143 12686
rect 13261 12746 13327 12749
rect 14089 12746 14155 12749
rect 19006 12746 19012 12748
rect 13261 12744 13922 12746
rect 13261 12688 13266 12744
rect 13322 12688 13922 12744
rect 13261 12686 13922 12688
rect 13261 12683 13327 12686
rect 12433 12608 12864 12610
rect 12433 12552 12438 12608
rect 12494 12552 12864 12608
rect 12433 12550 12864 12552
rect 13862 12610 13922 12686
rect 14089 12744 19012 12746
rect 14089 12688 14094 12744
rect 14150 12688 19012 12744
rect 14089 12686 19012 12688
rect 14089 12683 14155 12686
rect 19006 12684 19012 12686
rect 19076 12684 19082 12748
rect 19149 12746 19215 12749
rect 22645 12746 22711 12749
rect 19149 12744 19258 12746
rect 19149 12688 19154 12744
rect 19210 12688 19258 12744
rect 19149 12683 19258 12688
rect 15193 12610 15259 12613
rect 13862 12608 15259 12610
rect 13862 12552 15198 12608
rect 15254 12552 15259 12608
rect 13862 12550 15259 12552
rect 12433 12547 12499 12550
rect 15193 12547 15259 12550
rect 15469 12610 15535 12613
rect 18873 12612 18939 12613
rect 15469 12608 18154 12610
rect 15469 12552 15474 12608
rect 15530 12552 18154 12608
rect 15469 12550 18154 12552
rect 15469 12547 15535 12550
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 6913 12472 8954 12474
rect 6913 12416 6918 12472
rect 6974 12416 8954 12472
rect 6913 12414 8954 12416
rect 6913 12411 6979 12414
rect 9990 12412 9996 12476
rect 10060 12474 10066 12476
rect 11513 12474 11579 12477
rect 12341 12476 12407 12477
rect 12341 12474 12388 12476
rect 10060 12472 11579 12474
rect 10060 12416 11518 12472
rect 11574 12416 11579 12472
rect 10060 12414 11579 12416
rect 12296 12472 12388 12474
rect 12296 12416 12346 12472
rect 12296 12414 12388 12416
rect 10060 12412 10066 12414
rect 11513 12411 11579 12414
rect 12341 12412 12388 12414
rect 12452 12412 12458 12476
rect 13997 12474 14063 12477
rect 17861 12474 17927 12477
rect 13997 12472 17927 12474
rect 13997 12416 14002 12472
rect 14058 12416 17866 12472
rect 17922 12416 17927 12472
rect 13997 12414 17927 12416
rect 18094 12474 18154 12550
rect 18822 12548 18828 12612
rect 18892 12610 18939 12612
rect 19198 12610 19258 12683
rect 19428 12744 22711 12746
rect 19428 12688 22650 12744
rect 22706 12688 22711 12744
rect 19428 12686 22711 12688
rect 19428 12613 19488 12686
rect 22645 12683 22711 12686
rect 18892 12608 19258 12610
rect 18934 12552 19258 12608
rect 18892 12550 19258 12552
rect 19425 12608 19491 12613
rect 19425 12552 19430 12608
rect 19486 12552 19491 12608
rect 18892 12548 18939 12550
rect 18873 12547 18939 12548
rect 19425 12547 19491 12552
rect 22185 12610 22251 12613
rect 22645 12610 22711 12613
rect 22185 12608 22711 12610
rect 22185 12552 22190 12608
rect 22246 12552 22650 12608
rect 22706 12552 22711 12608
rect 22185 12550 22711 12552
rect 22185 12547 22251 12550
rect 22645 12547 22711 12550
rect 24669 12610 24735 12613
rect 24894 12610 24900 12612
rect 24669 12608 24900 12610
rect 24669 12552 24674 12608
rect 24730 12552 24900 12608
rect 24669 12550 24900 12552
rect 24669 12547 24735 12550
rect 24894 12548 24900 12550
rect 24964 12548 24970 12612
rect 25129 12610 25195 12613
rect 26200 12610 27000 12640
rect 25129 12608 27000 12610
rect 25129 12552 25134 12608
rect 25190 12552 27000 12608
rect 25129 12550 27000 12552
rect 25129 12547 25195 12550
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 26200 12520 27000 12550
rect 22946 12479 23262 12480
rect 19701 12474 19767 12477
rect 18094 12472 19767 12474
rect 18094 12416 19706 12472
rect 19762 12416 19767 12472
rect 18094 12414 19767 12416
rect 12341 12411 12407 12412
rect 13997 12411 14063 12414
rect 17861 12411 17927 12414
rect 19701 12411 19767 12414
rect 3509 12338 3575 12341
rect 6310 12338 6316 12340
rect 3509 12336 6316 12338
rect 3509 12280 3514 12336
rect 3570 12280 6316 12336
rect 3509 12278 6316 12280
rect 3509 12275 3575 12278
rect 6310 12276 6316 12278
rect 6380 12276 6386 12340
rect 7557 12338 7623 12341
rect 7833 12338 7899 12341
rect 12525 12340 12591 12341
rect 12525 12338 12572 12340
rect 7557 12336 7899 12338
rect 7557 12280 7562 12336
rect 7618 12280 7838 12336
rect 7894 12280 7899 12336
rect 7557 12278 7899 12280
rect 12480 12336 12572 12338
rect 12480 12280 12530 12336
rect 12480 12278 12572 12280
rect 7557 12275 7623 12278
rect 7833 12275 7899 12278
rect 12525 12276 12572 12278
rect 12636 12276 12642 12340
rect 12801 12338 12867 12341
rect 15285 12338 15351 12341
rect 12801 12336 15351 12338
rect 12801 12280 12806 12336
rect 12862 12280 15290 12336
rect 15346 12280 15351 12336
rect 12801 12278 15351 12280
rect 12525 12275 12591 12276
rect 12801 12275 12867 12278
rect 15285 12275 15351 12278
rect 16757 12338 16823 12341
rect 17534 12338 17540 12340
rect 16757 12336 17540 12338
rect 16757 12280 16762 12336
rect 16818 12280 17540 12336
rect 16757 12278 17540 12280
rect 16757 12275 16823 12278
rect 17534 12276 17540 12278
rect 17604 12338 17610 12340
rect 18505 12338 18571 12341
rect 17604 12336 18571 12338
rect 17604 12280 18510 12336
rect 18566 12280 18571 12336
rect 17604 12278 18571 12280
rect 17604 12276 17610 12278
rect 18505 12275 18571 12278
rect 19006 12276 19012 12340
rect 19076 12338 19082 12340
rect 20345 12338 20411 12341
rect 19076 12336 20411 12338
rect 19076 12280 20350 12336
rect 20406 12280 20411 12336
rect 19076 12278 20411 12280
rect 19076 12276 19082 12278
rect 20345 12275 20411 12278
rect 21541 12338 21607 12341
rect 21817 12338 21883 12341
rect 21541 12336 21883 12338
rect 21541 12280 21546 12336
rect 21602 12280 21822 12336
rect 21878 12280 21883 12336
rect 21541 12278 21883 12280
rect 21541 12275 21607 12278
rect 21817 12275 21883 12278
rect 2589 12202 2655 12205
rect 24117 12202 24183 12205
rect 2589 12200 24183 12202
rect 2589 12144 2594 12200
rect 2650 12144 24122 12200
rect 24178 12144 24183 12200
rect 2589 12142 24183 12144
rect 2589 12139 2655 12142
rect 24117 12139 24183 12142
rect 25037 12202 25103 12205
rect 26200 12202 27000 12232
rect 25037 12200 27000 12202
rect 25037 12144 25042 12200
rect 25098 12144 27000 12200
rect 25037 12142 27000 12144
rect 25037 12139 25103 12142
rect 26200 12112 27000 12142
rect 10542 12004 10548 12068
rect 10612 12066 10618 12068
rect 10961 12066 11027 12069
rect 12750 12066 12756 12068
rect 10612 12064 11027 12066
rect 10612 12008 10966 12064
rect 11022 12008 11027 12064
rect 10612 12006 11027 12008
rect 10612 12004 10618 12006
rect 10961 12003 11027 12006
rect 12390 12006 12756 12066
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 9673 11930 9739 11933
rect 11237 11930 11303 11933
rect 11462 11930 11468 11932
rect 9673 11928 11468 11930
rect 9673 11872 9678 11928
rect 9734 11872 11242 11928
rect 11298 11872 11468 11928
rect 9673 11870 11468 11872
rect 9673 11867 9739 11870
rect 11237 11867 11303 11870
rect 11462 11868 11468 11870
rect 11532 11868 11538 11932
rect 5165 11794 5231 11797
rect 5758 11794 5764 11796
rect 5165 11792 5764 11794
rect 5165 11736 5170 11792
rect 5226 11736 5764 11792
rect 5165 11734 5764 11736
rect 5165 11731 5231 11734
rect 5758 11732 5764 11734
rect 5828 11732 5834 11796
rect 6177 11794 6243 11797
rect 12390 11794 12450 12006
rect 12750 12004 12756 12006
rect 12820 12004 12826 12068
rect 16062 12004 16068 12068
rect 16132 12066 16138 12068
rect 16757 12066 16823 12069
rect 16132 12064 16823 12066
rect 16132 12008 16762 12064
rect 16818 12008 16823 12064
rect 16132 12006 16823 12008
rect 16132 12004 16138 12006
rect 16757 12003 16823 12006
rect 19609 12066 19675 12069
rect 24669 12066 24735 12069
rect 19609 12064 24735 12066
rect 19609 12008 19614 12064
rect 19670 12008 24674 12064
rect 24730 12008 24735 12064
rect 19609 12006 24735 12008
rect 19609 12003 19675 12006
rect 24669 12003 24735 12006
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 23565 11930 23631 11933
rect 23790 11930 23796 11932
rect 23565 11928 23796 11930
rect 23565 11872 23570 11928
rect 23626 11872 23796 11928
rect 23565 11870 23796 11872
rect 23565 11867 23631 11870
rect 23790 11868 23796 11870
rect 23860 11868 23866 11932
rect 6177 11792 12450 11794
rect 6177 11736 6182 11792
rect 6238 11736 12450 11792
rect 6177 11734 12450 11736
rect 6177 11731 6243 11734
rect 17718 11732 17724 11796
rect 17788 11794 17794 11796
rect 17861 11794 17927 11797
rect 17788 11792 17927 11794
rect 17788 11736 17866 11792
rect 17922 11736 17927 11792
rect 17788 11734 17927 11736
rect 17788 11732 17794 11734
rect 17861 11731 17927 11734
rect 18045 11794 18111 11797
rect 19190 11794 19196 11796
rect 18045 11792 19196 11794
rect 18045 11736 18050 11792
rect 18106 11736 19196 11792
rect 18045 11734 19196 11736
rect 18045 11731 18111 11734
rect 19190 11732 19196 11734
rect 19260 11732 19266 11796
rect 23933 11794 23999 11797
rect 19566 11792 23999 11794
rect 19566 11736 23938 11792
rect 23994 11736 23999 11792
rect 19566 11734 23999 11736
rect 1853 11658 1919 11661
rect 10726 11658 10732 11660
rect 1853 11656 10732 11658
rect 1853 11600 1858 11656
rect 1914 11600 10732 11656
rect 1853 11598 10732 11600
rect 1853 11595 1919 11598
rect 10726 11596 10732 11598
rect 10796 11596 10802 11660
rect 16849 11658 16915 11661
rect 19374 11658 19380 11660
rect 12390 11656 19380 11658
rect 12390 11600 16854 11656
rect 16910 11600 19380 11656
rect 12390 11598 19380 11600
rect 3550 11460 3556 11524
rect 3620 11522 3626 11524
rect 3785 11522 3851 11525
rect 3620 11520 3851 11522
rect 3620 11464 3790 11520
rect 3846 11464 3851 11520
rect 3620 11462 3851 11464
rect 3620 11460 3626 11462
rect 3785 11459 3851 11462
rect 4613 11522 4679 11525
rect 10358 11522 10364 11524
rect 4613 11520 10364 11522
rect 4613 11464 4618 11520
rect 4674 11464 10364 11520
rect 4613 11462 10364 11464
rect 4613 11459 4679 11462
rect 10358 11460 10364 11462
rect 10428 11460 10434 11524
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 1853 11388 1919 11389
rect 1853 11386 1900 11388
rect 1808 11384 1900 11386
rect 1808 11328 1858 11384
rect 1808 11326 1900 11328
rect 1853 11324 1900 11326
rect 1964 11324 1970 11388
rect 8385 11386 8451 11389
rect 8518 11386 8524 11388
rect 8385 11384 8524 11386
rect 8385 11328 8390 11384
rect 8446 11328 8524 11384
rect 8385 11326 8524 11328
rect 1853 11323 1919 11324
rect 8385 11323 8451 11326
rect 8518 11324 8524 11326
rect 8588 11324 8594 11388
rect 2037 11250 2103 11253
rect 3417 11250 3483 11253
rect 6913 11252 6979 11253
rect 2037 11248 3483 11250
rect 2037 11192 2042 11248
rect 2098 11192 3422 11248
rect 3478 11192 3483 11248
rect 2037 11190 3483 11192
rect 2037 11187 2103 11190
rect 3417 11187 3483 11190
rect 6862 11188 6868 11252
rect 6932 11250 6979 11252
rect 6932 11248 7024 11250
rect 6974 11192 7024 11248
rect 6932 11190 7024 11192
rect 6932 11188 6979 11190
rect 6913 11187 6979 11188
rect 2405 11114 2471 11117
rect 12390 11114 12450 11598
rect 16849 11595 16915 11598
rect 19374 11596 19380 11598
rect 19444 11596 19450 11660
rect 13445 11522 13511 11525
rect 19566 11522 19626 11734
rect 23933 11731 23999 11734
rect 24761 11794 24827 11797
rect 26200 11794 27000 11824
rect 24761 11792 27000 11794
rect 24761 11736 24766 11792
rect 24822 11736 27000 11792
rect 24761 11734 27000 11736
rect 24761 11731 24827 11734
rect 26200 11704 27000 11734
rect 21214 11596 21220 11660
rect 21284 11658 21290 11660
rect 25078 11658 25084 11660
rect 21284 11598 25084 11658
rect 21284 11596 21290 11598
rect 25078 11596 25084 11598
rect 25148 11596 25154 11660
rect 21725 11524 21791 11525
rect 21725 11522 21772 11524
rect 13445 11520 19626 11522
rect 13445 11464 13450 11520
rect 13506 11464 19626 11520
rect 13445 11462 19626 11464
rect 21680 11520 21772 11522
rect 21680 11464 21730 11520
rect 21680 11462 21772 11464
rect 13445 11459 13511 11462
rect 21725 11460 21772 11462
rect 21836 11460 21842 11524
rect 21725 11459 21791 11460
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 14365 11386 14431 11389
rect 18505 11386 18571 11389
rect 19609 11386 19675 11389
rect 14365 11384 18571 11386
rect 14365 11328 14370 11384
rect 14426 11328 18510 11384
rect 18566 11328 18571 11384
rect 14365 11326 18571 11328
rect 14365 11323 14431 11326
rect 18505 11323 18571 11326
rect 18646 11384 19675 11386
rect 18646 11328 19614 11384
rect 19670 11328 19675 11384
rect 18646 11326 19675 11328
rect 13813 11250 13879 11253
rect 15878 11250 15884 11252
rect 13813 11248 15884 11250
rect 13813 11192 13818 11248
rect 13874 11192 15884 11248
rect 13813 11190 15884 11192
rect 13813 11187 13879 11190
rect 15878 11188 15884 11190
rect 15948 11188 15954 11252
rect 17033 11250 17099 11253
rect 18646 11250 18706 11326
rect 19609 11323 19675 11326
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 17033 11248 18706 11250
rect 17033 11192 17038 11248
rect 17094 11192 18706 11248
rect 17033 11190 18706 11192
rect 19333 11250 19399 11253
rect 25446 11250 25452 11252
rect 19333 11248 25452 11250
rect 19333 11192 19338 11248
rect 19394 11192 25452 11248
rect 19333 11190 25452 11192
rect 17033 11187 17099 11190
rect 19333 11187 19399 11190
rect 25446 11188 25452 11190
rect 25516 11188 25522 11252
rect 14774 11114 14780 11116
rect 2405 11112 12450 11114
rect 2405 11056 2410 11112
rect 2466 11056 12450 11112
rect 2405 11054 12450 11056
rect 12528 11054 14780 11114
rect 2405 11051 2471 11054
rect 4429 10978 4495 10981
rect 4654 10978 4660 10980
rect 4429 10976 4660 10978
rect 4429 10920 4434 10976
rect 4490 10920 4660 10976
rect 4429 10918 4660 10920
rect 4429 10915 4495 10918
rect 4654 10916 4660 10918
rect 4724 10916 4730 10980
rect 12341 10978 12407 10981
rect 12528 10978 12588 11054
rect 14774 11052 14780 11054
rect 14844 11052 14850 11116
rect 15193 11114 15259 11117
rect 16246 11114 16252 11116
rect 15193 11112 16252 11114
rect 15193 11056 15198 11112
rect 15254 11056 16252 11112
rect 15193 11054 16252 11056
rect 15193 11051 15259 11054
rect 16246 11052 16252 11054
rect 16316 11052 16322 11116
rect 16430 11052 16436 11116
rect 16500 11114 16506 11116
rect 17953 11114 18019 11117
rect 16500 11112 18019 11114
rect 16500 11056 17958 11112
rect 18014 11056 18019 11112
rect 16500 11054 18019 11056
rect 16500 11052 16506 11054
rect 17953 11051 18019 11054
rect 18321 11114 18387 11117
rect 18454 11114 18460 11116
rect 18321 11112 18460 11114
rect 18321 11056 18326 11112
rect 18382 11056 18460 11112
rect 18321 11054 18460 11056
rect 18321 11051 18387 11054
rect 18454 11052 18460 11054
rect 18524 11052 18530 11116
rect 19190 11052 19196 11116
rect 19260 11114 19266 11116
rect 20846 11114 20852 11116
rect 19260 11054 20852 11114
rect 19260 11052 19266 11054
rect 20846 11052 20852 11054
rect 20916 11052 20922 11116
rect 21173 11114 21239 11117
rect 24025 11114 24091 11117
rect 21173 11112 24091 11114
rect 21173 11056 21178 11112
rect 21234 11056 24030 11112
rect 24086 11056 24091 11112
rect 21173 11054 24091 11056
rect 21173 11051 21239 11054
rect 24025 11051 24091 11054
rect 20110 10978 20116 10980
rect 12341 10976 12588 10978
rect 12341 10920 12346 10976
rect 12402 10920 12588 10976
rect 12341 10918 12588 10920
rect 18462 10918 20116 10978
rect 12341 10915 12407 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 4337 10842 4403 10845
rect 5574 10842 5580 10844
rect 4337 10840 5580 10842
rect 4337 10784 4342 10840
rect 4398 10784 5580 10840
rect 4337 10782 5580 10784
rect 4337 10779 4403 10782
rect 5574 10780 5580 10782
rect 5644 10780 5650 10844
rect 7097 10842 7163 10845
rect 7230 10842 7236 10844
rect 7097 10840 7236 10842
rect 7097 10784 7102 10840
rect 7158 10784 7236 10840
rect 7097 10782 7236 10784
rect 7097 10779 7163 10782
rect 7230 10780 7236 10782
rect 7300 10780 7306 10844
rect 16614 10842 16620 10844
rect 9630 10782 16620 10842
rect 7782 10644 7788 10708
rect 7852 10706 7858 10708
rect 9213 10706 9279 10709
rect 7852 10704 9279 10706
rect 7852 10648 9218 10704
rect 9274 10648 9279 10704
rect 7852 10646 9279 10648
rect 7852 10644 7858 10646
rect 9213 10643 9279 10646
rect 4245 10570 4311 10573
rect 9630 10570 9690 10782
rect 16614 10780 16620 10782
rect 16684 10780 16690 10844
rect 17166 10780 17172 10844
rect 17236 10842 17242 10844
rect 17493 10842 17559 10845
rect 17236 10840 17559 10842
rect 17236 10784 17498 10840
rect 17554 10784 17559 10840
rect 17236 10782 17559 10784
rect 17236 10780 17242 10782
rect 17493 10779 17559 10782
rect 10593 10706 10659 10709
rect 13854 10706 13860 10708
rect 10593 10704 13860 10706
rect 10593 10648 10598 10704
rect 10654 10648 13860 10704
rect 10593 10646 13860 10648
rect 10593 10643 10659 10646
rect 13854 10644 13860 10646
rect 13924 10644 13930 10708
rect 18462 10706 18522 10918
rect 20110 10916 20116 10918
rect 20180 10916 20186 10980
rect 20529 10978 20595 10981
rect 22318 10978 22324 10980
rect 20529 10976 22324 10978
rect 20529 10920 20534 10976
rect 20590 10920 22324 10976
rect 20529 10918 22324 10920
rect 20529 10915 20595 10918
rect 22318 10916 22324 10918
rect 22388 10916 22394 10980
rect 25129 10978 25195 10981
rect 26200 10978 27000 11008
rect 25129 10976 27000 10978
rect 25129 10920 25134 10976
rect 25190 10920 27000 10976
rect 25129 10918 27000 10920
rect 25129 10915 25195 10918
rect 26200 10888 27000 10918
rect 19374 10780 19380 10844
rect 19444 10842 19450 10844
rect 21398 10842 21404 10844
rect 19444 10782 21404 10842
rect 19444 10780 19450 10782
rect 21398 10780 21404 10782
rect 21468 10780 21474 10844
rect 22502 10706 22508 10708
rect 14000 10646 18522 10706
rect 19566 10646 22508 10706
rect 4245 10568 9690 10570
rect 4245 10512 4250 10568
rect 4306 10512 9690 10568
rect 4245 10510 9690 10512
rect 4245 10507 4311 10510
rect 3785 10434 3851 10437
rect 10910 10434 10916 10436
rect 3785 10432 10916 10434
rect 3785 10376 3790 10432
rect 3846 10376 10916 10432
rect 3785 10374 10916 10376
rect 3785 10371 3851 10374
rect 10910 10372 10916 10374
rect 10980 10372 10986 10436
rect 13445 10434 13511 10437
rect 14000 10434 14060 10646
rect 14549 10570 14615 10573
rect 19425 10570 19491 10573
rect 14549 10568 19491 10570
rect 14549 10512 14554 10568
rect 14610 10512 19430 10568
rect 19486 10512 19491 10568
rect 14549 10510 19491 10512
rect 14549 10507 14615 10510
rect 19425 10507 19491 10510
rect 13445 10432 14060 10434
rect 13445 10376 13450 10432
rect 13506 10376 14060 10432
rect 13445 10374 14060 10376
rect 15193 10434 15259 10437
rect 18965 10434 19031 10437
rect 15193 10432 19031 10434
rect 15193 10376 15198 10432
rect 15254 10376 18970 10432
rect 19026 10376 19031 10432
rect 15193 10374 19031 10376
rect 13445 10371 13511 10374
rect 15193 10371 15259 10374
rect 18965 10371 19031 10374
rect 19425 10434 19491 10437
rect 19566 10434 19626 10646
rect 22502 10644 22508 10646
rect 22572 10644 22578 10708
rect 25129 10570 25195 10573
rect 26200 10570 27000 10600
rect 25129 10568 27000 10570
rect 25129 10512 25134 10568
rect 25190 10512 27000 10568
rect 25129 10510 27000 10512
rect 25129 10507 25195 10510
rect 26200 10480 27000 10510
rect 19425 10432 19626 10434
rect 19425 10376 19430 10432
rect 19486 10376 19626 10432
rect 19425 10374 19626 10376
rect 24209 10434 24275 10437
rect 25630 10434 25636 10436
rect 24209 10432 25636 10434
rect 24209 10376 24214 10432
rect 24270 10376 25636 10432
rect 24209 10374 25636 10376
rect 19425 10371 19491 10374
rect 24209 10371 24275 10374
rect 25630 10372 25636 10374
rect 25700 10372 25706 10436
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 6085 10298 6151 10301
rect 12525 10298 12591 10301
rect 6085 10296 12591 10298
rect 6085 10240 6090 10296
rect 6146 10240 12530 10296
rect 12586 10240 12591 10296
rect 6085 10238 12591 10240
rect 6085 10235 6151 10238
rect 12525 10235 12591 10238
rect 15285 10298 15351 10301
rect 19333 10298 19399 10301
rect 23974 10298 23980 10300
rect 15285 10296 19399 10298
rect 15285 10240 15290 10296
rect 15346 10240 19338 10296
rect 19394 10240 19399 10296
rect 15285 10238 19399 10240
rect 15285 10235 15351 10238
rect 19333 10235 19399 10238
rect 23384 10238 23980 10298
rect 7414 10100 7420 10164
rect 7484 10162 7490 10164
rect 10593 10162 10659 10165
rect 13997 10162 14063 10165
rect 7484 10160 14063 10162
rect 7484 10104 10598 10160
rect 10654 10104 14002 10160
rect 14058 10104 14063 10160
rect 7484 10102 14063 10104
rect 7484 10100 7490 10102
rect 10593 10099 10659 10102
rect 13997 10099 14063 10102
rect 17534 10100 17540 10164
rect 17604 10162 17610 10164
rect 18822 10162 18828 10164
rect 17604 10102 18828 10162
rect 17604 10100 17610 10102
rect 18822 10100 18828 10102
rect 18892 10100 18898 10164
rect 18965 10162 19031 10165
rect 23384 10162 23444 10238
rect 23974 10236 23980 10238
rect 24044 10236 24050 10300
rect 24342 10236 24348 10300
rect 24412 10298 24418 10300
rect 25037 10298 25103 10301
rect 24412 10296 25103 10298
rect 24412 10240 25042 10296
rect 25098 10240 25103 10296
rect 24412 10238 25103 10240
rect 24412 10236 24418 10238
rect 25037 10235 25103 10238
rect 24209 10162 24275 10165
rect 18965 10160 23444 10162
rect 18965 10104 18970 10160
rect 19026 10104 23444 10160
rect 18965 10102 23444 10104
rect 23982 10160 24275 10162
rect 23982 10104 24214 10160
rect 24270 10104 24275 10160
rect 23982 10102 24275 10104
rect 18965 10099 19031 10102
rect 2773 10026 2839 10029
rect 23982 10026 24042 10102
rect 24209 10099 24275 10102
rect 24853 10162 24919 10165
rect 26200 10162 27000 10192
rect 24853 10160 27000 10162
rect 24853 10104 24858 10160
rect 24914 10104 27000 10160
rect 24853 10102 27000 10104
rect 24853 10099 24919 10102
rect 26200 10072 27000 10102
rect 2773 10024 24042 10026
rect 2773 9968 2778 10024
rect 2834 9968 24042 10024
rect 2773 9966 24042 9968
rect 2773 9963 2839 9966
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 13670 9692 13676 9756
rect 13740 9754 13746 9756
rect 15469 9754 15535 9757
rect 26200 9754 27000 9784
rect 13740 9752 15535 9754
rect 13740 9696 15474 9752
rect 15530 9696 15535 9752
rect 13740 9694 15535 9696
rect 13740 9692 13746 9694
rect 15469 9691 15535 9694
rect 24672 9694 27000 9754
rect 24672 9621 24732 9694
rect 26200 9664 27000 9694
rect 5165 9620 5231 9621
rect 5165 9618 5212 9620
rect 5120 9616 5212 9618
rect 5120 9560 5170 9616
rect 5120 9558 5212 9560
rect 5165 9556 5212 9558
rect 5276 9556 5282 9620
rect 7598 9556 7604 9620
rect 7668 9618 7674 9620
rect 7741 9618 7807 9621
rect 7668 9616 7807 9618
rect 7668 9560 7746 9616
rect 7802 9560 7807 9616
rect 7668 9558 7807 9560
rect 7668 9556 7674 9558
rect 5165 9555 5231 9556
rect 7741 9555 7807 9558
rect 10593 9618 10659 9621
rect 22645 9618 22711 9621
rect 10593 9616 22711 9618
rect 10593 9560 10598 9616
rect 10654 9560 22650 9616
rect 22706 9560 22711 9616
rect 10593 9558 22711 9560
rect 10593 9555 10659 9558
rect 22645 9555 22711 9558
rect 24669 9616 24735 9621
rect 24669 9560 24674 9616
rect 24730 9560 24735 9616
rect 24669 9555 24735 9560
rect 2313 9482 2379 9485
rect 8569 9482 8635 9485
rect 16430 9482 16436 9484
rect 2313 9480 3802 9482
rect 2313 9424 2318 9480
rect 2374 9424 3802 9480
rect 2313 9422 3802 9424
rect 2313 9419 2379 9422
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 606 9148 612 9212
rect 676 9210 682 9212
rect 1577 9210 1643 9213
rect 676 9208 1643 9210
rect 676 9152 1582 9208
rect 1638 9152 1643 9208
rect 676 9150 1643 9152
rect 3742 9210 3802 9422
rect 8569 9480 16436 9482
rect 8569 9424 8574 9480
rect 8630 9424 16436 9480
rect 8569 9422 16436 9424
rect 8569 9419 8635 9422
rect 16430 9420 16436 9422
rect 16500 9420 16506 9484
rect 3918 9284 3924 9348
rect 3988 9346 3994 9348
rect 12709 9346 12775 9349
rect 3988 9344 12775 9346
rect 3988 9288 12714 9344
rect 12770 9288 12775 9344
rect 3988 9286 12775 9288
rect 3988 9284 3994 9286
rect 12709 9283 12775 9286
rect 24853 9346 24919 9349
rect 26200 9346 27000 9376
rect 24853 9344 27000 9346
rect 24853 9288 24858 9344
rect 24914 9288 27000 9344
rect 24853 9286 27000 9288
rect 24853 9283 24919 9286
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 26200 9256 27000 9286
rect 22946 9215 23262 9216
rect 4705 9210 4771 9213
rect 9806 9210 9812 9212
rect 3742 9150 4354 9210
rect 676 9148 682 9150
rect 1577 9147 1643 9150
rect 974 9012 980 9076
rect 1044 9074 1050 9076
rect 4153 9074 4219 9077
rect 1044 9072 4219 9074
rect 1044 9016 4158 9072
rect 4214 9016 4219 9072
rect 1044 9014 4219 9016
rect 4294 9074 4354 9150
rect 4705 9208 9812 9210
rect 4705 9152 4710 9208
rect 4766 9152 9812 9208
rect 4705 9150 9812 9152
rect 4705 9147 4771 9150
rect 9806 9148 9812 9150
rect 9876 9148 9882 9212
rect 12198 9074 12204 9076
rect 4294 9014 12204 9074
rect 1044 9012 1050 9014
rect 4153 9011 4219 9014
rect 12198 9012 12204 9014
rect 12268 9012 12274 9076
rect 12566 9012 12572 9076
rect 12636 9074 12642 9076
rect 22093 9074 22159 9077
rect 12636 9072 22159 9074
rect 12636 9016 22098 9072
rect 22154 9016 22159 9072
rect 12636 9014 22159 9016
rect 12636 9012 12642 9014
rect 22093 9011 22159 9014
rect 3734 8876 3740 8940
rect 3804 8938 3810 8940
rect 8477 8938 8543 8941
rect 3804 8936 8543 8938
rect 3804 8880 8482 8936
rect 8538 8880 8543 8936
rect 3804 8878 8543 8880
rect 3804 8876 3810 8878
rect 8477 8875 8543 8878
rect 14457 8938 14523 8941
rect 19374 8938 19380 8940
rect 14457 8936 19380 8938
rect 14457 8880 14462 8936
rect 14518 8880 19380 8936
rect 14457 8878 19380 8880
rect 14457 8875 14523 8878
rect 19374 8876 19380 8878
rect 19444 8876 19450 8940
rect 24945 8938 25011 8941
rect 26200 8938 27000 8968
rect 24945 8936 27000 8938
rect 24945 8880 24950 8936
rect 25006 8880 27000 8936
rect 24945 8878 27000 8880
rect 24945 8875 25011 8878
rect 26200 8848 27000 8878
rect 2262 8740 2268 8804
rect 2332 8802 2338 8804
rect 3233 8802 3299 8805
rect 2332 8800 3299 8802
rect 2332 8744 3238 8800
rect 3294 8744 3299 8800
rect 2332 8742 3299 8744
rect 2332 8740 2338 8742
rect 3233 8739 3299 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 2589 8668 2655 8669
rect 2589 8666 2636 8668
rect 2544 8664 2636 8666
rect 2544 8608 2594 8664
rect 2544 8606 2636 8608
rect 2589 8604 2636 8606
rect 2700 8604 2706 8668
rect 16113 8666 16179 8669
rect 17166 8666 17172 8668
rect 16113 8664 17172 8666
rect 16113 8608 16118 8664
rect 16174 8608 17172 8664
rect 16113 8606 17172 8608
rect 2589 8603 2655 8604
rect 16113 8603 16179 8606
rect 17166 8604 17172 8606
rect 17236 8604 17242 8668
rect 790 8468 796 8532
rect 860 8530 866 8532
rect 4153 8530 4219 8533
rect 860 8528 4219 8530
rect 860 8472 4158 8528
rect 4214 8472 4219 8528
rect 860 8470 4219 8472
rect 860 8468 866 8470
rect 4153 8467 4219 8470
rect 6678 8468 6684 8532
rect 6748 8530 6754 8532
rect 8753 8530 8819 8533
rect 6748 8528 8819 8530
rect 6748 8472 8758 8528
rect 8814 8472 8819 8528
rect 6748 8470 8819 8472
rect 6748 8468 6754 8470
rect 8753 8467 8819 8470
rect 10869 8530 10935 8533
rect 23933 8530 23999 8533
rect 10869 8528 23999 8530
rect 10869 8472 10874 8528
rect 10930 8472 23938 8528
rect 23994 8472 23999 8528
rect 10869 8470 23999 8472
rect 10869 8467 10935 8470
rect 23933 8467 23999 8470
rect 24761 8530 24827 8533
rect 26200 8530 27000 8560
rect 24761 8528 27000 8530
rect 24761 8472 24766 8528
rect 24822 8472 27000 8528
rect 24761 8470 27000 8472
rect 24761 8467 24827 8470
rect 26200 8440 27000 8470
rect 16297 8394 16363 8397
rect 22686 8394 22692 8396
rect 16297 8392 22692 8394
rect 16297 8336 16302 8392
rect 16358 8336 22692 8392
rect 16297 8334 22692 8336
rect 16297 8331 16363 8334
rect 22686 8332 22692 8334
rect 22756 8332 22762 8396
rect 13997 8258 14063 8261
rect 19006 8258 19012 8260
rect 13997 8256 19012 8258
rect 13997 8200 14002 8256
rect 14058 8200 19012 8256
rect 13997 8198 19012 8200
rect 13997 8195 14063 8198
rect 19006 8196 19012 8198
rect 19076 8196 19082 8260
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 9254 8060 9260 8124
rect 9324 8122 9330 8124
rect 12157 8122 12223 8125
rect 9324 8120 12223 8122
rect 9324 8064 12162 8120
rect 12218 8064 12223 8120
rect 9324 8062 12223 8064
rect 9324 8060 9330 8062
rect 12157 8059 12223 8062
rect 23381 8122 23447 8125
rect 26200 8122 27000 8152
rect 23381 8120 27000 8122
rect 23381 8064 23386 8120
rect 23442 8064 27000 8120
rect 23381 8062 27000 8064
rect 23381 8059 23447 8062
rect 26200 8032 27000 8062
rect 2589 7986 2655 7989
rect 4102 7986 4108 7988
rect 2589 7984 4108 7986
rect 2589 7928 2594 7984
rect 2650 7928 4108 7984
rect 2589 7926 4108 7928
rect 2589 7923 2655 7926
rect 4102 7924 4108 7926
rect 4172 7924 4178 7988
rect 5165 7986 5231 7989
rect 15101 7986 15167 7989
rect 5165 7984 15167 7986
rect 5165 7928 5170 7984
rect 5226 7928 15106 7984
rect 15162 7928 15167 7984
rect 5165 7926 15167 7928
rect 5165 7923 5231 7926
rect 15101 7923 15167 7926
rect 15285 7986 15351 7989
rect 24301 7986 24367 7989
rect 15285 7984 24367 7986
rect 15285 7928 15290 7984
rect 15346 7928 24306 7984
rect 24362 7928 24367 7984
rect 15285 7926 24367 7928
rect 15285 7923 15351 7926
rect 24301 7923 24367 7926
rect 4981 7850 5047 7853
rect 19241 7850 19307 7853
rect 4981 7848 19307 7850
rect 4981 7792 4986 7848
rect 5042 7792 19246 7848
rect 19302 7792 19307 7848
rect 4981 7790 19307 7792
rect 4981 7787 5047 7790
rect 19241 7787 19307 7790
rect 22829 7850 22895 7853
rect 25262 7850 25268 7852
rect 22829 7848 25268 7850
rect 22829 7792 22834 7848
rect 22890 7792 25268 7848
rect 22829 7790 25268 7792
rect 22829 7787 22895 7790
rect 25262 7788 25268 7790
rect 25332 7788 25338 7852
rect 24945 7714 25011 7717
rect 26200 7714 27000 7744
rect 24945 7712 27000 7714
rect 24945 7656 24950 7712
rect 25006 7656 27000 7712
rect 24945 7654 27000 7656
rect 24945 7651 25011 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 10409 7442 10475 7445
rect 23933 7442 23999 7445
rect 25998 7442 26004 7444
rect 10409 7440 23999 7442
rect 10409 7384 10414 7440
rect 10470 7384 23938 7440
rect 23994 7384 23999 7440
rect 10409 7382 23999 7384
rect 10409 7379 10475 7382
rect 23933 7379 23999 7382
rect 24166 7382 26004 7442
rect 3693 7306 3759 7309
rect 13813 7306 13879 7309
rect 16573 7306 16639 7309
rect 24166 7306 24226 7382
rect 25998 7380 26004 7382
rect 26068 7380 26074 7444
rect 3693 7304 13554 7306
rect 3693 7248 3698 7304
rect 3754 7248 13554 7304
rect 3693 7246 13554 7248
rect 3693 7243 3759 7246
rect 13494 7170 13554 7246
rect 13813 7304 24226 7306
rect 13813 7248 13818 7304
rect 13874 7248 16578 7304
rect 16634 7248 24226 7304
rect 13813 7246 24226 7248
rect 24669 7306 24735 7309
rect 26200 7306 27000 7336
rect 24669 7304 27000 7306
rect 24669 7248 24674 7304
rect 24730 7248 27000 7304
rect 24669 7246 27000 7248
rect 13813 7243 13879 7246
rect 16573 7243 16639 7246
rect 24669 7243 24735 7246
rect 26200 7216 27000 7246
rect 18413 7170 18479 7173
rect 13494 7168 18479 7170
rect 13494 7112 18418 7168
rect 18474 7112 18479 7168
rect 13494 7110 18479 7112
rect 18413 7107 18479 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 8845 6898 8911 6901
rect 15694 6898 15700 6900
rect 8845 6896 15700 6898
rect 8845 6840 8850 6896
rect 8906 6840 15700 6896
rect 8845 6838 15700 6840
rect 8845 6835 8911 6838
rect 15694 6836 15700 6838
rect 15764 6836 15770 6900
rect 23289 6898 23355 6901
rect 26200 6898 27000 6928
rect 23289 6896 27000 6898
rect 23289 6840 23294 6896
rect 23350 6840 27000 6896
rect 23289 6838 27000 6840
rect 23289 6835 23355 6838
rect 26200 6808 27000 6838
rect 4061 6762 4127 6765
rect 14406 6762 14412 6764
rect 4061 6760 14412 6762
rect 4061 6704 4066 6760
rect 4122 6704 14412 6760
rect 4061 6702 14412 6704
rect 4061 6699 4127 6702
rect 14406 6700 14412 6702
rect 14476 6700 14482 6764
rect 15377 6762 15443 6765
rect 15510 6762 15516 6764
rect 15377 6760 15516 6762
rect 15377 6704 15382 6760
rect 15438 6704 15516 6760
rect 15377 6702 15516 6704
rect 15377 6699 15443 6702
rect 15510 6700 15516 6702
rect 15580 6700 15586 6764
rect 25814 6762 25820 6764
rect 15702 6702 25820 6762
rect 12893 6626 12959 6629
rect 15702 6626 15762 6702
rect 25814 6700 25820 6702
rect 25884 6700 25890 6764
rect 12893 6624 15762 6626
rect 12893 6568 12898 6624
rect 12954 6568 15762 6624
rect 12893 6566 15762 6568
rect 12893 6563 12959 6566
rect 19742 6564 19748 6628
rect 19812 6626 19818 6628
rect 23933 6626 23999 6629
rect 19812 6624 23999 6626
rect 19812 6568 23938 6624
rect 23994 6568 23999 6624
rect 19812 6566 23999 6568
rect 19812 6564 19818 6566
rect 23933 6563 23999 6566
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 12341 6490 12407 6493
rect 17769 6490 17835 6493
rect 12341 6488 17835 6490
rect 12341 6432 12346 6488
rect 12402 6432 17774 6488
rect 17830 6432 17835 6488
rect 12341 6430 17835 6432
rect 12341 6427 12407 6430
rect 17769 6427 17835 6430
rect 25681 6490 25747 6493
rect 26200 6490 27000 6520
rect 25681 6488 27000 6490
rect 25681 6432 25686 6488
rect 25742 6432 27000 6488
rect 25681 6430 27000 6432
rect 25681 6427 25747 6430
rect 26200 6400 27000 6430
rect 1761 6354 1827 6357
rect 20805 6354 20871 6357
rect 1761 6352 20871 6354
rect 1761 6296 1766 6352
rect 1822 6296 20810 6352
rect 20866 6296 20871 6352
rect 1761 6294 20871 6296
rect 1761 6291 1827 6294
rect 20805 6291 20871 6294
rect 7465 6218 7531 6221
rect 19977 6218 20043 6221
rect 7465 6216 20043 6218
rect 7465 6160 7470 6216
rect 7526 6160 19982 6216
rect 20038 6160 20043 6216
rect 7465 6158 20043 6160
rect 7465 6155 7531 6158
rect 19977 6155 20043 6158
rect 13537 6082 13603 6085
rect 18505 6082 18571 6085
rect 13537 6080 18571 6082
rect 13537 6024 13542 6080
rect 13598 6024 18510 6080
rect 18566 6024 18571 6080
rect 13537 6022 18571 6024
rect 13537 6019 13603 6022
rect 18505 6019 18571 6022
rect 24761 6082 24827 6085
rect 26200 6082 27000 6112
rect 24761 6080 27000 6082
rect 24761 6024 24766 6080
rect 24822 6024 27000 6080
rect 24761 6022 27000 6024
rect 24761 6019 24827 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 26200 5992 27000 6022
rect 22946 5951 23262 5952
rect 16941 5948 17007 5949
rect 16941 5946 16988 5948
rect 16896 5944 16988 5946
rect 16896 5888 16946 5944
rect 16896 5886 16988 5888
rect 16941 5884 16988 5886
rect 17052 5884 17058 5948
rect 16941 5883 17007 5884
rect 6494 5748 6500 5812
rect 6564 5810 6570 5812
rect 16021 5810 16087 5813
rect 6564 5808 16087 5810
rect 6564 5752 16026 5808
rect 16082 5752 16087 5808
rect 6564 5750 16087 5752
rect 6564 5748 6570 5750
rect 16021 5747 16087 5750
rect 16297 5810 16363 5813
rect 19057 5810 19123 5813
rect 16297 5808 19123 5810
rect 16297 5752 16302 5808
rect 16358 5752 19062 5808
rect 19118 5752 19123 5808
rect 16297 5750 19123 5752
rect 16297 5747 16363 5750
rect 19057 5747 19123 5750
rect 6913 5674 6979 5677
rect 18873 5674 18939 5677
rect 6913 5672 18939 5674
rect 6913 5616 6918 5672
rect 6974 5616 18878 5672
rect 18934 5616 18939 5672
rect 6913 5614 18939 5616
rect 6913 5611 6979 5614
rect 18873 5611 18939 5614
rect 19057 5674 19123 5677
rect 23422 5674 23428 5676
rect 19057 5672 23428 5674
rect 19057 5616 19062 5672
rect 19118 5616 23428 5672
rect 19057 5614 23428 5616
rect 19057 5611 19123 5614
rect 23422 5612 23428 5614
rect 23492 5612 23498 5676
rect 24945 5674 25011 5677
rect 26200 5674 27000 5704
rect 24945 5672 27000 5674
rect 24945 5616 24950 5672
rect 25006 5616 27000 5672
rect 24945 5614 27000 5616
rect 24945 5611 25011 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 13537 5402 13603 5405
rect 16665 5402 16731 5405
rect 13537 5400 16731 5402
rect 13537 5344 13542 5400
rect 13598 5344 16670 5400
rect 16726 5344 16731 5400
rect 13537 5342 16731 5344
rect 13537 5339 13603 5342
rect 16665 5339 16731 5342
rect 17493 5266 17559 5269
rect 20294 5266 20300 5268
rect 17493 5264 20300 5266
rect 17493 5208 17498 5264
rect 17554 5208 20300 5264
rect 17493 5206 20300 5208
rect 17493 5203 17559 5206
rect 20294 5204 20300 5206
rect 20364 5204 20370 5268
rect 24577 5266 24643 5269
rect 26200 5266 27000 5296
rect 24577 5264 27000 5266
rect 24577 5208 24582 5264
rect 24638 5208 27000 5264
rect 24577 5206 27000 5208
rect 24577 5203 24643 5206
rect 26200 5176 27000 5206
rect 16481 5130 16547 5133
rect 24526 5130 24532 5132
rect 16481 5128 24532 5130
rect 16481 5072 16486 5128
rect 16542 5072 24532 5128
rect 16481 5070 24532 5072
rect 16481 5067 16547 5070
rect 24526 5068 24532 5070
rect 24596 5068 24602 5132
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 14590 4796 14596 4860
rect 14660 4858 14666 4860
rect 17125 4858 17191 4861
rect 14660 4856 17191 4858
rect 14660 4800 17130 4856
rect 17186 4800 17191 4856
rect 14660 4798 17191 4800
rect 14660 4796 14666 4798
rect 17125 4795 17191 4798
rect 24853 4858 24919 4861
rect 26200 4858 27000 4888
rect 24853 4856 27000 4858
rect 24853 4800 24858 4856
rect 24914 4800 27000 4856
rect 24853 4798 27000 4800
rect 24853 4795 24919 4798
rect 26200 4768 27000 4798
rect 8702 4524 8708 4588
rect 8772 4586 8778 4588
rect 17953 4586 18019 4589
rect 8772 4584 18019 4586
rect 8772 4528 17958 4584
rect 18014 4528 18019 4584
rect 8772 4526 18019 4528
rect 8772 4524 8778 4526
rect 17953 4523 18019 4526
rect 24945 4450 25011 4453
rect 26200 4450 27000 4480
rect 24945 4448 27000 4450
rect 24945 4392 24950 4448
rect 25006 4392 27000 4448
rect 24945 4390 27000 4392
rect 24945 4387 25011 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 26200 4360 27000 4390
rect 17946 4319 18262 4320
rect 17493 4316 17559 4317
rect 17493 4314 17540 4316
rect 17448 4312 17540 4314
rect 17448 4256 17498 4312
rect 17448 4254 17540 4256
rect 17493 4252 17540 4254
rect 17604 4252 17610 4316
rect 17493 4251 17559 4252
rect 11145 4178 11211 4181
rect 25630 4178 25636 4180
rect 11145 4176 25636 4178
rect 11145 4120 11150 4176
rect 11206 4120 25636 4176
rect 11145 4118 25636 4120
rect 11145 4115 11211 4118
rect 25630 4116 25636 4118
rect 25700 4116 25706 4180
rect 17033 4042 17099 4045
rect 18638 4042 18644 4044
rect 17033 4040 18644 4042
rect 17033 3984 17038 4040
rect 17094 3984 18644 4040
rect 17033 3982 18644 3984
rect 17033 3979 17099 3982
rect 18638 3980 18644 3982
rect 18708 3980 18714 4044
rect 18873 4042 18939 4045
rect 20662 4042 20668 4044
rect 18873 4040 20668 4042
rect 18873 3984 18878 4040
rect 18934 3984 20668 4040
rect 18873 3982 20668 3984
rect 18873 3979 18939 3982
rect 20662 3980 20668 3982
rect 20732 3980 20738 4044
rect 23381 4042 23447 4045
rect 26200 4042 27000 4072
rect 23381 4040 27000 4042
rect 23381 3984 23386 4040
rect 23442 3984 27000 4040
rect 23381 3982 27000 3984
rect 23381 3979 23447 3982
rect 26200 3952 27000 3982
rect 18597 3906 18663 3909
rect 19190 3906 19196 3908
rect 18597 3904 19196 3906
rect 18597 3848 18602 3904
rect 18658 3848 19196 3904
rect 18597 3846 19196 3848
rect 18597 3843 18663 3846
rect 19190 3844 19196 3846
rect 19260 3844 19266 3908
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 18229 3770 18295 3773
rect 21950 3770 21956 3772
rect 18229 3768 21956 3770
rect 18229 3712 18234 3768
rect 18290 3712 21956 3768
rect 18229 3710 21956 3712
rect 18229 3707 18295 3710
rect 21950 3708 21956 3710
rect 22020 3708 22026 3772
rect 13353 3634 13419 3637
rect 21030 3634 21036 3636
rect 13353 3632 21036 3634
rect 13353 3576 13358 3632
rect 13414 3576 21036 3632
rect 13353 3574 21036 3576
rect 13353 3571 13419 3574
rect 21030 3572 21036 3574
rect 21100 3572 21106 3636
rect 24945 3634 25011 3637
rect 26200 3634 27000 3664
rect 24945 3632 27000 3634
rect 24945 3576 24950 3632
rect 25006 3576 27000 3632
rect 24945 3574 27000 3576
rect 24945 3571 25011 3574
rect 26200 3544 27000 3574
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 25681 3226 25747 3229
rect 26200 3226 27000 3256
rect 25681 3224 27000 3226
rect 25681 3168 25686 3224
rect 25742 3168 27000 3224
rect 25681 3166 27000 3168
rect 25681 3163 25747 3166
rect 26200 3136 27000 3166
rect 8293 3090 8359 3093
rect 19057 3090 19123 3093
rect 8293 3088 19123 3090
rect 8293 3032 8298 3088
rect 8354 3032 19062 3088
rect 19118 3032 19123 3088
rect 8293 3030 19123 3032
rect 8293 3027 8359 3030
rect 19057 3027 19123 3030
rect 11830 2892 11836 2956
rect 11900 2954 11906 2956
rect 19425 2954 19491 2957
rect 11900 2952 19491 2954
rect 11900 2896 19430 2952
rect 19486 2896 19491 2952
rect 11900 2894 19491 2896
rect 11900 2892 11906 2894
rect 19425 2891 19491 2894
rect 24853 2818 24919 2821
rect 26200 2818 27000 2848
rect 24853 2816 27000 2818
rect 24853 2760 24858 2816
rect 24914 2760 27000 2816
rect 24853 2758 27000 2760
rect 24853 2755 24919 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 26200 2728 27000 2758
rect 22946 2687 23262 2688
rect 19609 2546 19675 2549
rect 24710 2546 24716 2548
rect 19609 2544 24716 2546
rect 19609 2488 19614 2544
rect 19670 2488 24716 2544
rect 19609 2486 24716 2488
rect 19609 2483 19675 2486
rect 24710 2484 24716 2486
rect 24780 2484 24786 2548
rect 10133 2410 10199 2413
rect 21214 2410 21220 2412
rect 10133 2408 21220 2410
rect 10133 2352 10138 2408
rect 10194 2352 21220 2408
rect 10133 2350 21220 2352
rect 10133 2347 10199 2350
rect 21214 2348 21220 2350
rect 21284 2348 21290 2412
rect 24945 2410 25011 2413
rect 26200 2410 27000 2440
rect 24945 2408 27000 2410
rect 24945 2352 24950 2408
rect 25006 2352 27000 2408
rect 24945 2350 27000 2352
rect 24945 2347 25011 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 22185 2002 22251 2005
rect 26200 2002 27000 2032
rect 22185 2000 27000 2002
rect 22185 1944 22190 2000
rect 22246 1944 27000 2000
rect 22185 1942 27000 1944
rect 22185 1939 22251 1942
rect 26200 1912 27000 1942
rect 22277 1594 22343 1597
rect 26200 1594 27000 1624
rect 22277 1592 27000 1594
rect 22277 1536 22282 1592
rect 22338 1536 27000 1592
rect 22277 1534 27000 1536
rect 22277 1531 22343 1534
rect 26200 1504 27000 1534
rect 23381 1186 23447 1189
rect 26200 1186 27000 1216
rect 23381 1184 27000 1186
rect 23381 1128 23386 1184
rect 23442 1128 27000 1184
rect 23381 1126 27000 1128
rect 23381 1123 23447 1126
rect 26200 1096 27000 1126
rect 25037 778 25103 781
rect 26200 778 27000 808
rect 25037 776 27000 778
rect 25037 720 25042 776
rect 25098 720 27000 776
rect 25037 718 27000 720
rect 25037 715 25103 718
rect 26200 688 27000 718
rect 24853 370 24919 373
rect 26200 370 27000 400
rect 24853 368 27000 370
rect 24853 312 24858 368
rect 24914 312 27000 368
rect 24853 310 27000 312
rect 24853 307 24919 310
rect 26200 280 27000 310
<< via3 >>
rect 9260 26692 9324 26756
rect 18460 26556 18524 26620
rect 18828 26420 18892 26484
rect 6132 26284 6196 26348
rect 796 26148 860 26212
rect 5212 25876 5276 25940
rect 796 25604 860 25668
rect 980 25468 1044 25532
rect 15148 25468 15212 25532
rect 4660 25332 4724 25396
rect 8340 25332 8404 25396
rect 11100 25332 11164 25396
rect 9444 25196 9508 25260
rect 9812 25060 9876 25124
rect 20668 25060 20732 25124
rect 9628 24924 9692 24988
rect 10548 24788 10612 24852
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7236 24380 7300 24444
rect 19012 24304 19076 24308
rect 19012 24248 19062 24304
rect 19062 24248 19076 24304
rect 19012 24244 19076 24248
rect 3556 24108 3620 24172
rect 2636 24032 2700 24036
rect 2636 23976 2650 24032
rect 2650 23976 2700 24032
rect 2636 23972 2700 23976
rect 11652 24108 11716 24172
rect 16620 24108 16684 24172
rect 12204 23972 12268 24036
rect 13860 23972 13924 24036
rect 24716 23972 24780 24036
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 5028 23836 5092 23900
rect 12756 23700 12820 23764
rect 2452 23564 2516 23628
rect 7604 23564 7668 23628
rect 16436 23564 16500 23628
rect 25452 23624 25516 23628
rect 25452 23568 25466 23624
rect 25466 23568 25516 23624
rect 25452 23564 25516 23568
rect 5948 23428 6012 23492
rect 12572 23488 12636 23492
rect 12572 23432 12622 23488
rect 12622 23432 12636 23488
rect 12572 23428 12636 23432
rect 20852 23488 20916 23492
rect 20852 23432 20902 23488
rect 20902 23432 20916 23488
rect 20852 23428 20916 23432
rect 25268 23488 25332 23492
rect 25268 23432 25282 23488
rect 25282 23432 25332 23488
rect 25268 23428 25332 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 12756 23292 12820 23356
rect 16252 23292 16316 23356
rect 26004 23020 26068 23084
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 9812 22748 9876 22812
rect 13492 22612 13556 22676
rect 18460 22748 18524 22812
rect 20668 22612 20732 22676
rect 9260 22340 9324 22404
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 3924 22204 3988 22268
rect 3740 22068 3804 22132
rect 12572 22068 12636 22132
rect 14596 22340 14660 22404
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 18460 22068 18524 22132
rect 18828 22128 18892 22132
rect 18828 22072 18878 22128
rect 18878 22072 18892 22128
rect 18828 22068 18892 22072
rect 19932 22128 19996 22132
rect 19932 22072 19982 22128
rect 19982 22072 19996 22128
rect 19932 22068 19996 22072
rect 1900 21660 1964 21724
rect 6500 21524 6564 21588
rect 7420 21932 7484 21996
rect 19196 21932 19260 21996
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 15148 21660 15212 21724
rect 18460 21796 18524 21860
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 20852 21524 20916 21588
rect 7420 21388 7484 21452
rect 8524 21312 8588 21316
rect 8524 21256 8574 21312
rect 8574 21256 8588 21312
rect 8524 21252 8588 21256
rect 21220 21252 21284 21316
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 12204 21116 12268 21180
rect 12020 21040 12084 21044
rect 12020 20984 12070 21040
rect 12070 20984 12084 21040
rect 12020 20980 12084 20984
rect 15884 20844 15948 20908
rect 8708 20768 8772 20772
rect 8708 20712 8758 20768
rect 8758 20712 8772 20768
rect 8708 20708 8772 20712
rect 9812 20708 9876 20772
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 13676 20708 13740 20772
rect 16804 20768 16868 20772
rect 16804 20712 16854 20768
rect 16854 20712 16868 20768
rect 16804 20708 16868 20712
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 24532 20980 24596 21044
rect 22508 20844 22572 20908
rect 21588 20708 21652 20772
rect 23612 20768 23676 20772
rect 23612 20712 23626 20768
rect 23626 20712 23676 20768
rect 23612 20708 23676 20712
rect 10180 20300 10244 20364
rect 17356 20436 17420 20500
rect 20668 20436 20732 20500
rect 16988 20300 17052 20364
rect 22324 20300 22388 20364
rect 11652 20224 11716 20228
rect 11652 20168 11702 20224
rect 11702 20168 11716 20224
rect 11652 20164 11716 20168
rect 19380 20224 19444 20228
rect 19380 20168 19394 20224
rect 19394 20168 19444 20224
rect 19380 20164 19444 20168
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 6684 19892 6748 19956
rect 10548 19892 10612 19956
rect 12572 20028 12636 20092
rect 23796 19952 23860 19956
rect 23796 19896 23810 19952
rect 23810 19896 23860 19952
rect 23796 19892 23860 19896
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 10364 19544 10428 19548
rect 21220 19620 21284 19684
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 10364 19488 10378 19544
rect 10378 19488 10428 19544
rect 10364 19484 10428 19488
rect 15700 19484 15764 19548
rect 12204 19348 12268 19412
rect 14044 19348 14108 19412
rect 15148 19348 15212 19412
rect 5580 19212 5644 19276
rect 6316 19212 6380 19276
rect 11836 19272 11900 19276
rect 11836 19216 11886 19272
rect 11886 19216 11900 19272
rect 11836 19212 11900 19216
rect 22140 19212 22204 19276
rect 23428 19348 23492 19412
rect 25636 19348 25700 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 10916 18940 10980 19004
rect 19932 19136 19996 19140
rect 19932 19080 19982 19136
rect 19982 19080 19996 19136
rect 19932 19076 19996 19080
rect 21404 19076 21468 19140
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 16436 18940 16500 19004
rect 17724 18940 17788 19004
rect 22692 18940 22756 19004
rect 16436 18804 16500 18868
rect 16068 18532 16132 18596
rect 19564 18532 19628 18596
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 5948 18396 6012 18460
rect 9076 18396 9140 18460
rect 20484 18396 20548 18460
rect 2268 18124 2332 18188
rect 9260 18124 9324 18188
rect 11284 18124 11348 18188
rect 15700 17988 15764 18052
rect 18460 18048 18524 18052
rect 18460 17992 18510 18048
rect 18510 17992 18524 18048
rect 18460 17988 18524 17992
rect 19748 18048 19812 18052
rect 19748 17992 19762 18048
rect 19762 17992 19812 18048
rect 19748 17988 19812 17992
rect 24716 17988 24780 18052
rect 24900 18048 24964 18052
rect 24900 17992 24950 18048
rect 24950 17992 24964 18048
rect 24900 17988 24964 17992
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 7788 17852 7852 17916
rect 8892 17852 8956 17916
rect 17172 17852 17236 17916
rect 21956 17716 22020 17780
rect 22140 17716 22204 17780
rect 9444 17444 9508 17508
rect 9996 17444 10060 17508
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 10548 17308 10612 17372
rect 8340 17036 8404 17100
rect 8340 16900 8404 16964
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 10732 16628 10796 16692
rect 22324 16764 22388 16828
rect 10180 16492 10244 16556
rect 15516 16628 15580 16692
rect 17724 16628 17788 16692
rect 14596 16492 14660 16556
rect 19196 16492 19260 16556
rect 20300 16492 20364 16556
rect 18828 16356 18892 16420
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 9444 16084 9508 16148
rect 12756 15948 12820 16012
rect 14044 15948 14108 16012
rect 14228 15948 14292 16012
rect 16252 15948 16316 16012
rect 9812 15812 9876 15876
rect 23428 15948 23492 16012
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 13860 15736 13924 15740
rect 13860 15680 13874 15736
rect 13874 15680 13924 15736
rect 13860 15676 13924 15680
rect 16252 15676 16316 15740
rect 16620 15736 16684 15740
rect 16620 15680 16634 15736
rect 16634 15680 16684 15736
rect 16620 15676 16684 15680
rect 5764 15540 5828 15604
rect 19012 15676 19076 15740
rect 20852 15676 20916 15740
rect 23980 15676 24044 15740
rect 9076 15464 9140 15468
rect 9076 15408 9126 15464
rect 9126 15408 9140 15464
rect 9076 15404 9140 15408
rect 9444 15464 9508 15468
rect 9444 15408 9494 15464
rect 9494 15408 9508 15464
rect 9444 15404 9508 15408
rect 20668 15404 20732 15468
rect 23428 15404 23492 15468
rect 9812 15268 9876 15332
rect 11284 15328 11348 15332
rect 11284 15272 11298 15328
rect 11298 15272 11348 15328
rect 11284 15268 11348 15272
rect 12020 15268 12084 15332
rect 20668 15268 20732 15332
rect 22140 15268 22204 15332
rect 25084 15268 25148 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 5028 15132 5092 15196
rect 10916 15132 10980 15196
rect 18644 15132 18708 15196
rect 26004 15132 26068 15196
rect 8340 14996 8404 15060
rect 15516 14996 15580 15060
rect 16804 14996 16868 15060
rect 18828 14996 18892 15060
rect 15148 14860 15212 14924
rect 17540 14724 17604 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 11468 14512 11532 14516
rect 11468 14456 11518 14512
rect 11518 14456 11532 14512
rect 11468 14452 11532 14456
rect 14412 14588 14476 14652
rect 16436 14588 16500 14652
rect 21772 14648 21836 14652
rect 21772 14592 21822 14648
rect 21822 14592 21836 14648
rect 21772 14588 21836 14592
rect 25084 14860 25148 14924
rect 17172 14452 17236 14516
rect 19380 14452 19444 14516
rect 21956 14316 22020 14380
rect 24348 14452 24412 14516
rect 13492 14180 13556 14244
rect 19012 14180 19076 14244
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 4108 13908 4172 13972
rect 11652 13908 11716 13972
rect 19564 14044 19628 14108
rect 16620 13772 16684 13836
rect 22324 13832 22388 13836
rect 22324 13776 22374 13832
rect 22374 13776 22388 13832
rect 22324 13772 22388 13776
rect 25820 13772 25884 13836
rect 19932 13636 19996 13700
rect 20116 13636 20180 13700
rect 21220 13636 21284 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 8892 13500 8956 13564
rect 9628 13500 9692 13564
rect 21588 13364 21652 13428
rect 16620 13228 16684 13292
rect 20484 13228 20548 13292
rect 23612 13228 23676 13292
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 6868 13016 6932 13020
rect 6868 12960 6918 13016
rect 6918 12960 6932 13016
rect 6868 12956 6932 12960
rect 23796 13092 23860 13156
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2452 12820 2516 12884
rect 16620 12956 16684 13020
rect 14228 12820 14292 12884
rect 17540 12820 17604 12884
rect 17724 12820 17788 12884
rect 21036 12956 21100 13020
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 6132 12412 6196 12476
rect 19012 12684 19076 12748
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 9996 12412 10060 12476
rect 12388 12472 12452 12476
rect 12388 12416 12402 12472
rect 12402 12416 12452 12472
rect 12388 12412 12452 12416
rect 18828 12608 18892 12612
rect 18828 12552 18878 12608
rect 18878 12552 18892 12608
rect 18828 12548 18892 12552
rect 24900 12548 24964 12612
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 6316 12276 6380 12340
rect 12572 12336 12636 12340
rect 12572 12280 12586 12336
rect 12586 12280 12636 12336
rect 12572 12276 12636 12280
rect 17540 12276 17604 12340
rect 19012 12276 19076 12340
rect 10548 12004 10612 12068
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 11468 11868 11532 11932
rect 5764 11732 5828 11796
rect 12756 12004 12820 12068
rect 16068 12004 16132 12068
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 23796 11868 23860 11932
rect 17724 11732 17788 11796
rect 19196 11732 19260 11796
rect 10732 11596 10796 11660
rect 3556 11460 3620 11524
rect 10364 11460 10428 11524
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 1900 11384 1964 11388
rect 1900 11328 1914 11384
rect 1914 11328 1964 11384
rect 1900 11324 1964 11328
rect 8524 11324 8588 11388
rect 6868 11248 6932 11252
rect 6868 11192 6918 11248
rect 6918 11192 6932 11248
rect 6868 11188 6932 11192
rect 19380 11596 19444 11660
rect 21220 11596 21284 11660
rect 25084 11596 25148 11660
rect 21772 11520 21836 11524
rect 21772 11464 21786 11520
rect 21786 11464 21836 11520
rect 21772 11460 21836 11464
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 15884 11188 15948 11252
rect 25452 11188 25516 11252
rect 4660 10916 4724 10980
rect 14780 11052 14844 11116
rect 16252 11052 16316 11116
rect 16436 11052 16500 11116
rect 18460 11052 18524 11116
rect 19196 11052 19260 11116
rect 20852 11052 20916 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 5580 10780 5644 10844
rect 7236 10780 7300 10844
rect 7788 10644 7852 10708
rect 16620 10780 16684 10844
rect 17172 10780 17236 10844
rect 13860 10644 13924 10708
rect 20116 10916 20180 10980
rect 22324 10916 22388 10980
rect 19380 10780 19444 10844
rect 21404 10780 21468 10844
rect 10916 10372 10980 10436
rect 22508 10644 22572 10708
rect 25636 10372 25700 10436
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7420 10100 7484 10164
rect 17540 10100 17604 10164
rect 18828 10100 18892 10164
rect 23980 10236 24044 10300
rect 24348 10236 24412 10300
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 13676 9692 13740 9756
rect 5212 9616 5276 9620
rect 5212 9560 5226 9616
rect 5226 9560 5276 9616
rect 5212 9556 5276 9560
rect 7604 9556 7668 9620
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 612 9148 676 9212
rect 16436 9420 16500 9484
rect 3924 9284 3988 9348
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 980 9012 1044 9076
rect 9812 9148 9876 9212
rect 12204 9012 12268 9076
rect 12572 9012 12636 9076
rect 3740 8876 3804 8940
rect 19380 8876 19444 8940
rect 2268 8740 2332 8804
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2636 8664 2700 8668
rect 2636 8608 2650 8664
rect 2650 8608 2700 8664
rect 2636 8604 2700 8608
rect 17172 8604 17236 8668
rect 796 8468 860 8532
rect 6684 8468 6748 8532
rect 22692 8332 22756 8396
rect 19012 8196 19076 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 9260 8060 9324 8124
rect 4108 7924 4172 7988
rect 25268 7788 25332 7852
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 26004 7380 26068 7444
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 15700 6836 15764 6900
rect 14412 6700 14476 6764
rect 15516 6700 15580 6764
rect 25820 6700 25884 6764
rect 19748 6564 19812 6628
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 16988 5944 17052 5948
rect 16988 5888 17002 5944
rect 17002 5888 17052 5944
rect 16988 5884 17052 5888
rect 6500 5748 6564 5812
rect 23428 5612 23492 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 20300 5204 20364 5268
rect 24532 5068 24596 5132
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 14596 4796 14660 4860
rect 8708 4524 8772 4588
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 17540 4312 17604 4316
rect 17540 4256 17554 4312
rect 17554 4256 17604 4312
rect 17540 4252 17604 4256
rect 25636 4116 25700 4180
rect 18644 3980 18708 4044
rect 20668 3980 20732 4044
rect 19196 3844 19260 3908
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 21956 3708 22020 3772
rect 21036 3572 21100 3636
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 11836 2892 11900 2956
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 24716 2484 24780 2548
rect 21220 2348 21284 2412
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 9259 26756 9325 26757
rect 9259 26692 9260 26756
rect 9324 26692 9325 26756
rect 9259 26691 9325 26692
rect 6131 26348 6197 26349
rect 6131 26284 6132 26348
rect 6196 26284 6197 26348
rect 6131 26283 6197 26284
rect 795 26212 861 26213
rect 795 26210 796 26212
rect 614 26150 796 26210
rect 614 9213 674 26150
rect 795 26148 796 26150
rect 860 26148 861 26212
rect 795 26147 861 26148
rect 5211 25940 5277 25941
rect 5211 25876 5212 25940
rect 5276 25876 5277 25940
rect 5211 25875 5277 25876
rect 795 25668 861 25669
rect 795 25604 796 25668
rect 860 25604 861 25668
rect 795 25603 861 25604
rect 611 9212 677 9213
rect 611 9148 612 9212
rect 676 9148 677 9212
rect 611 9147 677 9148
rect 798 8533 858 25603
rect 979 25532 1045 25533
rect 979 25468 980 25532
rect 1044 25468 1045 25532
rect 979 25467 1045 25468
rect 982 9077 1042 25467
rect 4659 25396 4725 25397
rect 4659 25332 4660 25396
rect 4724 25332 4725 25396
rect 4659 25331 4725 25332
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2635 24036 2701 24037
rect 2635 23972 2636 24036
rect 2700 23972 2701 24036
rect 2635 23971 2701 23972
rect 2451 23628 2517 23629
rect 2451 23564 2452 23628
rect 2516 23564 2517 23628
rect 2451 23563 2517 23564
rect 1899 21724 1965 21725
rect 1899 21660 1900 21724
rect 1964 21660 1965 21724
rect 1899 21659 1965 21660
rect 1902 11389 1962 21659
rect 2267 18188 2333 18189
rect 2267 18124 2268 18188
rect 2332 18124 2333 18188
rect 2267 18123 2333 18124
rect 1899 11388 1965 11389
rect 1899 11324 1900 11388
rect 1964 11324 1965 11388
rect 1899 11323 1965 11324
rect 979 9076 1045 9077
rect 979 9012 980 9076
rect 1044 9012 1045 9076
rect 979 9011 1045 9012
rect 2270 8805 2330 18123
rect 2454 12885 2514 23563
rect 2451 12884 2517 12885
rect 2451 12820 2452 12884
rect 2516 12820 2517 12884
rect 2451 12819 2517 12820
rect 2267 8804 2333 8805
rect 2267 8740 2268 8804
rect 2332 8740 2333 8804
rect 2267 8739 2333 8740
rect 2638 8669 2698 23971
rect 2944 23424 3264 24448
rect 3555 24172 3621 24173
rect 3555 24108 3556 24172
rect 3620 24108 3621 24172
rect 3555 24107 3621 24108
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 3558 11525 3618 24107
rect 3923 22268 3989 22269
rect 3923 22204 3924 22268
rect 3988 22204 3989 22268
rect 3923 22203 3989 22204
rect 3739 22132 3805 22133
rect 3739 22068 3740 22132
rect 3804 22068 3805 22132
rect 3739 22067 3805 22068
rect 3555 11524 3621 11525
rect 3555 11460 3556 11524
rect 3620 11460 3621 11524
rect 3555 11459 3621 11460
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2635 8668 2701 8669
rect 2635 8604 2636 8668
rect 2700 8604 2701 8668
rect 2635 8603 2701 8604
rect 795 8532 861 8533
rect 795 8468 796 8532
rect 860 8468 861 8532
rect 795 8467 861 8468
rect 2944 8192 3264 9216
rect 3742 8941 3802 22067
rect 3926 9349 3986 22203
rect 4107 13972 4173 13973
rect 4107 13908 4108 13972
rect 4172 13908 4173 13972
rect 4107 13907 4173 13908
rect 3923 9348 3989 9349
rect 3923 9284 3924 9348
rect 3988 9284 3989 9348
rect 3923 9283 3989 9284
rect 3739 8940 3805 8941
rect 3739 8876 3740 8940
rect 3804 8876 3805 8940
rect 3739 8875 3805 8876
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 4110 7989 4170 13907
rect 4662 10981 4722 25331
rect 5027 23900 5093 23901
rect 5027 23836 5028 23900
rect 5092 23836 5093 23900
rect 5027 23835 5093 23836
rect 5030 15197 5090 23835
rect 5027 15196 5093 15197
rect 5027 15132 5028 15196
rect 5092 15132 5093 15196
rect 5027 15131 5093 15132
rect 4659 10980 4725 10981
rect 4659 10916 4660 10980
rect 4724 10916 4725 10980
rect 4659 10915 4725 10916
rect 5214 9621 5274 25875
rect 5947 23492 6013 23493
rect 5947 23428 5948 23492
rect 6012 23428 6013 23492
rect 5947 23427 6013 23428
rect 5579 19276 5645 19277
rect 5579 19212 5580 19276
rect 5644 19212 5645 19276
rect 5579 19211 5645 19212
rect 5582 10845 5642 19211
rect 5950 18461 6010 23427
rect 5947 18460 6013 18461
rect 5947 18396 5948 18460
rect 6012 18396 6013 18460
rect 5947 18395 6013 18396
rect 5763 15604 5829 15605
rect 5763 15540 5764 15604
rect 5828 15540 5829 15604
rect 5763 15539 5829 15540
rect 5766 11797 5826 15539
rect 6134 12477 6194 26283
rect 8339 25396 8405 25397
rect 8339 25332 8340 25396
rect 8404 25332 8405 25396
rect 8339 25331 8405 25332
rect 7235 24444 7301 24445
rect 7235 24380 7236 24444
rect 7300 24380 7301 24444
rect 7235 24379 7301 24380
rect 6499 21588 6565 21589
rect 6499 21524 6500 21588
rect 6564 21524 6565 21588
rect 6499 21523 6565 21524
rect 6315 19276 6381 19277
rect 6315 19212 6316 19276
rect 6380 19212 6381 19276
rect 6315 19211 6381 19212
rect 6131 12476 6197 12477
rect 6131 12412 6132 12476
rect 6196 12412 6197 12476
rect 6131 12411 6197 12412
rect 6318 12341 6378 19211
rect 6315 12340 6381 12341
rect 6315 12276 6316 12340
rect 6380 12276 6381 12340
rect 6315 12275 6381 12276
rect 5763 11796 5829 11797
rect 5763 11732 5764 11796
rect 5828 11732 5829 11796
rect 5763 11731 5829 11732
rect 5579 10844 5645 10845
rect 5579 10780 5580 10844
rect 5644 10780 5645 10844
rect 5579 10779 5645 10780
rect 5211 9620 5277 9621
rect 5211 9556 5212 9620
rect 5276 9556 5277 9620
rect 5211 9555 5277 9556
rect 4107 7988 4173 7989
rect 4107 7924 4108 7988
rect 4172 7924 4173 7988
rect 4107 7923 4173 7924
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 6502 5813 6562 21523
rect 6683 19956 6749 19957
rect 6683 19892 6684 19956
rect 6748 19892 6749 19956
rect 6683 19891 6749 19892
rect 6686 8533 6746 19891
rect 6867 13020 6933 13021
rect 6867 12956 6868 13020
rect 6932 12956 6933 13020
rect 6867 12955 6933 12956
rect 6870 11253 6930 12955
rect 6867 11252 6933 11253
rect 6867 11188 6868 11252
rect 6932 11188 6933 11252
rect 6867 11187 6933 11188
rect 7238 10845 7298 24379
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7603 23628 7669 23629
rect 7603 23564 7604 23628
rect 7668 23564 7669 23628
rect 7603 23563 7669 23564
rect 7419 21996 7485 21997
rect 7419 21932 7420 21996
rect 7484 21932 7485 21996
rect 7419 21931 7485 21932
rect 7422 21453 7482 21931
rect 7419 21452 7485 21453
rect 7419 21388 7420 21452
rect 7484 21388 7485 21452
rect 7419 21387 7485 21388
rect 7235 10844 7301 10845
rect 7235 10780 7236 10844
rect 7300 10780 7301 10844
rect 7235 10779 7301 10780
rect 7422 10165 7482 21387
rect 7419 10164 7485 10165
rect 7419 10100 7420 10164
rect 7484 10100 7485 10164
rect 7419 10099 7485 10100
rect 7606 9621 7666 23563
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7787 17916 7853 17917
rect 7787 17852 7788 17916
rect 7852 17852 7853 17916
rect 7787 17851 7853 17852
rect 7790 10709 7850 17851
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 8342 17101 8402 25331
rect 9262 22405 9322 26691
rect 18459 26620 18525 26621
rect 18459 26556 18460 26620
rect 18524 26556 18525 26620
rect 18459 26555 18525 26556
rect 15147 25532 15213 25533
rect 15147 25468 15148 25532
rect 15212 25468 15213 25532
rect 15147 25467 15213 25468
rect 11099 25396 11165 25397
rect 11099 25332 11100 25396
rect 11164 25332 11165 25396
rect 11099 25331 11165 25332
rect 9443 25260 9509 25261
rect 9443 25196 9444 25260
rect 9508 25196 9509 25260
rect 9443 25195 9509 25196
rect 9259 22404 9325 22405
rect 9259 22340 9260 22404
rect 9324 22340 9325 22404
rect 9259 22339 9325 22340
rect 8523 21316 8589 21317
rect 8523 21252 8524 21316
rect 8588 21252 8589 21316
rect 8523 21251 8589 21252
rect 8339 17100 8405 17101
rect 8339 17036 8340 17100
rect 8404 17036 8405 17100
rect 8339 17035 8405 17036
rect 8339 16964 8405 16965
rect 8339 16900 8340 16964
rect 8404 16900 8405 16964
rect 8339 16899 8405 16900
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 8342 15061 8402 16899
rect 8339 15060 8405 15061
rect 8339 14996 8340 15060
rect 8404 14996 8405 15060
rect 8339 14995 8405 14996
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 8526 11389 8586 21251
rect 8707 20772 8773 20773
rect 8707 20708 8708 20772
rect 8772 20708 8773 20772
rect 8707 20707 8773 20708
rect 8523 11388 8589 11389
rect 8523 11324 8524 11388
rect 8588 11324 8589 11388
rect 8523 11323 8589 11324
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7787 10708 7853 10709
rect 7787 10644 7788 10708
rect 7852 10644 7853 10708
rect 7787 10643 7853 10644
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7603 9620 7669 9621
rect 7603 9556 7604 9620
rect 7668 9556 7669 9620
rect 7603 9555 7669 9556
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 6683 8532 6749 8533
rect 6683 8468 6684 8532
rect 6748 8468 6749 8532
rect 6683 8467 6749 8468
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 6499 5812 6565 5813
rect 6499 5748 6500 5812
rect 6564 5748 6565 5812
rect 6499 5747 6565 5748
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 8710 4589 8770 20707
rect 9075 18460 9141 18461
rect 9075 18396 9076 18460
rect 9140 18396 9141 18460
rect 9075 18395 9141 18396
rect 8891 17916 8957 17917
rect 8891 17852 8892 17916
rect 8956 17852 8957 17916
rect 8891 17851 8957 17852
rect 8894 13565 8954 17851
rect 9078 15469 9138 18395
rect 9259 18188 9325 18189
rect 9259 18124 9260 18188
rect 9324 18124 9325 18188
rect 9259 18123 9325 18124
rect 9075 15468 9141 15469
rect 9075 15404 9076 15468
rect 9140 15404 9141 15468
rect 9075 15403 9141 15404
rect 8891 13564 8957 13565
rect 8891 13500 8892 13564
rect 8956 13500 8957 13564
rect 8891 13499 8957 13500
rect 9262 8125 9322 18123
rect 9446 17509 9506 25195
rect 9811 25124 9877 25125
rect 9811 25060 9812 25124
rect 9876 25060 9877 25124
rect 9811 25059 9877 25060
rect 9627 24988 9693 24989
rect 9627 24924 9628 24988
rect 9692 24924 9693 24988
rect 9627 24923 9693 24924
rect 9443 17508 9509 17509
rect 9443 17444 9444 17508
rect 9508 17444 9509 17508
rect 9443 17443 9509 17444
rect 9443 16148 9509 16149
rect 9443 16084 9444 16148
rect 9508 16084 9509 16148
rect 9443 16083 9509 16084
rect 9446 15469 9506 16083
rect 9443 15468 9509 15469
rect 9443 15404 9444 15468
rect 9508 15404 9509 15468
rect 9443 15403 9509 15404
rect 9630 13565 9690 24923
rect 9814 22813 9874 25059
rect 10547 24852 10613 24853
rect 10547 24788 10548 24852
rect 10612 24788 10613 24852
rect 10547 24787 10613 24788
rect 9811 22812 9877 22813
rect 9811 22748 9812 22812
rect 9876 22748 9877 22812
rect 9811 22747 9877 22748
rect 9811 20772 9877 20773
rect 9811 20708 9812 20772
rect 9876 20708 9877 20772
rect 9811 20707 9877 20708
rect 9814 15877 9874 20707
rect 10179 20364 10245 20365
rect 10179 20300 10180 20364
rect 10244 20300 10245 20364
rect 10179 20299 10245 20300
rect 9995 17508 10061 17509
rect 9995 17444 9996 17508
rect 10060 17444 10061 17508
rect 9995 17443 10061 17444
rect 9811 15876 9877 15877
rect 9811 15812 9812 15876
rect 9876 15812 9877 15876
rect 9811 15811 9877 15812
rect 9811 15332 9877 15333
rect 9811 15268 9812 15332
rect 9876 15268 9877 15332
rect 9811 15267 9877 15268
rect 9627 13564 9693 13565
rect 9627 13500 9628 13564
rect 9692 13500 9693 13564
rect 9627 13499 9693 13500
rect 9814 9213 9874 15267
rect 9998 12477 10058 17443
rect 10182 16557 10242 20299
rect 10550 19957 10610 24787
rect 10547 19956 10613 19957
rect 10547 19892 10548 19956
rect 10612 19892 10613 19956
rect 10547 19891 10613 19892
rect 10363 19548 10429 19549
rect 10363 19484 10364 19548
rect 10428 19484 10429 19548
rect 10363 19483 10429 19484
rect 10179 16556 10245 16557
rect 10179 16492 10180 16556
rect 10244 16492 10245 16556
rect 10179 16491 10245 16492
rect 9995 12476 10061 12477
rect 9995 12412 9996 12476
rect 10060 12412 10061 12476
rect 9995 12411 10061 12412
rect 10366 11525 10426 19483
rect 11102 19410 11162 25331
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 11651 24172 11717 24173
rect 11651 24108 11652 24172
rect 11716 24108 11717 24172
rect 11651 24107 11717 24108
rect 11654 20229 11714 24107
rect 12203 24036 12269 24037
rect 12203 23972 12204 24036
rect 12268 23972 12269 24036
rect 12203 23971 12269 23972
rect 12206 21181 12266 23971
rect 12755 23764 12821 23765
rect 12755 23700 12756 23764
rect 12820 23700 12821 23764
rect 12755 23699 12821 23700
rect 12571 23492 12637 23493
rect 12571 23428 12572 23492
rect 12636 23428 12637 23492
rect 12571 23427 12637 23428
rect 12574 22133 12634 23427
rect 12758 23357 12818 23699
rect 12944 23424 13264 24448
rect 13859 24036 13925 24037
rect 13859 23972 13860 24036
rect 13924 23972 13925 24036
rect 13859 23971 13925 23972
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12755 23356 12821 23357
rect 12755 23292 12756 23356
rect 12820 23292 12821 23356
rect 12755 23291 12821 23292
rect 12944 22336 13264 23360
rect 13491 22676 13557 22677
rect 13491 22612 13492 22676
rect 13556 22612 13557 22676
rect 13491 22611 13557 22612
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12571 22132 12637 22133
rect 12571 22068 12572 22132
rect 12636 22068 12637 22132
rect 12571 22067 12637 22068
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12203 21180 12269 21181
rect 12203 21116 12204 21180
rect 12268 21116 12269 21180
rect 12203 21115 12269 21116
rect 12019 21044 12085 21045
rect 12019 20980 12020 21044
rect 12084 20980 12085 21044
rect 12019 20979 12085 20980
rect 11651 20228 11717 20229
rect 11651 20164 11652 20228
rect 11716 20164 11717 20228
rect 11651 20163 11717 20164
rect 10918 19350 11162 19410
rect 10918 19005 10978 19350
rect 10915 19004 10981 19005
rect 10915 18940 10916 19004
rect 10980 18940 10981 19004
rect 10915 18939 10981 18940
rect 11283 18188 11349 18189
rect 11283 18124 11284 18188
rect 11348 18124 11349 18188
rect 11283 18123 11349 18124
rect 10547 17372 10613 17373
rect 10547 17308 10548 17372
rect 10612 17308 10613 17372
rect 10547 17307 10613 17308
rect 10550 12069 10610 17307
rect 10731 16692 10797 16693
rect 10731 16628 10732 16692
rect 10796 16628 10797 16692
rect 10731 16627 10797 16628
rect 10547 12068 10613 12069
rect 10547 12004 10548 12068
rect 10612 12004 10613 12068
rect 10547 12003 10613 12004
rect 10734 11661 10794 16627
rect 11286 15333 11346 18123
rect 11283 15332 11349 15333
rect 11283 15268 11284 15332
rect 11348 15268 11349 15332
rect 11283 15267 11349 15268
rect 10915 15196 10981 15197
rect 10915 15132 10916 15196
rect 10980 15132 10981 15196
rect 10915 15131 10981 15132
rect 10731 11660 10797 11661
rect 10731 11596 10732 11660
rect 10796 11596 10797 11660
rect 10731 11595 10797 11596
rect 10363 11524 10429 11525
rect 10363 11460 10364 11524
rect 10428 11460 10429 11524
rect 10363 11459 10429 11460
rect 10918 10437 10978 15131
rect 11467 14516 11533 14517
rect 11467 14452 11468 14516
rect 11532 14452 11533 14516
rect 11467 14451 11533 14452
rect 11470 11933 11530 14451
rect 11654 13973 11714 20163
rect 11835 19276 11901 19277
rect 11835 19212 11836 19276
rect 11900 19212 11901 19276
rect 11835 19211 11901 19212
rect 11651 13972 11717 13973
rect 11651 13908 11652 13972
rect 11716 13908 11717 13972
rect 11651 13907 11717 13908
rect 11467 11932 11533 11933
rect 11467 11868 11468 11932
rect 11532 11868 11533 11932
rect 11467 11867 11533 11868
rect 10915 10436 10981 10437
rect 10915 10372 10916 10436
rect 10980 10372 10981 10436
rect 10915 10371 10981 10372
rect 9811 9212 9877 9213
rect 9811 9148 9812 9212
rect 9876 9148 9877 9212
rect 9811 9147 9877 9148
rect 9259 8124 9325 8125
rect 9259 8060 9260 8124
rect 9324 8060 9325 8124
rect 9259 8059 9325 8060
rect 8707 4588 8773 4589
rect 8707 4524 8708 4588
rect 8772 4524 8773 4588
rect 8707 4523 8773 4524
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 11838 2957 11898 19211
rect 12022 15333 12082 20979
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12571 20092 12637 20093
rect 12571 20028 12572 20092
rect 12636 20028 12637 20092
rect 12571 20027 12637 20028
rect 12203 19412 12269 19413
rect 12203 19348 12204 19412
rect 12268 19348 12269 19412
rect 12203 19347 12269 19348
rect 12019 15332 12085 15333
rect 12019 15268 12020 15332
rect 12084 15268 12085 15332
rect 12019 15267 12085 15268
rect 12206 9077 12266 19347
rect 12387 12476 12453 12477
rect 12387 12412 12388 12476
rect 12452 12412 12453 12476
rect 12387 12411 12453 12412
rect 12390 11930 12450 12411
rect 12574 12341 12634 20027
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12755 16012 12821 16013
rect 12755 15948 12756 16012
rect 12820 15948 12821 16012
rect 12755 15947 12821 15948
rect 12571 12340 12637 12341
rect 12571 12276 12572 12340
rect 12636 12276 12637 12340
rect 12571 12275 12637 12276
rect 12758 12069 12818 15947
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 13494 14245 13554 22611
rect 13675 20772 13741 20773
rect 13675 20708 13676 20772
rect 13740 20708 13741 20772
rect 13675 20707 13741 20708
rect 13491 14244 13557 14245
rect 13491 14180 13492 14244
rect 13556 14180 13557 14244
rect 13491 14179 13557 14180
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12755 12068 12821 12069
rect 12755 12004 12756 12068
rect 12820 12004 12821 12068
rect 12755 12003 12821 12004
rect 12390 11870 12634 11930
rect 12574 9077 12634 11870
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 13678 9757 13738 20707
rect 13862 15741 13922 23971
rect 14595 22404 14661 22405
rect 14595 22340 14596 22404
rect 14660 22340 14661 22404
rect 14595 22339 14661 22340
rect 14043 19412 14109 19413
rect 14043 19348 14044 19412
rect 14108 19348 14109 19412
rect 14043 19347 14109 19348
rect 14598 19350 14658 22339
rect 15150 21725 15210 25467
rect 16619 24172 16685 24173
rect 16619 24108 16620 24172
rect 16684 24108 16685 24172
rect 16619 24107 16685 24108
rect 16435 23628 16501 23629
rect 16435 23564 16436 23628
rect 16500 23564 16501 23628
rect 16435 23563 16501 23564
rect 16251 23356 16317 23357
rect 16251 23292 16252 23356
rect 16316 23292 16317 23356
rect 16251 23291 16317 23292
rect 15147 21724 15213 21725
rect 15147 21660 15148 21724
rect 15212 21660 15213 21724
rect 15147 21659 15213 21660
rect 15883 20908 15949 20909
rect 15883 20844 15884 20908
rect 15948 20844 15949 20908
rect 15883 20843 15949 20844
rect 15699 19548 15765 19549
rect 15699 19484 15700 19548
rect 15764 19484 15765 19548
rect 15699 19483 15765 19484
rect 15147 19412 15213 19413
rect 14046 16013 14106 19347
rect 14598 19290 14842 19350
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 14595 16556 14661 16557
rect 14595 16492 14596 16556
rect 14660 16492 14661 16556
rect 14595 16491 14661 16492
rect 14043 16012 14109 16013
rect 14043 15948 14044 16012
rect 14108 15948 14109 16012
rect 14043 15947 14109 15948
rect 14227 16012 14293 16013
rect 14227 15948 14228 16012
rect 14292 15948 14293 16012
rect 14227 15947 14293 15948
rect 13859 15740 13925 15741
rect 13859 15676 13860 15740
rect 13924 15676 13925 15740
rect 13859 15675 13925 15676
rect 13862 10709 13922 15675
rect 14230 12885 14290 15947
rect 14411 14652 14477 14653
rect 14411 14588 14412 14652
rect 14476 14588 14477 14652
rect 14411 14587 14477 14588
rect 14227 12884 14293 12885
rect 14227 12820 14228 12884
rect 14292 12820 14293 12884
rect 14227 12819 14293 12820
rect 13859 10708 13925 10709
rect 13859 10644 13860 10708
rect 13924 10644 13925 10708
rect 13859 10643 13925 10644
rect 13675 9756 13741 9757
rect 13675 9692 13676 9756
rect 13740 9692 13741 9756
rect 13675 9691 13741 9692
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12203 9076 12269 9077
rect 12203 9012 12204 9076
rect 12268 9012 12269 9076
rect 12203 9011 12269 9012
rect 12571 9076 12637 9077
rect 12571 9012 12572 9076
rect 12636 9012 12637 9076
rect 12571 9011 12637 9012
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 14414 6765 14474 14587
rect 14411 6764 14477 6765
rect 14411 6700 14412 6764
rect 14476 6700 14477 6764
rect 14411 6699 14477 6700
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 14598 4861 14658 16491
rect 14782 11117 14842 19290
rect 15150 14925 15210 19347
rect 15702 18730 15762 19483
rect 15518 18670 15762 18730
rect 15518 16693 15578 18670
rect 15699 18052 15765 18053
rect 15699 17988 15700 18052
rect 15764 17988 15765 18052
rect 15699 17987 15765 17988
rect 15515 16692 15581 16693
rect 15515 16628 15516 16692
rect 15580 16628 15581 16692
rect 15515 16627 15581 16628
rect 15515 15060 15581 15061
rect 15515 14996 15516 15060
rect 15580 14996 15581 15060
rect 15515 14995 15581 14996
rect 15147 14924 15213 14925
rect 15147 14860 15148 14924
rect 15212 14860 15213 14924
rect 15147 14859 15213 14860
rect 14779 11116 14845 11117
rect 14779 11052 14780 11116
rect 14844 11052 14845 11116
rect 14779 11051 14845 11052
rect 15518 6765 15578 14995
rect 15702 6901 15762 17987
rect 15886 11253 15946 20843
rect 16067 18596 16133 18597
rect 16067 18532 16068 18596
rect 16132 18532 16133 18596
rect 16067 18531 16133 18532
rect 16070 12069 16130 18531
rect 16254 16013 16314 23291
rect 16438 19005 16498 23563
rect 16435 19004 16501 19005
rect 16435 18940 16436 19004
rect 16500 18940 16501 19004
rect 16435 18939 16501 18940
rect 16435 18868 16501 18869
rect 16435 18804 16436 18868
rect 16500 18804 16501 18868
rect 16435 18803 16501 18804
rect 16251 16012 16317 16013
rect 16251 15948 16252 16012
rect 16316 15948 16317 16012
rect 16251 15947 16317 15948
rect 16251 15740 16317 15741
rect 16251 15676 16252 15740
rect 16316 15676 16317 15740
rect 16251 15675 16317 15676
rect 16067 12068 16133 12069
rect 16067 12004 16068 12068
rect 16132 12004 16133 12068
rect 16067 12003 16133 12004
rect 15883 11252 15949 11253
rect 15883 11188 15884 11252
rect 15948 11188 15949 11252
rect 15883 11187 15949 11188
rect 16254 11117 16314 15675
rect 16438 14653 16498 18803
rect 16622 15741 16682 24107
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 18462 22813 18522 26555
rect 18827 26484 18893 26485
rect 18827 26420 18828 26484
rect 18892 26420 18893 26484
rect 18827 26419 18893 26420
rect 18459 22812 18525 22813
rect 18459 22748 18460 22812
rect 18524 22748 18525 22812
rect 18459 22747 18525 22748
rect 18830 22133 18890 26419
rect 20667 25124 20733 25125
rect 20667 25060 20668 25124
rect 20732 25060 20733 25124
rect 20667 25059 20733 25060
rect 19011 24308 19077 24309
rect 19011 24244 19012 24308
rect 19076 24244 19077 24308
rect 19011 24243 19077 24244
rect 18459 22132 18525 22133
rect 18459 22068 18460 22132
rect 18524 22068 18525 22132
rect 18459 22067 18525 22068
rect 18827 22132 18893 22133
rect 18827 22068 18828 22132
rect 18892 22068 18893 22132
rect 18827 22067 18893 22068
rect 18462 21861 18522 22067
rect 18459 21860 18525 21861
rect 18459 21796 18460 21860
rect 18524 21796 18525 21860
rect 18459 21795 18525 21796
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 16803 20772 16869 20773
rect 16803 20708 16804 20772
rect 16868 20708 16869 20772
rect 16803 20707 16869 20708
rect 16619 15740 16685 15741
rect 16619 15676 16620 15740
rect 16684 15676 16685 15740
rect 16619 15675 16685 15676
rect 16806 15061 16866 20707
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17355 20500 17421 20501
rect 17355 20436 17356 20500
rect 17420 20436 17421 20500
rect 17355 20435 17421 20436
rect 16987 20364 17053 20365
rect 16987 20300 16988 20364
rect 17052 20300 17053 20364
rect 16987 20299 17053 20300
rect 16803 15060 16869 15061
rect 16803 14996 16804 15060
rect 16868 14996 16869 15060
rect 16803 14995 16869 14996
rect 16435 14652 16501 14653
rect 16435 14588 16436 14652
rect 16500 14588 16501 14652
rect 16435 14587 16501 14588
rect 16619 13836 16685 13837
rect 16619 13772 16620 13836
rect 16684 13772 16685 13836
rect 16619 13771 16685 13772
rect 16622 13293 16682 13771
rect 16619 13292 16685 13293
rect 16619 13228 16620 13292
rect 16684 13228 16685 13292
rect 16619 13227 16685 13228
rect 16619 13020 16685 13021
rect 16619 12956 16620 13020
rect 16684 12956 16685 13020
rect 16619 12955 16685 12956
rect 16251 11116 16317 11117
rect 16251 11052 16252 11116
rect 16316 11052 16317 11116
rect 16251 11051 16317 11052
rect 16435 11116 16501 11117
rect 16435 11052 16436 11116
rect 16500 11052 16501 11116
rect 16435 11051 16501 11052
rect 16438 9485 16498 11051
rect 16622 10845 16682 12955
rect 16619 10844 16685 10845
rect 16619 10780 16620 10844
rect 16684 10780 16685 10844
rect 16619 10779 16685 10780
rect 16435 9484 16501 9485
rect 16435 9420 16436 9484
rect 16500 9420 16501 9484
rect 16435 9419 16501 9420
rect 15699 6900 15765 6901
rect 15699 6836 15700 6900
rect 15764 6836 15765 6900
rect 15699 6835 15765 6836
rect 15515 6764 15581 6765
rect 15515 6700 15516 6764
rect 15580 6700 15581 6764
rect 15515 6699 15581 6700
rect 16990 5949 17050 20299
rect 17171 17916 17237 17917
rect 17171 17852 17172 17916
rect 17236 17852 17237 17916
rect 17171 17851 17237 17852
rect 17174 14517 17234 17851
rect 17171 14516 17237 14517
rect 17171 14452 17172 14516
rect 17236 14452 17237 14516
rect 17171 14451 17237 14452
rect 17358 12746 17418 20435
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17723 19004 17789 19005
rect 17723 18940 17724 19004
rect 17788 18940 17789 19004
rect 17723 18939 17789 18940
rect 17726 16693 17786 18939
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 18459 18052 18525 18053
rect 18459 17988 18460 18052
rect 18524 17988 18525 18052
rect 18459 17987 18525 17988
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17723 16692 17789 16693
rect 17723 16628 17724 16692
rect 17788 16628 17789 16692
rect 17723 16627 17789 16628
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17539 14788 17605 14789
rect 17539 14724 17540 14788
rect 17604 14724 17605 14788
rect 17539 14723 17605 14724
rect 17542 12885 17602 14723
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17539 12884 17605 12885
rect 17539 12820 17540 12884
rect 17604 12820 17605 12884
rect 17539 12819 17605 12820
rect 17723 12884 17789 12885
rect 17723 12820 17724 12884
rect 17788 12820 17789 12884
rect 17723 12819 17789 12820
rect 17358 12686 17602 12746
rect 17542 12341 17602 12686
rect 17539 12340 17605 12341
rect 17539 12276 17540 12340
rect 17604 12276 17605 12340
rect 17539 12275 17605 12276
rect 17726 11797 17786 12819
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17723 11796 17789 11797
rect 17723 11732 17724 11796
rect 17788 11732 17789 11796
rect 17723 11731 17789 11732
rect 17944 10912 18264 11936
rect 18462 11117 18522 17987
rect 18827 16420 18893 16421
rect 18827 16356 18828 16420
rect 18892 16356 18893 16420
rect 18827 16355 18893 16356
rect 18643 15196 18709 15197
rect 18643 15132 18644 15196
rect 18708 15132 18709 15196
rect 18643 15131 18709 15132
rect 18459 11116 18525 11117
rect 18459 11052 18460 11116
rect 18524 11052 18525 11116
rect 18459 11051 18525 11052
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17171 10844 17237 10845
rect 17171 10780 17172 10844
rect 17236 10780 17237 10844
rect 17171 10779 17237 10780
rect 17174 8669 17234 10779
rect 17539 10164 17605 10165
rect 17539 10100 17540 10164
rect 17604 10100 17605 10164
rect 17539 10099 17605 10100
rect 17171 8668 17237 8669
rect 17171 8604 17172 8668
rect 17236 8604 17237 8668
rect 17171 8603 17237 8604
rect 16987 5948 17053 5949
rect 16987 5884 16988 5948
rect 17052 5884 17053 5948
rect 16987 5883 17053 5884
rect 14595 4860 14661 4861
rect 14595 4796 14596 4860
rect 14660 4796 14661 4860
rect 14595 4795 14661 4796
rect 17542 4317 17602 10099
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17539 4316 17605 4317
rect 17539 4252 17540 4316
rect 17604 4252 17605 4316
rect 17539 4251 17605 4252
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 11835 2956 11901 2957
rect 11835 2892 11836 2956
rect 11900 2892 11901 2956
rect 11835 2891 11901 2892
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 3296 18264 4320
rect 18646 4045 18706 15131
rect 18830 15061 18890 16355
rect 19014 15741 19074 24243
rect 20670 22677 20730 25059
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 20851 23492 20917 23493
rect 20851 23428 20852 23492
rect 20916 23428 20917 23492
rect 20851 23427 20917 23428
rect 20667 22676 20733 22677
rect 20667 22612 20668 22676
rect 20732 22612 20733 22676
rect 20667 22611 20733 22612
rect 19931 22132 19997 22133
rect 19931 22068 19932 22132
rect 19996 22068 19997 22132
rect 19931 22067 19997 22068
rect 19195 21996 19261 21997
rect 19195 21932 19196 21996
rect 19260 21932 19261 21996
rect 19195 21931 19261 21932
rect 19198 16557 19258 21931
rect 19379 20228 19445 20229
rect 19379 20164 19380 20228
rect 19444 20164 19445 20228
rect 19379 20163 19445 20164
rect 19195 16556 19261 16557
rect 19195 16492 19196 16556
rect 19260 16492 19261 16556
rect 19195 16491 19261 16492
rect 19382 16010 19442 20163
rect 19934 19141 19994 22067
rect 20854 21589 20914 23427
rect 22944 23424 23264 24448
rect 24715 24036 24781 24037
rect 24715 23972 24716 24036
rect 24780 23972 24781 24036
rect 24715 23971 24781 23972
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 20851 21588 20917 21589
rect 20851 21524 20852 21588
rect 20916 21524 20917 21588
rect 20851 21523 20917 21524
rect 21219 21316 21285 21317
rect 21219 21252 21220 21316
rect 21284 21252 21285 21316
rect 21219 21251 21285 21252
rect 20667 20500 20733 20501
rect 20667 20436 20668 20500
rect 20732 20436 20733 20500
rect 20667 20435 20733 20436
rect 19931 19140 19997 19141
rect 19931 19076 19932 19140
rect 19996 19076 19997 19140
rect 19931 19075 19997 19076
rect 19563 18596 19629 18597
rect 19563 18532 19564 18596
rect 19628 18532 19629 18596
rect 19563 18531 19629 18532
rect 19198 15950 19442 16010
rect 19011 15740 19077 15741
rect 19011 15676 19012 15740
rect 19076 15676 19077 15740
rect 19011 15675 19077 15676
rect 18827 15060 18893 15061
rect 18827 14996 18828 15060
rect 18892 14996 18893 15060
rect 18827 14995 18893 14996
rect 19011 14244 19077 14245
rect 19011 14180 19012 14244
rect 19076 14180 19077 14244
rect 19011 14179 19077 14180
rect 19014 12749 19074 14179
rect 19011 12748 19077 12749
rect 19011 12684 19012 12748
rect 19076 12684 19077 12748
rect 19011 12683 19077 12684
rect 18827 12612 18893 12613
rect 18827 12548 18828 12612
rect 18892 12548 18893 12612
rect 18827 12547 18893 12548
rect 18830 10165 18890 12547
rect 19011 12340 19077 12341
rect 19011 12276 19012 12340
rect 19076 12276 19077 12340
rect 19011 12275 19077 12276
rect 18827 10164 18893 10165
rect 18827 10100 18828 10164
rect 18892 10100 18893 10164
rect 18827 10099 18893 10100
rect 19014 8261 19074 12275
rect 19198 11797 19258 15950
rect 19379 14516 19445 14517
rect 19379 14452 19380 14516
rect 19444 14452 19445 14516
rect 19379 14451 19445 14452
rect 19195 11796 19261 11797
rect 19195 11732 19196 11796
rect 19260 11732 19261 11796
rect 19195 11731 19261 11732
rect 19382 11661 19442 14451
rect 19566 14109 19626 18531
rect 19747 18052 19813 18053
rect 19747 17988 19748 18052
rect 19812 17988 19813 18052
rect 19747 17987 19813 17988
rect 19563 14108 19629 14109
rect 19563 14044 19564 14108
rect 19628 14044 19629 14108
rect 19563 14043 19629 14044
rect 19379 11660 19445 11661
rect 19379 11596 19380 11660
rect 19444 11596 19445 11660
rect 19379 11595 19445 11596
rect 19195 11116 19261 11117
rect 19195 11052 19196 11116
rect 19260 11052 19261 11116
rect 19195 11051 19261 11052
rect 19011 8260 19077 8261
rect 19011 8196 19012 8260
rect 19076 8196 19077 8260
rect 19011 8195 19077 8196
rect 18643 4044 18709 4045
rect 18643 3980 18644 4044
rect 18708 3980 18709 4044
rect 18643 3979 18709 3980
rect 19198 3909 19258 11051
rect 19379 10844 19445 10845
rect 19379 10780 19380 10844
rect 19444 10780 19445 10844
rect 19379 10779 19445 10780
rect 19382 8941 19442 10779
rect 19379 8940 19445 8941
rect 19379 8876 19380 8940
rect 19444 8876 19445 8940
rect 19379 8875 19445 8876
rect 19750 6629 19810 17987
rect 19934 13701 19994 19075
rect 20483 18460 20549 18461
rect 20483 18396 20484 18460
rect 20548 18396 20549 18460
rect 20483 18395 20549 18396
rect 20299 16556 20365 16557
rect 20299 16492 20300 16556
rect 20364 16492 20365 16556
rect 20299 16491 20365 16492
rect 19931 13700 19997 13701
rect 19931 13636 19932 13700
rect 19996 13636 19997 13700
rect 19931 13635 19997 13636
rect 20115 13700 20181 13701
rect 20115 13636 20116 13700
rect 20180 13636 20181 13700
rect 20115 13635 20181 13636
rect 20118 10981 20178 13635
rect 20115 10980 20181 10981
rect 20115 10916 20116 10980
rect 20180 10916 20181 10980
rect 20115 10915 20181 10916
rect 19747 6628 19813 6629
rect 19747 6564 19748 6628
rect 19812 6564 19813 6628
rect 19747 6563 19813 6564
rect 20302 5269 20362 16491
rect 20486 13293 20546 18395
rect 20670 15469 20730 20435
rect 21222 19685 21282 21251
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22507 20908 22573 20909
rect 22507 20844 22508 20908
rect 22572 20844 22573 20908
rect 22507 20843 22573 20844
rect 21587 20772 21653 20773
rect 21587 20708 21588 20772
rect 21652 20708 21653 20772
rect 21587 20707 21653 20708
rect 21219 19684 21285 19685
rect 21219 19620 21220 19684
rect 21284 19620 21285 19684
rect 21219 19619 21285 19620
rect 20851 15740 20917 15741
rect 20851 15676 20852 15740
rect 20916 15676 20917 15740
rect 20851 15675 20917 15676
rect 20667 15468 20733 15469
rect 20667 15404 20668 15468
rect 20732 15404 20733 15468
rect 20667 15403 20733 15404
rect 20667 15332 20733 15333
rect 20667 15268 20668 15332
rect 20732 15268 20733 15332
rect 20667 15267 20733 15268
rect 20483 13292 20549 13293
rect 20483 13228 20484 13292
rect 20548 13228 20549 13292
rect 20483 13227 20549 13228
rect 20299 5268 20365 5269
rect 20299 5204 20300 5268
rect 20364 5204 20365 5268
rect 20299 5203 20365 5204
rect 20670 4045 20730 15267
rect 20854 11117 20914 15675
rect 21222 13701 21282 19619
rect 21403 19140 21469 19141
rect 21403 19076 21404 19140
rect 21468 19076 21469 19140
rect 21403 19075 21469 19076
rect 21219 13700 21285 13701
rect 21219 13636 21220 13700
rect 21284 13636 21285 13700
rect 21219 13635 21285 13636
rect 21035 13020 21101 13021
rect 21035 12956 21036 13020
rect 21100 12956 21101 13020
rect 21035 12955 21101 12956
rect 20851 11116 20917 11117
rect 20851 11052 20852 11116
rect 20916 11052 20917 11116
rect 20851 11051 20917 11052
rect 20667 4044 20733 4045
rect 20667 3980 20668 4044
rect 20732 3980 20733 4044
rect 20667 3979 20733 3980
rect 19195 3908 19261 3909
rect 19195 3844 19196 3908
rect 19260 3844 19261 3908
rect 19195 3843 19261 3844
rect 21038 3637 21098 12955
rect 21219 11660 21285 11661
rect 21219 11596 21220 11660
rect 21284 11596 21285 11660
rect 21219 11595 21285 11596
rect 21035 3636 21101 3637
rect 21035 3572 21036 3636
rect 21100 3572 21101 3636
rect 21035 3571 21101 3572
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 21222 2413 21282 11595
rect 21406 10845 21466 19075
rect 21590 13429 21650 20707
rect 22323 20364 22389 20365
rect 22323 20300 22324 20364
rect 22388 20300 22389 20364
rect 22323 20299 22389 20300
rect 22139 19276 22205 19277
rect 22139 19212 22140 19276
rect 22204 19212 22205 19276
rect 22139 19211 22205 19212
rect 22142 17781 22202 19211
rect 21955 17780 22021 17781
rect 21955 17716 21956 17780
rect 22020 17716 22021 17780
rect 21955 17715 22021 17716
rect 22139 17780 22205 17781
rect 22139 17716 22140 17780
rect 22204 17716 22205 17780
rect 22139 17715 22205 17716
rect 21771 14652 21837 14653
rect 21771 14588 21772 14652
rect 21836 14588 21837 14652
rect 21771 14587 21837 14588
rect 21587 13428 21653 13429
rect 21587 13364 21588 13428
rect 21652 13364 21653 13428
rect 21587 13363 21653 13364
rect 21774 11525 21834 14587
rect 21958 14381 22018 17715
rect 22326 16829 22386 20299
rect 22323 16828 22389 16829
rect 22323 16764 22324 16828
rect 22388 16764 22389 16828
rect 22323 16763 22389 16764
rect 22139 15332 22205 15333
rect 22139 15268 22140 15332
rect 22204 15268 22205 15332
rect 22139 15267 22205 15268
rect 21955 14380 22021 14381
rect 21955 14316 21956 14380
rect 22020 14316 22021 14380
rect 21955 14315 22021 14316
rect 21771 11524 21837 11525
rect 21771 11460 21772 11524
rect 21836 11460 21837 11524
rect 22142 11522 22202 15267
rect 22323 13836 22389 13837
rect 22323 13772 22324 13836
rect 22388 13772 22389 13836
rect 22323 13771 22389 13772
rect 21771 11459 21837 11460
rect 21958 11462 22202 11522
rect 21403 10844 21469 10845
rect 21403 10780 21404 10844
rect 21468 10780 21469 10844
rect 21403 10779 21469 10780
rect 21958 3773 22018 11462
rect 22326 10981 22386 13771
rect 22323 10980 22389 10981
rect 22323 10916 22324 10980
rect 22388 10916 22389 10980
rect 22323 10915 22389 10916
rect 22510 10709 22570 20843
rect 22944 20160 23264 21184
rect 24531 21044 24597 21045
rect 24531 20980 24532 21044
rect 24596 20980 24597 21044
rect 24531 20979 24597 20980
rect 23611 20772 23677 20773
rect 23611 20708 23612 20772
rect 23676 20708 23677 20772
rect 23611 20707 23677 20708
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 23427 19412 23493 19413
rect 23427 19348 23428 19412
rect 23492 19348 23493 19412
rect 23427 19347 23493 19348
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22691 19004 22757 19005
rect 22691 18940 22692 19004
rect 22756 18940 22757 19004
rect 22691 18939 22757 18940
rect 22507 10708 22573 10709
rect 22507 10644 22508 10708
rect 22572 10644 22573 10708
rect 22507 10643 22573 10644
rect 22694 8397 22754 18939
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 23430 16013 23490 19347
rect 23427 16012 23493 16013
rect 23427 15948 23428 16012
rect 23492 15948 23493 16012
rect 23427 15947 23493 15948
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 23427 15468 23493 15469
rect 23427 15404 23428 15468
rect 23492 15404 23493 15468
rect 23427 15403 23493 15404
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22691 8396 22757 8397
rect 22691 8332 22692 8396
rect 22756 8332 22757 8396
rect 22691 8331 22757 8332
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 23430 5677 23490 15403
rect 23614 13293 23674 20707
rect 23795 19956 23861 19957
rect 23795 19892 23796 19956
rect 23860 19892 23861 19956
rect 23795 19891 23861 19892
rect 23611 13292 23677 13293
rect 23611 13228 23612 13292
rect 23676 13228 23677 13292
rect 23611 13227 23677 13228
rect 23798 13157 23858 19891
rect 23979 15740 24045 15741
rect 23979 15676 23980 15740
rect 24044 15676 24045 15740
rect 23979 15675 24045 15676
rect 23795 13156 23861 13157
rect 23795 13092 23796 13156
rect 23860 13092 23861 13156
rect 23795 13091 23861 13092
rect 23798 11933 23858 13091
rect 23795 11932 23861 11933
rect 23795 11868 23796 11932
rect 23860 11868 23861 11932
rect 23795 11867 23861 11868
rect 23982 10301 24042 15675
rect 24347 14516 24413 14517
rect 24347 14452 24348 14516
rect 24412 14452 24413 14516
rect 24347 14451 24413 14452
rect 24350 10301 24410 14451
rect 23979 10300 24045 10301
rect 23979 10236 23980 10300
rect 24044 10236 24045 10300
rect 23979 10235 24045 10236
rect 24347 10300 24413 10301
rect 24347 10236 24348 10300
rect 24412 10236 24413 10300
rect 24347 10235 24413 10236
rect 23427 5676 23493 5677
rect 23427 5612 23428 5676
rect 23492 5612 23493 5676
rect 23427 5611 23493 5612
rect 24534 5133 24594 20979
rect 24718 18730 24778 23971
rect 25451 23628 25517 23629
rect 25451 23564 25452 23628
rect 25516 23564 25517 23628
rect 25451 23563 25517 23564
rect 25267 23492 25333 23493
rect 25267 23428 25268 23492
rect 25332 23428 25333 23492
rect 25267 23427 25333 23428
rect 24718 18670 25146 18730
rect 24715 18052 24781 18053
rect 24715 17988 24716 18052
rect 24780 17988 24781 18052
rect 24715 17987 24781 17988
rect 24899 18052 24965 18053
rect 24899 17988 24900 18052
rect 24964 17988 24965 18052
rect 24899 17987 24965 17988
rect 24531 5132 24597 5133
rect 24531 5068 24532 5132
rect 24596 5068 24597 5132
rect 24531 5067 24597 5068
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 21955 3772 22021 3773
rect 21955 3708 21956 3772
rect 22020 3708 22021 3772
rect 21955 3707 22021 3708
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 21219 2412 21285 2413
rect 21219 2348 21220 2412
rect 21284 2348 21285 2412
rect 21219 2347 21285 2348
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 2128 23264 2688
rect 24718 2549 24778 17987
rect 24902 12613 24962 17987
rect 25086 15333 25146 18670
rect 25083 15332 25149 15333
rect 25083 15268 25084 15332
rect 25148 15268 25149 15332
rect 25083 15267 25149 15268
rect 25083 14924 25149 14925
rect 25083 14860 25084 14924
rect 25148 14860 25149 14924
rect 25083 14859 25149 14860
rect 24899 12612 24965 12613
rect 24899 12548 24900 12612
rect 24964 12548 24965 12612
rect 24899 12547 24965 12548
rect 25086 11661 25146 14859
rect 25083 11660 25149 11661
rect 25083 11596 25084 11660
rect 25148 11596 25149 11660
rect 25083 11595 25149 11596
rect 25270 7853 25330 23427
rect 25454 11253 25514 23563
rect 26003 23084 26069 23085
rect 26003 23020 26004 23084
rect 26068 23020 26069 23084
rect 26003 23019 26069 23020
rect 26006 22110 26066 23019
rect 26006 22050 26250 22110
rect 25635 19412 25701 19413
rect 25635 19348 25636 19412
rect 25700 19348 25701 19412
rect 25635 19347 25701 19348
rect 25451 11252 25517 11253
rect 25451 11188 25452 11252
rect 25516 11188 25517 11252
rect 25451 11187 25517 11188
rect 25638 10437 25698 19347
rect 26003 15196 26069 15197
rect 26003 15132 26004 15196
rect 26068 15132 26069 15196
rect 26003 15131 26069 15132
rect 25819 13836 25885 13837
rect 25819 13772 25820 13836
rect 25884 13772 25885 13836
rect 25819 13771 25885 13772
rect 25635 10436 25701 10437
rect 25635 10372 25636 10436
rect 25700 10372 25701 10436
rect 25635 10371 25701 10372
rect 25822 9210 25882 13771
rect 25638 9150 25882 9210
rect 25267 7852 25333 7853
rect 25267 7788 25268 7852
rect 25332 7788 25333 7852
rect 25267 7787 25333 7788
rect 25638 4181 25698 9150
rect 26006 8530 26066 15131
rect 25822 8470 26066 8530
rect 25822 6765 25882 8470
rect 26190 7850 26250 22050
rect 26006 7790 26250 7850
rect 26006 7445 26066 7790
rect 26003 7444 26069 7445
rect 26003 7380 26004 7444
rect 26068 7380 26069 7444
rect 26003 7379 26069 7380
rect 25819 6764 25885 6765
rect 25819 6700 25820 6764
rect 25884 6700 25885 6764
rect 25819 6699 25885 6700
rect 25635 4180 25701 4181
rect 25635 4116 25636 4180
rect 25700 4116 25701 4180
rect 25635 4115 25701 4116
rect 24715 2548 24781 2549
rect 24715 2484 24716 2548
rect 24780 2484 24781 2548
rect 24715 2483 24781 2484
use sky130_fd_sc_hd__clkbuf_2  _072_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21620 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1679235063
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp 1679235063
transform 1 0 16008 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp 1679235063
transform 1 0 20884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _076_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14720 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _077_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _078_
timestamp 1679235063
transform 1 0 18584 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1679235063
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp 1679235063
transform 1 0 23552 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1679235063
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1679235063
transform 1 0 23644 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1679235063
transform 1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _085_
timestamp 1679235063
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _086_
timestamp 1679235063
transform 1 0 10304 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _087_
timestamp 1679235063
transform 1 0 14260 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1679235063
transform 1 0 11776 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1679235063
transform 1 0 24932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1679235063
transform 1 0 11776 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1679235063
transform 1 0 19504 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _092_
timestamp 1679235063
transform 1 0 15548 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _093_
timestamp 1679235063
transform 1 0 10948 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _094_
timestamp 1679235063
transform 1 0 9384 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _095_
timestamp 1679235063
transform 1 0 12420 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _096_
timestamp 1679235063
transform 1 0 9108 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _097_
timestamp 1679235063
transform 1 0 12420 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _098_
timestamp 1679235063
transform 1 0 16836 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _099_
timestamp 1679235063
transform 1 0 14168 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_
timestamp 1679235063
transform 1 0 10304 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _101_
timestamp 1679235063
transform 1 0 11684 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1679235063
transform 1 0 11776 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1679235063
transform 1 0 16008 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _106_
timestamp 1679235063
transform 1 0 4692 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1679235063
transform 1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _108_
timestamp 1679235063
transform 1 0 5152 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_
timestamp 1679235063
transform 1 0 3220 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 15824 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1679235063
transform 1 0 18400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _114_
timestamp 1679235063
transform 1 0 6532 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _115_
timestamp 1679235063
transform 1 0 3404 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _116_
timestamp 1679235063
transform 1 0 3956 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _117_
timestamp 1679235063
transform 1 0 2576 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1679235063
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 9200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 6808 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _122_
timestamp 1679235063
transform 1 0 6348 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _123_
timestamp 1679235063
transform 1 0 1564 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _124_
timestamp 1679235063
transform 1 0 4048 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_
timestamp 1679235063
transform 1 0 1840 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1679235063
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1679235063
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1679235063
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1679235063
transform 1 0 7728 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1679235063
transform 1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 5612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 9752 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 17940 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1679235063
transform 1 0 17572 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1679235063
transform 1 0 19964 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1679235063
transform 1 0 20240 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1679235063
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1679235063
transform 1 0 20700 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1679235063
transform 1 0 17296 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1679235063
transform 1 0 18860 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1679235063
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1679235063
transform 1 0 16744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1679235063
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1679235063
transform 1 0 11592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1679235063
transform 1 0 20608 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1679235063
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1679235063
transform 1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1679235063
transform 1 0 22172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1679235063
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1679235063
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1679235063
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1679235063
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1679235063
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1679235063
transform 1 0 19320 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1679235063
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1679235063
transform 1 0 1472 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout125_A
timestamp 1679235063
transform 1 0 18032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout126_A
timestamp 1679235063
transform 1 0 13248 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout127_A
timestamp 1679235063
transform 1 0 19044 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout128_A
timestamp 1679235063
transform 1 0 21160 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout129_A
timestamp 1679235063
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold6_A
timestamp 1679235063
transform 1 0 1656 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold20_A
timestamp 1679235063
transform 1 0 20148 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold32_A
timestamp 1679235063
transform 1 0 25116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold49_A
timestamp 1679235063
transform 1 0 5152 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold66_A
timestamp 1679235063
transform 1 0 1656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold68_A
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold78_A
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold84_A
timestamp 1679235063
transform 1 0 22908 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold100_A
timestamp 1679235063
transform 1 0 1472 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold104_A
timestamp 1679235063
transform 1 0 16008 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold112_A
timestamp 1679235063
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold113_A
timestamp 1679235063
transform 1 0 1656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold132_A
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold133_A
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold136_A
timestamp 1679235063
transform 1 0 1656 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold152_A
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold160_A
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold162_A
timestamp 1679235063
transform 1 0 16100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold184_A
timestamp 1679235063
transform 1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold186_A
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold194_A
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold198_A
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold204_A
timestamp 1679235063
transform 1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold211_A
timestamp 1679235063
transform 1 0 5336 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold212_A
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold213_A
timestamp 1679235063
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold214_A
timestamp 1679235063
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1679235063
transform 1 0 19320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 1472 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 1656 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 4324 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 18124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 16652 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 12788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 2668 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 9016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 21896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 3220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 1472 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 2852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 5152 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 12328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 6716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 11592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 16468 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 6808 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 5152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1679235063
transform 1 0 23552 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1679235063
transform 1 0 6440 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1679235063
transform 1 0 6716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1679235063
transform 1 0 12696 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1679235063
transform 1 0 9108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 1656 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 1472 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 1656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20700 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21620 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 21896 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 20424 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20884 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20332 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17848 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16192 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13064 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21160 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 19320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 16284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21344 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 15272 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 3864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_14.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_14.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 24012 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21896 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22724 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 25300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 24012 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21344 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_32.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 22356 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17572 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18860 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14996 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 12604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 22724 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 1472 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 6440 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 9108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 17848 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 3864 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 25300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22540 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 2760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_12.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 2576 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 13616 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 5520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15272 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17204 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15180 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17020 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1679235063
transform 1 0 9476 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1679235063
transform 1 0 15640 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1679235063
transform 1 0 10396 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1679235063
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1679235063
transform 1 0 18216 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1679235063
transform 1 0 20792 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1679235063
transform 1 0 18216 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout124 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15824 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout125 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout126
timestamp 1679235063
transform 1 0 14260 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout127
timestamp 1679235063
transform 1 0 18400 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout128 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23092 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout129
timestamp 1679235063
transform 1 0 20608 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1679235063
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45
timestamp 1679235063
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1679235063
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95
timestamp 1679235063
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1679235063
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1679235063
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1679235063
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1679235063
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_165
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1679235063
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1679235063
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1679235063
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1679235063
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_263
timestamp 1679235063
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1679235063
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1679235063
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1679235063
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1679235063
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_65
timestamp 1679235063
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1679235063
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_88
timestamp 1679235063
transform 1 0 9200 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_100
timestamp 1679235063
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1679235063
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1679235063
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1679235063
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_161
timestamp 1679235063
transform 1 0 15916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_165
timestamp 1679235063
transform 1 0 16284 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1679235063
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1679235063
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1679235063
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1679235063
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1679235063
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1679235063
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 1679235063
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1679235063
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1679235063
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1679235063
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1679235063
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1679235063
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1679235063
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_168
timestamp 1679235063
transform 1 0 16560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1679235063
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1679235063
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1679235063
transform 1 0 18308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1679235063
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_200
timestamp 1679235063
transform 1 0 19504 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1679235063
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1679235063
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp 1679235063
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1679235063
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1679235063
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1679235063
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1679235063
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_70
timestamp 1679235063
transform 1 0 7544 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_82
timestamp 1679235063
transform 1 0 8648 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_94
timestamp 1679235063
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1679235063
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_161
timestamp 1679235063
transform 1 0 15916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1679235063
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_174
timestamp 1679235063
transform 1 0 17112 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1679235063
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1679235063
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1679235063
transform 1 0 19044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_202
timestamp 1679235063
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1679235063
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1679235063
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1679235063
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1679235063
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1679235063
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp 1679235063
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1679235063
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp 1679235063
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_158
timestamp 1679235063
transform 1 0 15640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_172
timestamp 1679235063
transform 1 0 16928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1679235063
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1679235063
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1679235063
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_199
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1679235063
transform 1 0 20424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1679235063
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_263
timestamp 1679235063
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_133
timestamp 1679235063
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_138
timestamp 1679235063
transform 1 0 13800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_142
timestamp 1679235063
transform 1 0 14168 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1679235063
transform 1 0 15180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_160
timestamp 1679235063
transform 1 0 15824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1679235063
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_174
timestamp 1679235063
transform 1 0 17112 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1679235063
transform 1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp 1679235063
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1679235063
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_210
timestamp 1679235063
transform 1 0 20424 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1679235063
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_127
timestamp 1679235063
transform 1 0 12788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1679235063
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1679235063
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_167
timestamp 1679235063
transform 1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_174
timestamp 1679235063
transform 1 0 17112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1679235063
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_199
timestamp 1679235063
transform 1 0 19412 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_216
timestamp 1679235063
transform 1 0 20976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1679235063
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1679235063
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_263
timestamp 1679235063
transform 1 0 25300 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1679235063
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1679235063
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_90
timestamp 1679235063
transform 1 0 9384 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1679235063
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1679235063
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1679235063
transform 1 0 11684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_124
timestamp 1679235063
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_131
timestamp 1679235063
transform 1 0 13156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_138
timestamp 1679235063
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_152
timestamp 1679235063
transform 1 0 15088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_159
timestamp 1679235063
transform 1 0 15732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1679235063
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_173
timestamp 1679235063
transform 1 0 17020 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1679235063
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_197
timestamp 1679235063
transform 1 0 19228 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_205
timestamp 1679235063
transform 1 0 19964 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_209
timestamp 1679235063
transform 1 0 20332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1679235063
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_235
timestamp 1679235063
transform 1 0 22724 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_239
timestamp 1679235063
transform 1 0 23092 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1679235063
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_246
timestamp 1679235063
transform 1 0 23736 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_112
timestamp 1679235063
transform 1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_119
timestamp 1679235063
transform 1 0 12052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_146
timestamp 1679235063
transform 1 0 14536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_151
timestamp 1679235063
transform 1 0 14996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1679235063
transform 1 0 15640 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_171
timestamp 1679235063
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_182
timestamp 1679235063
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1679235063
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_199
timestamp 1679235063
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1679235063
transform 1 0 20424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_222
timestamp 1679235063
transform 1 0 21528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_229
timestamp 1679235063
transform 1 0 22172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_233
timestamp 1679235063
transform 1 0 22540 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_263
timestamp 1679235063
transform 1 0 25300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1679235063
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_103
timestamp 1679235063
transform 1 0 10580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1679235063
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_119
timestamp 1679235063
transform 1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_133
timestamp 1679235063
transform 1 0 13340 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_147
timestamp 1679235063
transform 1 0 14628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1679235063
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1679235063
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1679235063
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1679235063
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1679235063
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1679235063
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1679235063
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1679235063
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_14
timestamp 1679235063
transform 1 0 2392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_18
timestamp 1679235063
transform 1 0 2760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_21
timestamp 1679235063
transform 1 0 3036 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_25
timestamp 1679235063
transform 1 0 3404 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1679235063
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1679235063
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1679235063
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_117
timestamp 1679235063
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1679235063
transform 1 0 12604 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 1679235063
transform 1 0 12972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1679235063
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_143
timestamp 1679235063
transform 1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_165
timestamp 1679235063
transform 1 0 16284 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1679235063
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1679235063
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1679235063
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_207
timestamp 1679235063
transform 1 0 20148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_211
timestamp 1679235063
transform 1 0 20516 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1679235063
transform 1 0 21160 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1679235063
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_263
timestamp 1679235063
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_12
timestamp 1679235063
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_19
timestamp 1679235063
transform 1 0 2852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_26
timestamp 1679235063
transform 1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1679235063
transform 1 0 3864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1679235063
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_40
timestamp 1679235063
transform 1 0 4784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1679235063
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1679235063
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_64
timestamp 1679235063
transform 1 0 6992 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_76
timestamp 1679235063
transform 1 0 8096 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp 1679235063
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_91
timestamp 1679235063
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_96
timestamp 1679235063
transform 1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1679235063
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_133
timestamp 1679235063
transform 1 0 13340 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1679235063
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_154
timestamp 1679235063
transform 1 0 15272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1679235063
transform 1 0 17572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1679235063
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_203
timestamp 1679235063
transform 1 0 19780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1679235063
transform 1 0 20884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1679235063
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1679235063
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1679235063
transform 1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_12
timestamp 1679235063
transform 1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_19
timestamp 1679235063
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1679235063
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1679235063
transform 1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1679235063
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_42
timestamp 1679235063
transform 1 0 4968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_46
timestamp 1679235063
transform 1 0 5336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_50
timestamp 1679235063
transform 1 0 5704 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_54
timestamp 1679235063
transform 1 0 6072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_58
timestamp 1679235063
transform 1 0 6440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1679235063
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_66
timestamp 1679235063
transform 1 0 7176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_70
timestamp 1679235063
transform 1 0 7544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_74
timestamp 1679235063
transform 1 0 7912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1679235063
transform 1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1679235063
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1679235063
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_92
timestamp 1679235063
transform 1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_96
timestamp 1679235063
transform 1 0 9936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1679235063
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_124
timestamp 1679235063
transform 1 0 12512 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1679235063
transform 1 0 14628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_151
timestamp 1679235063
transform 1 0 14996 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_160
timestamp 1679235063
transform 1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_172
timestamp 1679235063
transform 1 0 16928 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_184
timestamp 1679235063
transform 1 0 18032 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_207
timestamp 1679235063
transform 1 0 20148 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1679235063
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_227
timestamp 1679235063
transform 1 0 21988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_231
timestamp 1679235063
transform 1 0 22356 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_263
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1679235063
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_14
timestamp 1679235063
transform 1 0 2392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1679235063
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1679235063
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_35
timestamp 1679235063
transform 1 0 4324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1679235063
transform 1 0 4968 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1679235063
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1679235063
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_63
timestamp 1679235063
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_67
timestamp 1679235063
transform 1 0 7268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_71
timestamp 1679235063
transform 1 0 7636 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1679235063
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1679235063
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1679235063
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1679235063
transform 1 0 11960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_130
timestamp 1679235063
transform 1 0 13064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1679235063
transform 1 0 14168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_154
timestamp 1679235063
transform 1 0 15272 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1679235063
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1679235063
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1679235063
transform 1 0 18860 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_197
timestamp 1679235063
transform 1 0 19228 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1679235063
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_219
timestamp 1679235063
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1679235063
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1679235063
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1679235063
transform 1 0 2392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1679235063
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1679235063
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_50
timestamp 1679235063
transform 1 0 5704 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_55
timestamp 1679235063
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_63
timestamp 1679235063
transform 1 0 6900 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_74
timestamp 1679235063
transform 1 0 7912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1679235063
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1679235063
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_100
timestamp 1679235063
transform 1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1679235063
transform 1 0 11408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1679235063
transform 1 0 11776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_126
timestamp 1679235063
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_143
timestamp 1679235063
transform 1 0 14260 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 1679235063
transform 1 0 14628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_156
timestamp 1679235063
transform 1 0 15456 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_168
timestamp 1679235063
transform 1 0 16560 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1679235063
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_192
timestamp 1679235063
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_200
timestamp 1679235063
transform 1 0 19504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_210
timestamp 1679235063
transform 1 0 20424 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1679235063
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_240
timestamp 1679235063
transform 1 0 23184 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_248
timestamp 1679235063
transform 1 0 23920 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_264
timestamp 1679235063
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_21
timestamp 1679235063
transform 1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_25
timestamp 1679235063
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1679235063
transform 1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_46
timestamp 1679235063
transform 1 0 5336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1679235063
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_63
timestamp 1679235063
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1679235063
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 1679235063
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_82
timestamp 1679235063
transform 1 0 8648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_89
timestamp 1679235063
transform 1 0 9292 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1679235063
transform 1 0 9936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1679235063
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_124
timestamp 1679235063
transform 1 0 12512 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_136
timestamp 1679235063
transform 1 0 13616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1679235063
transform 1 0 14720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 1679235063
transform 1 0 15824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1679235063
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1679235063
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_183
timestamp 1679235063
transform 1 0 17940 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1679235063
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_204
timestamp 1679235063
transform 1 0 19872 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_216
timestamp 1679235063
transform 1 0 20976 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1679235063
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1679235063
transform 1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_20
timestamp 1679235063
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1679235063
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_31
timestamp 1679235063
transform 1 0 3956 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_47
timestamp 1679235063
transform 1 0 5428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_51
timestamp 1679235063
transform 1 0 5796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1679235063
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1679235063
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1679235063
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_103
timestamp 1679235063
transform 1 0 10580 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_108
timestamp 1679235063
transform 1 0 11040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1679235063
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1679235063
transform 1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1679235063
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1679235063
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1679235063
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1679235063
transform 1 0 17480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_190
timestamp 1679235063
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1679235063
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1679235063
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_227
timestamp 1679235063
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_231
timestamp 1679235063
transform 1 0 22356 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1679235063
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1679235063
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_6
timestamp 1679235063
transform 1 0 1656 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1679235063
transform 1 0 2116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_18
timestamp 1679235063
transform 1 0 2760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_25
timestamp 1679235063
transform 1 0 3404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1679235063
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1679235063
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_73
timestamp 1679235063
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1679235063
transform 1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1679235063
transform 1 0 9016 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1679235063
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1679235063
transform 1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1679235063
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1679235063
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1679235063
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_154
timestamp 1679235063
transform 1 0 15272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1679235063
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_197
timestamp 1679235063
transform 1 0 19228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_218
timestamp 1679235063
transform 1 0 21160 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1679235063
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1679235063
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1679235063
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1679235063
transform 1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_19
timestamp 1679235063
transform 1 0 2852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1679235063
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_35
timestamp 1679235063
transform 1 0 4324 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_49
timestamp 1679235063
transform 1 0 5612 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp 1679235063
transform 1 0 6256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1679235063
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1679235063
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_90
timestamp 1679235063
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1679235063
transform 1 0 10488 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_114
timestamp 1679235063
transform 1 0 11592 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1679235063
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_151
timestamp 1679235063
transform 1 0 14996 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_156
timestamp 1679235063
transform 1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1679235063
transform 1 0 17480 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1679235063
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_219
timestamp 1679235063
transform 1 0 21252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_225
timestamp 1679235063
transform 1 0 21804 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_247
timestamp 1679235063
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_263
timestamp 1679235063
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1679235063
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1679235063
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_19
timestamp 1679235063
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_33
timestamp 1679235063
transform 1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_46
timestamp 1679235063
transform 1 0 5336 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_50
timestamp 1679235063
transform 1 0 5704 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1679235063
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1679235063
transform 1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_76
timestamp 1679235063
transform 1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_83
timestamp 1679235063
transform 1 0 8740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_88
timestamp 1679235063
transform 1 0 9200 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1679235063
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1679235063
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_128
timestamp 1679235063
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1679235063
transform 1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1679235063
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_191
timestamp 1679235063
transform 1 0 18676 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1679235063
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1679235063
transform 1 0 21068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_228
timestamp 1679235063
transform 1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1679235063
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_263
timestamp 1679235063
transform 1 0 25300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_14
timestamp 1679235063
transform 1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1679235063
transform 1 0 3036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1679235063
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1679235063
transform 1 0 5520 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1679235063
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1679235063
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1679235063
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_89
timestamp 1679235063
transform 1 0 9292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_111
timestamp 1679235063
transform 1 0 11316 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1679235063
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1679235063
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_152
timestamp 1679235063
transform 1 0 15088 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_156
timestamp 1679235063
transform 1 0 15456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1679235063
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_182
timestamp 1679235063
transform 1 0 17848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_192
timestamp 1679235063
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_200
timestamp 1679235063
transform 1 0 19504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1679235063
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_246
timestamp 1679235063
transform 1 0 23736 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_263
timestamp 1679235063
transform 1 0 25300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1679235063
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp 1679235063
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_35
timestamp 1679235063
transform 1 0 4324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_42
timestamp 1679235063
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1679235063
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1679235063
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_74
timestamp 1679235063
transform 1 0 7912 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1679235063
transform 1 0 9016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_120
timestamp 1679235063
transform 1 0 12144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1679235063
transform 1 0 13248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_156
timestamp 1679235063
transform 1 0 15456 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_179
timestamp 1679235063
transform 1 0 17572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1679235063
transform 1 0 18032 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_206
timestamp 1679235063
transform 1 0 20056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_228
timestamp 1679235063
transform 1 0 22080 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_250
timestamp 1679235063
transform 1 0 24104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_262
timestamp 1679235063
transform 1 0 25208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1679235063
transform 1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1679235063
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1679235063
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1679235063
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1679235063
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_70
timestamp 1679235063
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_89
timestamp 1679235063
transform 1 0 9292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1679235063
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_123
timestamp 1679235063
transform 1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_127
timestamp 1679235063
transform 1 0 12788 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1679235063
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1679235063
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1679235063
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1679235063
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1679235063
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_247
timestamp 1679235063
transform 1 0 23828 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1679235063
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_264
timestamp 1679235063
transform 1 0 25392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1679235063
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1679235063
transform 1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1679235063
transform 1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1679235063
transform 1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1679235063
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1679235063
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_74
timestamp 1679235063
transform 1 0 7912 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_86
timestamp 1679235063
transform 1 0 9016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_98
timestamp 1679235063
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_121
timestamp 1679235063
transform 1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_125
timestamp 1679235063
transform 1 0 12604 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_146
timestamp 1679235063
transform 1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_158
timestamp 1679235063
transform 1 0 15640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_191
timestamp 1679235063
transform 1 0 18676 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1679235063
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1679235063
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1679235063
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1679235063
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_6
timestamp 1679235063
transform 1 0 1656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1679235063
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1679235063
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1679235063
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_46
timestamp 1679235063
transform 1 0 5336 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_58
timestamp 1679235063
transform 1 0 6440 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1679235063
transform 1 0 7544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_96
timestamp 1679235063
transform 1 0 9936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_120
timestamp 1679235063
transform 1 0 12144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_133
timestamp 1679235063
transform 1 0 13340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1679235063
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_167
timestamp 1679235063
transform 1 0 16468 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1679235063
transform 1 0 16744 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1679235063
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1679235063
transform 1 0 20424 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1679235063
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_235
timestamp 1679235063
transform 1 0 22724 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_247
timestamp 1679235063
transform 1 0 23828 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1679235063
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_263
timestamp 1679235063
transform 1 0 25300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1679235063
transform 1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_18
timestamp 1679235063
transform 1 0 2760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1679235063
transform 1 0 3864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_42
timestamp 1679235063
transform 1 0 4968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1679235063
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_74
timestamp 1679235063
transform 1 0 7912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1679235063
transform 1 0 9016 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1679235063
transform 1 0 10120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1679235063
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_148
timestamp 1679235063
transform 1 0 14720 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_153
timestamp 1679235063
transform 1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1679235063
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_193
timestamp 1679235063
transform 1 0 18860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1679235063
transform 1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_219
timestamp 1679235063
transform 1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1679235063
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1679235063
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1679235063
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1679235063
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_263
timestamp 1679235063
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_14
timestamp 1679235063
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1679235063
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_39
timestamp 1679235063
transform 1 0 4692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_46
timestamp 1679235063
transform 1 0 5336 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_58
timestamp 1679235063
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_70
timestamp 1679235063
transform 1 0 7544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_91
timestamp 1679235063
transform 1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1679235063
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1679235063
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1679235063
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1679235063
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1679235063
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1679235063
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1679235063
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1679235063
transform 1 0 1840 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_18
timestamp 1679235063
transform 1 0 2760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_30
timestamp 1679235063
transform 1 0 3864 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_42
timestamp 1679235063
transform 1 0 4968 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_59
timestamp 1679235063
transform 1 0 6532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1679235063
transform 1 0 6808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_72
timestamp 1679235063
transform 1 0 7728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1679235063
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1679235063
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_120
timestamp 1679235063
transform 1 0 12144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1679235063
transform 1 0 14352 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_151
timestamp 1679235063
transform 1 0 14996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_164
timestamp 1679235063
transform 1 0 16192 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_180
timestamp 1679235063
transform 1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_186
timestamp 1679235063
transform 1 0 18216 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_208
timestamp 1679235063
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_220
timestamp 1679235063
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_230
timestamp 1679235063
transform 1 0 22264 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_252
timestamp 1679235063
transform 1 0 24288 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1679235063
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_14
timestamp 1679235063
transform 1 0 2392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1679235063
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_34
timestamp 1679235063
transform 1 0 4232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_46
timestamp 1679235063
transform 1 0 5336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1679235063
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_70
timestamp 1679235063
transform 1 0 7544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_89
timestamp 1679235063
transform 1 0 9292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_111
timestamp 1679235063
transform 1 0 11316 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_135
timestamp 1679235063
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1679235063
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1679235063
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1679235063
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_190
timestamp 1679235063
transform 1 0 18584 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1679235063
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1679235063
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1679235063
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_233
timestamp 1679235063
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_239
timestamp 1679235063
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_263
timestamp 1679235063
transform 1 0 25300 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1679235063
transform 1 0 1840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_18
timestamp 1679235063
transform 1 0 2760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_30
timestamp 1679235063
transform 1 0 3864 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_42
timestamp 1679235063
transform 1 0 4968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1679235063
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1679235063
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp 1679235063
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1679235063
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_155
timestamp 1679235063
transform 1 0 15364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_171
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_182
timestamp 1679235063
transform 1 0 17848 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1679235063
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_219
timestamp 1679235063
transform 1 0 21252 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1679235063
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1679235063
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_259
timestamp 1679235063
transform 1 0 24932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_265
timestamp 1679235063
transform 1 0 25484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_14
timestamp 1679235063
transform 1 0 2392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1679235063
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 1679235063
transform 1 0 4232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_46
timestamp 1679235063
transform 1 0 5336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1679235063
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_70
timestamp 1679235063
transform 1 0 7544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1679235063
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1679235063
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1679235063
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1679235063
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_156
timestamp 1679235063
transform 1 0 15456 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_177
timestamp 1679235063
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_181
timestamp 1679235063
transform 1 0 17756 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1679235063
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_204
timestamp 1679235063
transform 1 0 19872 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_228
timestamp 1679235063
transform 1 0 22080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_241
timestamp 1679235063
transform 1 0 23276 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1679235063
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1679235063
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_23
timestamp 1679235063
transform 1 0 3220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_30
timestamp 1679235063
transform 1 0 3864 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_42
timestamp 1679235063
transform 1 0 4968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_69
timestamp 1679235063
transform 1 0 7452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_81
timestamp 1679235063
transform 1 0 8556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_105
timestamp 1679235063
transform 1 0 10764 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_120
timestamp 1679235063
transform 1 0 12144 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_144
timestamp 1679235063
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1679235063
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_161
timestamp 1679235063
transform 1 0 15916 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1679235063
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1679235063
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_219
timestamp 1679235063
transform 1 0 21252 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1679235063
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1679235063
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1679235063
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_262
timestamp 1679235063
transform 1 0 25208 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_8
timestamp 1679235063
transform 1 0 1840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1679235063
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_34
timestamp 1679235063
transform 1 0 4232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_46
timestamp 1679235063
transform 1 0 5336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_58
timestamp 1679235063
transform 1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1679235063
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_96
timestamp 1679235063
transform 1 0 9936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1679235063
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_133
timestamp 1679235063
transform 1 0 13340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1679235063
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1679235063
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_172
timestamp 1679235063
transform 1 0 16928 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_190
timestamp 1679235063
transform 1 0 18584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_212
timestamp 1679235063
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_235
timestamp 1679235063
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_248
timestamp 1679235063
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1679235063
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_5
timestamp 1679235063
transform 1 0 1564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_35
timestamp 1679235063
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_42
timestamp 1679235063
transform 1 0 4968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1679235063
transform 1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1679235063
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_81
timestamp 1679235063
transform 1 0 8556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_105
timestamp 1679235063
transform 1 0 10764 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_109
timestamp 1679235063
transform 1 0 11132 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1679235063
transform 1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_128
timestamp 1679235063
transform 1 0 12880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_134
timestamp 1679235063
transform 1 0 13432 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_156
timestamp 1679235063
transform 1 0 15456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_164
timestamp 1679235063
transform 1 0 16192 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_171
timestamp 1679235063
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_194
timestamp 1679235063
transform 1 0 18952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_208
timestamp 1679235063
transform 1 0 20240 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1679235063
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1679235063
transform 1 0 22816 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_240
timestamp 1679235063
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_263
timestamp 1679235063
transform 1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_8
timestamp 1679235063
transform 1 0 1840 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1679235063
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_59
timestamp 1679235063
transform 1 0 6532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_79
timestamp 1679235063
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_92
timestamp 1679235063
transform 1 0 9568 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1679235063
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1679235063
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1679235063
transform 1 0 13340 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1679235063
transform 1 0 14812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_153
timestamp 1679235063
transform 1 0 15180 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1679235063
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1679235063
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1679235063
transform 1 0 18492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_193
timestamp 1679235063
transform 1 0 18860 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_219
timestamp 1679235063
transform 1 0 21252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_225
timestamp 1679235063
transform 1 0 21804 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1679235063
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1679235063
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1679235063
transform 1 0 2392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1679235063
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_63
timestamp 1679235063
transform 1 0 6900 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_81
timestamp 1679235063
transform 1 0 8556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_105
timestamp 1679235063
transform 1 0 10764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_109
timestamp 1679235063
transform 1 0 11132 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_119
timestamp 1679235063
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_130
timestamp 1679235063
transform 1 0 13064 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_154
timestamp 1679235063
transform 1 0 15272 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_180
timestamp 1679235063
transform 1 0 17664 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_184
timestamp 1679235063
transform 1 0 18032 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_207
timestamp 1679235063
transform 1 0 20148 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_211
timestamp 1679235063
transform 1 0 20516 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1679235063
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_8
timestamp 1679235063
transform 1 0 1840 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1679235063
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1679235063
transform 1 0 4048 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_42
timestamp 1679235063
transform 1 0 4968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1679235063
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_89
timestamp 1679235063
transform 1 0 9292 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1679235063
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1679235063
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_132
timestamp 1679235063
transform 1 0 13248 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_152
timestamp 1679235063
transform 1 0 15088 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_156
timestamp 1679235063
transform 1 0 15456 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1679235063
transform 1 0 17572 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_192
timestamp 1679235063
transform 1 0 18768 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1679235063
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1679235063
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_229
timestamp 1679235063
transform 1 0 22172 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_237
timestamp 1679235063
transform 1 0 22908 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1679235063
transform 1 0 2392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_60
timestamp 1679235063
transform 1 0 6624 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_66
timestamp 1679235063
transform 1 0 7176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1679235063
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_125
timestamp 1679235063
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1679235063
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1679235063
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1679235063
transform 1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_180
timestamp 1679235063
transform 1 0 17664 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1679235063
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1679235063
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_219
timestamp 1679235063
transform 1 0 21252 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1679235063
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_235
timestamp 1679235063
transform 1 0 22724 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_259
timestamp 1679235063
transform 1 0 24932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_265
timestamp 1679235063
transform 1 0 25484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_8
timestamp 1679235063
transform 1 0 1840 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1679235063
transform 1 0 4048 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1679235063
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_89
timestamp 1679235063
transform 1 0 9292 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_99
timestamp 1679235063
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_123
timestamp 1679235063
transform 1 0 12420 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_128
timestamp 1679235063
transform 1 0 12880 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1679235063
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1679235063
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_184
timestamp 1679235063
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_192
timestamp 1679235063
transform 1 0 18768 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1679235063
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1679235063
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_60
timestamp 1679235063
transform 1 0 6624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1679235063
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_117
timestamp 1679235063
transform 1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_135
timestamp 1679235063
transform 1 0 13524 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_139
timestamp 1679235063
transform 1 0 13892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_150
timestamp 1679235063
transform 1 0 14904 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_162
timestamp 1679235063
transform 1 0 16008 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1679235063
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1679235063
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_218
timestamp 1679235063
transform 1 0 21160 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1679235063
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1679235063
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_263
timestamp 1679235063
transform 1 0 25300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1679235063
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_159
timestamp 1679235063
transform 1 0 15732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_181
timestamp 1679235063
transform 1 0 17756 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_203
timestamp 1679235063
transform 1 0 19780 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_216
timestamp 1679235063
transform 1 0 20976 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1679235063
transform 1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 4232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 20332 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold5 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17388 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 3128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 4232 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold9
timestamp 1679235063
transform 1 0 20608 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold10
timestamp 1679235063
transform 1 0 24564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 23092 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold15
timestamp 1679235063
transform 1 0 6808 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold16
timestamp 1679235063
transform 1 0 19688 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 13984 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform 1 0 17940 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold20
timestamp 1679235063
transform 1 0 20516 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold21
timestamp 1679235063
transform 1 0 1656 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform 1 0 5704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold23
timestamp 1679235063
transform 1 0 5060 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 12512 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 4600 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold27
timestamp 1679235063
transform 1 0 6808 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 13892 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 4232 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold32
timestamp 1679235063
transform 1 0 24656 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 15088 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 1656 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold36
timestamp 1679235063
transform 1 0 16652 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 17848 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold38
timestamp 1679235063
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold39
timestamp 1679235063
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 9200 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold41
timestamp 1679235063
transform 1 0 17112 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 17296 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 15272 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 11684 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold45
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold46
timestamp 1679235063
transform 1 0 5704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 7820 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold48
timestamp 1679235063
transform 1 0 11408 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold49
timestamp 1679235063
transform 1 0 5704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold51
timestamp 1679235063
transform 1 0 6808 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 3956 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 8280 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 16928 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 18584 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 6808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold58
timestamp 1679235063
transform 1 0 1656 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 6992 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 19688 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 19412 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform 1 0 6808 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 24564 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 21528 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold65
timestamp 1679235063
transform 1 0 19596 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold66
timestamp 1679235063
transform 1 0 3128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 8280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold68
timestamp 1679235063
transform 1 0 9476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold69
timestamp 1679235063
transform 1 0 5704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform 1 0 6716 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1679235063
transform 1 0 2024 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold72
timestamp 1679235063
transform 1 0 7176 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold73
timestamp 1679235063
transform 1 0 11960 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1679235063
transform 1 0 6440 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1679235063
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold77
timestamp 1679235063
transform 1 0 9844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold78
timestamp 1679235063
transform 1 0 10672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold79
timestamp 1679235063
transform 1 0 2576 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold80
timestamp 1679235063
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold81
timestamp 1679235063
transform 1 0 19688 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold82
timestamp 1679235063
transform 1 0 9384 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 12144 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 19688 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform 1 0 12328 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold86
timestamp 1679235063
transform 1 0 1748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold87
timestamp 1679235063
transform 1 0 2024 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold88
timestamp 1679235063
transform 1 0 20240 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold89
timestamp 1679235063
transform 1 0 20516 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold90
timestamp 1679235063
transform 1 0 14904 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold91
timestamp 1679235063
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold92
timestamp 1679235063
transform 1 0 21344 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold93
timestamp 1679235063
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold95
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold96
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1679235063
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold99
timestamp 1679235063
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold100
timestamp 1679235063
transform 1 0 2024 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold101
timestamp 1679235063
transform 1 0 14536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold102
timestamp 1679235063
transform 1 0 19780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold103
timestamp 1679235063
transform 1 0 24472 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold104
timestamp 1679235063
transform 1 0 14720 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold105
timestamp 1679235063
transform 1 0 24564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold106
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold107
timestamp 1679235063
transform 1 0 24564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold108
timestamp 1679235063
transform 1 0 15824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold109
timestamp 1679235063
transform 1 0 16192 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold110
timestamp 1679235063
transform 1 0 17756 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold111
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold112
timestamp 1679235063
transform 1 0 7176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold113
timestamp 1679235063
transform 1 0 1656 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold114
timestamp 1679235063
transform 1 0 3128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold115
timestamp 1679235063
transform 1 0 7176 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold116
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold117
timestamp 1679235063
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold118
timestamp 1679235063
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold119
timestamp 1679235063
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold120
timestamp 1679235063
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold121
timestamp 1679235063
transform 1 0 4232 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold122
timestamp 1679235063
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold123
timestamp 1679235063
transform 1 0 12880 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold124
timestamp 1679235063
transform 1 0 4600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold125
timestamp 1679235063
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold126
timestamp 1679235063
transform 1 0 16836 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold127
timestamp 1679235063
transform 1 0 19688 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold128
timestamp 1679235063
transform 1 0 6716 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold129
timestamp 1679235063
transform 1 0 5704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold130
timestamp 1679235063
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold131
timestamp 1679235063
transform 1 0 4600 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold132
timestamp 1679235063
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold133
timestamp 1679235063
transform 1 0 19228 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold134
timestamp 1679235063
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold135
timestamp 1679235063
transform 1 0 13432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold136
timestamp 1679235063
transform 1 0 4232 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold137
timestamp 1679235063
transform 1 0 20516 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold138
timestamp 1679235063
transform 1 0 1656 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold139
timestamp 1679235063
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold140
timestamp 1679235063
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold141
timestamp 1679235063
transform 1 0 14352 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold142
timestamp 1679235063
transform 1 0 21988 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold143
timestamp 1679235063
transform 1 0 18032 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold144
timestamp 1679235063
transform 1 0 10856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold145
timestamp 1679235063
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold146
timestamp 1679235063
transform 1 0 14536 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold147
timestamp 1679235063
transform 1 0 17848 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold148
timestamp 1679235063
transform 1 0 17020 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold149
timestamp 1679235063
transform 1 0 18124 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold150
timestamp 1679235063
transform 1 0 11776 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold151
timestamp 1679235063
transform 1 0 18124 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold152
timestamp 1679235063
transform 1 0 3128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18216 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold154
timestamp 1679235063
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold155
timestamp 1679235063
transform 1 0 10304 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold156
timestamp 1679235063
transform 1 0 7820 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold157
timestamp 1679235063
transform 1 0 13064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold158
timestamp 1679235063
transform 1 0 7176 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold159
timestamp 1679235063
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold160
timestamp 1679235063
transform 1 0 7912 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold161
timestamp 1679235063
transform 1 0 9200 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold162
timestamp 1679235063
transform 1 0 14444 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold163
timestamp 1679235063
transform 1 0 10304 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold164
timestamp 1679235063
transform 1 0 14536 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold165
timestamp 1679235063
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold166
timestamp 1679235063
transform 1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  hold167
timestamp 1679235063
transform 1 0 15640 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold168
timestamp 1679235063
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold169
timestamp 1679235063
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold170
timestamp 1679235063
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold171
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold172
timestamp 1679235063
transform 1 0 5796 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold173
timestamp 1679235063
transform 1 0 6716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold174
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold175
timestamp 1679235063
transform 1 0 18032 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold176
timestamp 1679235063
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold177
timestamp 1679235063
transform 1 0 8280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold178
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold179
timestamp 1679235063
transform 1 0 21988 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold180
timestamp 1679235063
transform 1 0 6808 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold181
timestamp 1679235063
transform 1 0 9384 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold182
timestamp 1679235063
transform 1 0 9476 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold183
timestamp 1679235063
transform 1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold184
timestamp 1679235063
transform 1 0 1656 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold185
timestamp 1679235063
transform 1 0 1656 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold186
timestamp 1679235063
transform 1 0 13432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold187
timestamp 1679235063
transform 1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold188
timestamp 1679235063
transform 1 0 19044 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold189
timestamp 1679235063
transform 1 0 20148 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold190
timestamp 1679235063
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold191
timestamp 1679235063
transform 1 0 18492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold192
timestamp 1679235063
transform 1 0 6808 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold193
timestamp 1679235063
transform 1 0 6808 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold194
timestamp 1679235063
transform 1 0 4600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold195
timestamp 1679235063
transform 1 0 5704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold196
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold197
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold198
timestamp 1679235063
transform 1 0 15088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold199
timestamp 1679235063
transform 1 0 9752 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold200
timestamp 1679235063
transform 1 0 4600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold201
timestamp 1679235063
transform 1 0 5704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold202
timestamp 1679235063
transform 1 0 21988 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold203
timestamp 1679235063
transform 1 0 20792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold204
timestamp 1679235063
transform 1 0 15548 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1679235063
transform 1 0 11960 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold206
timestamp 1679235063
transform 1 0 9384 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold207
timestamp 1679235063
transform 1 0 4232 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold208
timestamp 1679235063
transform 1 0 9476 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold209
timestamp 1679235063
transform 1 0 7820 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold210
timestamp 1679235063
transform 1 0 24196 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold211
timestamp 1679235063
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold212
timestamp 1679235063
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold213
timestamp 1679235063
transform 1 0 12512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold214
timestamp 1679235063
transform 1 0 9108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold215
timestamp 1679235063
transform 1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold216
timestamp 1679235063
transform 1 0 7360 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold217
timestamp 1679235063
transform 1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold218
timestamp 1679235063
transform 1 0 7544 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 6716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 6532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1679235063
transform 1 0 3956 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 6532 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 4692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 9660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1679235063
transform 1 0 14720 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1679235063
transform 1 0 15364 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1679235063
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1679235063
transform 1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1679235063
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1679235063
transform 1 0 9016 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1679235063
transform 1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 4692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 12972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1679235063
transform 1 0 2116 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1679235063
transform 1 0 13524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 16100 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1679235063
transform 1 0 4416 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1679235063
transform 1 0 3772 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1679235063
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1679235063
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1679235063
transform 1 0 4048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 8464 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1679235063
transform 1 0 4508 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1679235063
transform 1 0 11684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1679235063
transform 1 0 3956 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1679235063
transform 1 0 6624 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1679235063
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1679235063
transform 1 0 7084 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1679235063
transform 1 0 9016 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1679235063
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1679235063
transform 1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1679235063
transform 1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 8372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1679235063
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input62 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  output63 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1679235063
transform 1 0 20056 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1679235063
transform 1 0 22080 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1679235063
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1679235063
transform 1 0 22632 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1679235063
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1679235063
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1679235063
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1679235063
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1679235063
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1679235063
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1679235063
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1679235063
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1679235063
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1679235063
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1679235063
transform 1 0 22080 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1679235063
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 22080 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 20792 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 1748 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 5336 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 7084 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 7176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 7544 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 10580 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 12052 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 2852 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 2760 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 2760 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 2024 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 4600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14904 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17020 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20332 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21620 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22632 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22172 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23092 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23276 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23460 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23276 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22448 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20884 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20240 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20700 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22724 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22356 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21896 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19320 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18400 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15640 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15640 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17020 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19320 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21252 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15548 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18308 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18032 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15732 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14996 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13616 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13432 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13616 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12512 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11500 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11132 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10580 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8924 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8924 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8924 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8924 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9200 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9476 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12512 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10304 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10580 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9384 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12696 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13248 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13616 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17664 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_0.mux_l1_in_1__157 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_2.mux_l2_in_0__163
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23092 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_4.mux_l2_in_0__132
timestamp 1679235063
transform 1 0 2760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_6.mux_l1_in_1__137
timestamp 1679235063
transform 1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_8.mux_l2_in_0__138
timestamp 1679235063
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_10.mux_l2_in_0__158
timestamp 1679235063
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_12.mux_l2_in_0__159
timestamp 1679235063
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_14.mux_l2_in_0__160
timestamp 1679235063
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22080 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_16.mux_l2_in_0__161
timestamp 1679235063
transform 1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22448 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23000 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_18.mux_l2_in_0__162
timestamp 1679235063
transform 1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_28.mux_l2_in_0__164
timestamp 1679235063
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20792 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_30.mux_l2_in_0__165
timestamp 1679235063
transform 1 0 11776 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20608 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19596 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_32.mux_l2_in_0__130
timestamp 1679235063
transform 1 0 5060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_34.mux_l2_in_0__131
timestamp 1679235063
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17940 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_44.mux_l2_in_0__133
timestamp 1679235063
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_46.mux_l2_in_0__134
timestamp 1679235063
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_48.mux_l2_in_0__135
timestamp 1679235063
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_50.mux_l2_in_0__136
timestamp 1679235063
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_0.mux_l1_in_1__139
timestamp 1679235063
transform 1 0 17296 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_2.mux_l2_in_0__145
timestamp 1679235063
transform 1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20332 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_4.mux_l2_in_0__150
timestamp 1679235063
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20148 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_6.mux_l1_in_1__155
timestamp 1679235063
transform 1 0 2576 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17204 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14076 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_8.mux_l2_in_0__156
timestamp 1679235063
transform 1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17940 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_10.mux_l2_in_0__140
timestamp 1679235063
transform 1 0 18308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16468 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_12.mux_l2_in_0__141
timestamp 1679235063
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12420 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_14.mux_l2_in_0__142
timestamp 1679235063
transform 1 0 3220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15272 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9936 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_16.mux_l2_in_0__143
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16100 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_18.mux_l2_in_0__144
timestamp 1679235063
transform 1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14720 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10304 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_28.mux_l2_in_0__146
timestamp 1679235063
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17756 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_30.mux_l2_in_0__147
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_32.mux_l2_in_0__148
timestamp 1679235063
transform 1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15364 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_34.mux_l2_in_0__149
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15364 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_44.mux_l2_in_0__151
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10764 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2576 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12512 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_46.mux_l2_in_0__152
timestamp 1679235063
transform 1 0 6532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_48.mux_l2_in_0__153
timestamp 1679235063
transform 1 0 14996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17112 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_50.mux_l2_in_0__154
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 26200 280 27000 400 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 26200 17416 27000 17536 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 26200 18232 27000 18352 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 26200 19048 27000 19168 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 26200 20680 27000 20800 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 26200 13336 27000 13456 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 16 nsew signal input
flabel metal3 s 26200 21496 27000 21616 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 17 nsew signal input
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 18 nsew signal input
flabel metal3 s 26200 22312 27000 22432 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 19 nsew signal input
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 20 nsew signal input
flabel metal3 s 26200 23128 27000 23248 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 21 nsew signal input
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 22 nsew signal input
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 23 nsew signal input
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 24 nsew signal input
flabel metal3 s 26200 24760 27000 24880 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 25 nsew signal input
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 26 nsew signal input
flabel metal3 s 26200 14152 27000 14272 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 27 nsew signal input
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 28 nsew signal input
flabel metal3 s 26200 14968 27000 15088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 29 nsew signal input
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 30 nsew signal input
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 31 nsew signal input
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 32 nsew signal input
flabel metal3 s 26200 16600 27000 16720 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 33 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 34 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 35 nsew signal tristate
flabel metal3 s 26200 5176 27000 5296 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 36 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 37 nsew signal tristate
flabel metal3 s 26200 5992 27000 6112 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 38 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 39 nsew signal tristate
flabel metal3 s 26200 6808 27000 6928 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 40 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 41 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 42 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 43 nsew signal tristate
flabel metal3 s 26200 8440 27000 8560 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 44 nsew signal tristate
flabel metal3 s 26200 1096 27000 1216 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 45 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 46 nsew signal tristate
flabel metal3 s 26200 9256 27000 9376 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 47 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 48 nsew signal tristate
flabel metal3 s 26200 10072 27000 10192 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 49 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 50 nsew signal tristate
flabel metal3 s 26200 10888 27000 11008 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 51 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 52 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 53 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 54 nsew signal tristate
flabel metal3 s 26200 12520 27000 12640 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 55 nsew signal tristate
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 56 nsew signal tristate
flabel metal3 s 26200 1912 27000 2032 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 57 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 58 nsew signal tristate
flabel metal3 s 26200 2728 27000 2848 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 59 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 60 nsew signal tristate
flabel metal3 s 26200 3544 27000 3664 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 61 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 62 nsew signal tristate
flabel metal3 s 26200 4360 27000 4480 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 63 nsew signal tristate
flabel metal2 s 12714 26200 12770 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 64 nsew signal input
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 65 nsew signal input
flabel metal2 s 16762 26200 16818 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 66 nsew signal input
flabel metal2 s 17130 26200 17186 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 67 nsew signal input
flabel metal2 s 17498 26200 17554 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 68 nsew signal input
flabel metal2 s 17866 26200 17922 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 69 nsew signal input
flabel metal2 s 18234 26200 18290 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 70 nsew signal input
flabel metal2 s 18602 26200 18658 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 71 nsew signal input
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 72 nsew signal input
flabel metal2 s 19338 26200 19394 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 73 nsew signal input
flabel metal2 s 19706 26200 19762 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 74 nsew signal input
flabel metal2 s 13082 26200 13138 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 75 nsew signal input
flabel metal2 s 20074 26200 20130 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 76 nsew signal input
flabel metal2 s 20442 26200 20498 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 77 nsew signal input
flabel metal2 s 20810 26200 20866 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 78 nsew signal input
flabel metal2 s 21178 26200 21234 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 79 nsew signal input
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 80 nsew signal input
flabel metal2 s 21914 26200 21970 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 81 nsew signal input
flabel metal2 s 22282 26200 22338 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 82 nsew signal input
flabel metal2 s 22650 26200 22706 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 83 nsew signal input
flabel metal2 s 23018 26200 23074 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 84 nsew signal input
flabel metal2 s 23386 26200 23442 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 85 nsew signal input
flabel metal2 s 13450 26200 13506 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 86 nsew signal input
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 87 nsew signal input
flabel metal2 s 14186 26200 14242 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 88 nsew signal input
flabel metal2 s 14554 26200 14610 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 89 nsew signal input
flabel metal2 s 14922 26200 14978 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 90 nsew signal input
flabel metal2 s 15290 26200 15346 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 91 nsew signal input
flabel metal2 s 15658 26200 15714 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 92 nsew signal input
flabel metal2 s 16026 26200 16082 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 93 nsew signal input
flabel metal2 s 1674 26200 1730 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 94 nsew signal tristate
flabel metal2 s 5354 26200 5410 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 95 nsew signal tristate
flabel metal2 s 5722 26200 5778 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 96 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 97 nsew signal tristate
flabel metal2 s 6458 26200 6514 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 98 nsew signal tristate
flabel metal2 s 6826 26200 6882 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 99 nsew signal tristate
flabel metal2 s 7194 26200 7250 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 100 nsew signal tristate
flabel metal2 s 7562 26200 7618 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 101 nsew signal tristate
flabel metal2 s 7930 26200 7986 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 102 nsew signal tristate
flabel metal2 s 8298 26200 8354 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 103 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 104 nsew signal tristate
flabel metal2 s 2042 26200 2098 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 105 nsew signal tristate
flabel metal2 s 9034 26200 9090 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 106 nsew signal tristate
flabel metal2 s 9402 26200 9458 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 107 nsew signal tristate
flabel metal2 s 9770 26200 9826 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 108 nsew signal tristate
flabel metal2 s 10138 26200 10194 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 109 nsew signal tristate
flabel metal2 s 10506 26200 10562 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 110 nsew signal tristate
flabel metal2 s 10874 26200 10930 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 111 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 112 nsew signal tristate
flabel metal2 s 11610 26200 11666 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 113 nsew signal tristate
flabel metal2 s 11978 26200 12034 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 114 nsew signal tristate
flabel metal2 s 12346 26200 12402 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 115 nsew signal tristate
flabel metal2 s 2410 26200 2466 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 116 nsew signal tristate
flabel metal2 s 2778 26200 2834 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 117 nsew signal tristate
flabel metal2 s 3146 26200 3202 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 118 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 119 nsew signal tristate
flabel metal2 s 3882 26200 3938 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 120 nsew signal tristate
flabel metal2 s 4250 26200 4306 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 121 nsew signal tristate
flabel metal2 s 4618 26200 4674 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 122 nsew signal tristate
flabel metal2 s 4986 26200 5042 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 123 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 prog_clk
port 124 nsew signal input
flabel metal2 s 24490 26200 24546 27000 0 FreeSans 224 90 0 0 prog_reset
port 125 nsew signal input
flabel metal2 s 24858 26200 24914 27000 0 FreeSans 224 90 0 0 reset
port 126 nsew signal input
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 26200 25576 27000 25696 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 26200 26392 27000 26512 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 25226 26200 25282 27000 0 FreeSans 224 90 0 0 test_enable
port 131 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
rlabel metal1 13478 23936 13478 23936 0 VGND
rlabel metal1 13478 24480 13478 24480 0 VPWR
rlabel metal1 8924 2414 8924 2414 0 ccff_head
rlabel metal3 25630 340 25630 340 0 ccff_tail
rlabel metal1 19826 4114 19826 4114 0 chanx_right_in[0]
rlabel metal1 4002 19346 4002 19346 0 chanx_right_in[10]
rlabel metal2 2898 15351 2898 15351 0 chanx_right_in[11]
rlabel metal3 20700 17816 20700 17816 0 chanx_right_in[12]
rlabel metal4 17204 16184 17204 16184 0 chanx_right_in[13]
rlabel metal2 2576 19108 2576 19108 0 chanx_right_in[14]
rlabel metal1 2277 19754 2277 19754 0 chanx_right_in[15]
rlabel metal4 21988 16048 21988 16048 0 chanx_right_in[16]
rlabel metal1 18768 4590 18768 4590 0 chanx_right_in[17]
rlabel metal2 20746 15844 20746 15844 0 chanx_right_in[18]
rlabel metal2 21022 24497 21022 24497 0 chanx_right_in[19]
rlabel metal1 19458 12614 19458 12614 0 chanx_right_in[1]
rlabel metal3 15709 2380 15709 2380 0 chanx_right_in[20]
rlabel metal2 14490 7769 14490 7769 0 chanx_right_in[21]
rlabel metal2 18952 12852 18952 12852 0 chanx_right_in[22]
rlabel metal3 26090 22372 26090 22372 0 chanx_right_in[23]
rlabel metal3 17871 11220 17871 11220 0 chanx_right_in[24]
rlabel metal4 16468 10268 16468 10268 0 chanx_right_in[25]
rlabel metal1 17894 6902 17894 6902 0 chanx_right_in[26]
rlabel metal3 15962 12444 15962 12444 0 chanx_right_in[27]
rlabel metal2 22034 25109 22034 25109 0 chanx_right_in[28]
rlabel metal4 15180 23596 15180 23596 0 chanx_right_in[29]
rlabel metal1 19504 6426 19504 6426 0 chanx_right_in[2]
rlabel metal1 17066 5134 17066 5134 0 chanx_right_in[3]
rlabel metal1 16882 15878 16882 15878 0 chanx_right_in[4]
rlabel metal1 19274 14858 19274 14858 0 chanx_right_in[5]
rlabel metal2 16974 4046 16974 4046 0 chanx_right_in[6]
rlabel metal1 6532 20230 6532 20230 0 chanx_right_in[7]
rlabel metal1 21942 16558 21942 16558 0 chanx_right_in[8]
rlabel metal2 23230 16711 23230 16711 0 chanx_right_in[9]
rlabel metal3 25722 748 25722 748 0 chanx_right_out[0]
rlabel metal1 24104 5270 24104 5270 0 chanx_right_out[10]
rlabel metal2 24610 4097 24610 4097 0 chanx_right_out[11]
rlabel metal3 25676 5644 25676 5644 0 chanx_right_out[12]
rlabel metal2 24794 5049 24794 5049 0 chanx_right_out[13]
rlabel metal3 26044 6460 26044 6460 0 chanx_right_out[14]
rlabel metal2 23322 7089 23322 7089 0 chanx_right_out[15]
rlabel metal2 24702 6205 24702 6205 0 chanx_right_out[16]
rlabel metal3 25676 7684 25676 7684 0 chanx_right_out[17]
rlabel metal1 23368 8398 23368 8398 0 chanx_right_out[18]
rlabel metal2 24794 7361 24794 7361 0 chanx_right_out[19]
rlabel metal3 24894 1156 24894 1156 0 chanx_right_out[1]
rlabel metal3 25676 8908 25676 8908 0 chanx_right_out[20]
rlabel metal1 24104 9622 24104 9622 0 chanx_right_out[21]
rlabel metal1 24794 7344 24794 7344 0 chanx_right_out[22]
rlabel metal1 24104 10574 24104 10574 0 chanx_right_out[23]
rlabel metal2 25162 9537 25162 9537 0 chanx_right_out[24]
rlabel metal2 25162 10829 25162 10829 0 chanx_right_out[25]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[26]
rlabel metal2 24794 10625 24794 10625 0 chanx_right_out[27]
rlabel metal1 24472 11186 24472 11186 0 chanx_right_out[28]
rlabel metal3 25768 12580 25768 12580 0 chanx_right_out[29]
rlabel metal3 24342 1564 24342 1564 0 chanx_right_out[2]
rlabel metal3 24296 1972 24296 1972 0 chanx_right_out[3]
rlabel metal3 25676 2380 25676 2380 0 chanx_right_out[4]
rlabel metal1 24104 3094 24104 3094 0 chanx_right_out[5]
rlabel metal3 26044 3196 26044 3196 0 chanx_right_out[6]
rlabel metal1 23322 4012 23322 4012 0 chanx_right_out[7]
rlabel metal2 23414 4267 23414 4267 0 chanx_right_out[8]
rlabel metal3 25676 4420 25676 4420 0 chanx_right_out[9]
rlabel metal1 12972 22610 12972 22610 0 chany_top_in[0]
rlabel metal1 2162 10710 2162 10710 0 chany_top_in[10]
rlabel metal3 736 25092 736 25092 0 chany_top_in[11]
rlabel metal2 12788 14212 12788 14212 0 chany_top_in[12]
rlabel metal2 1610 25262 1610 25262 0 chany_top_in[13]
rlabel metal1 16468 24174 16468 24174 0 chany_top_in[14]
rlabel metal2 17986 25789 17986 25789 0 chany_top_in[15]
rlabel metal2 18630 26037 18630 26037 0 chany_top_in[16]
rlabel metal2 2070 11475 2070 11475 0 chany_top_in[17]
rlabel metal2 2484 18972 2484 18972 0 chany_top_in[18]
rlabel metal4 736 26180 736 26180 0 chany_top_in[19]
rlabel metal2 782 16966 782 16966 0 chany_top_in[1]
rlabel metal2 20102 26105 20102 26105 0 chany_top_in[20]
rlabel metal2 1242 21148 1242 21148 0 chany_top_in[21]
rlabel metal3 18561 23324 18561 23324 0 chany_top_in[22]
rlabel metal2 20930 26027 20930 26027 0 chany_top_in[23]
rlabel metal2 21298 26265 21298 26265 0 chany_top_in[24]
rlabel metal2 21942 25629 21942 25629 0 chany_top_in[25]
rlabel metal3 2047 21692 2047 21692 0 chany_top_in[26]
rlabel metal1 2346 10608 2346 10608 0 chany_top_in[27]
rlabel metal1 10350 9418 10350 9418 0 chany_top_in[28]
rlabel metal2 16606 7021 16606 7021 0 chany_top_in[29]
rlabel metal4 1012 17272 1012 17272 0 chany_top_in[2]
rlabel metal4 828 17068 828 17068 0 chany_top_in[3]
rlabel metal2 14214 26122 14214 26122 0 chany_top_in[4]
rlabel metal2 1150 17340 1150 17340 0 chany_top_in[5]
rlabel metal2 1564 15572 1564 15572 0 chany_top_in[6]
rlabel metal1 17020 3502 17020 3502 0 chany_top_in[7]
rlabel metal2 15541 26316 15541 26316 0 chany_top_in[8]
rlabel metal2 12558 22984 12558 22984 0 chany_top_in[9]
rlabel metal1 1932 19278 1932 19278 0 chany_top_out[0]
rlabel metal1 4692 23630 4692 23630 0 chany_top_out[10]
rlabel metal2 5750 24490 5750 24490 0 chany_top_out[11]
rlabel metal1 6210 21930 6210 21930 0 chany_top_out[12]
rlabel metal1 4876 24242 4876 24242 0 chany_top_out[13]
rlabel metal1 7130 21454 7130 21454 0 chany_top_out[14]
rlabel metal1 7544 21454 7544 21454 0 chany_top_out[15]
rlabel metal1 6716 23630 6716 23630 0 chany_top_out[16]
rlabel metal1 7084 23154 7084 23154 0 chany_top_out[17]
rlabel metal1 8188 22066 8188 22066 0 chany_top_out[18]
rlabel metal1 7268 24106 7268 24106 0 chany_top_out[19]
rlabel metal2 2070 23538 2070 23538 0 chany_top_out[1]
rlabel metal2 8786 24497 8786 24497 0 chany_top_out[20]
rlabel metal1 8786 23154 8786 23154 0 chany_top_out[21]
rlabel metal1 9062 24242 9062 24242 0 chany_top_out[22]
rlabel metal1 9384 23698 9384 23698 0 chany_top_out[23]
rlabel metal1 11316 21930 11316 21930 0 chany_top_out[24]
rlabel metal2 10902 25000 10902 25000 0 chany_top_out[25]
rlabel metal1 11132 24242 11132 24242 0 chany_top_out[26]
rlabel metal2 14766 24582 14766 24582 0 chany_top_out[27]
rlabel metal2 12006 24966 12006 24966 0 chany_top_out[28]
rlabel via1 12466 24259 12466 24259 0 chany_top_out[29]
rlabel metal2 2714 24888 2714 24888 0 chany_top_out[2]
rlabel metal2 2944 20366 2944 20366 0 chany_top_out[3]
rlabel metal1 3312 22066 3312 22066 0 chany_top_out[4]
rlabel metal2 3542 23878 3542 23878 0 chany_top_out[5]
rlabel metal2 4140 21964 4140 21964 0 chany_top_out[6]
rlabel metal1 4094 22678 4094 22678 0 chany_top_out[7]
rlabel metal1 3956 23154 3956 23154 0 chany_top_out[8]
rlabel metal2 5067 26316 5067 26316 0 chany_top_out[9]
rlabel metal1 21206 18326 21206 18326 0 clknet_0_prog_clk
rlabel metal2 11730 16320 11730 16320 0 clknet_3_0__leaf_prog_clk
rlabel metal1 15640 15538 15640 15538 0 clknet_3_1__leaf_prog_clk
rlabel metal2 8970 20978 8970 20978 0 clknet_3_2__leaf_prog_clk
rlabel metal1 14950 18734 14950 18734 0 clknet_3_3__leaf_prog_clk
rlabel metal2 19366 14484 19366 14484 0 clknet_3_4__leaf_prog_clk
rlabel metal1 20884 16626 20884 16626 0 clknet_3_5__leaf_prog_clk
rlabel metal2 20286 19890 20286 19890 0 clknet_3_6__leaf_prog_clk
rlabel metal2 18446 17374 18446 17374 0 clknet_3_7__leaf_prog_clk
rlabel metal1 7176 2618 7176 2618 0 net1
rlabel metal2 17986 4505 17986 4505 0 net10
rlabel metal1 3496 14382 3496 14382 0 net100
rlabel metal1 19642 22066 19642 22066 0 net101
rlabel metal1 6026 23086 6026 23086 0 net102
rlabel metal2 7406 21556 7406 21556 0 net103
rlabel metal1 4830 24106 4830 24106 0 net104
rlabel metal1 4094 19924 4094 19924 0 net105
rlabel metal1 6992 22542 6992 22542 0 net106
rlabel metal2 1886 14348 1886 14348 0 net107
rlabel metal3 5727 19244 5727 19244 0 net108
rlabel metal2 3818 15453 3818 15453 0 net109
rlabel metal1 6716 12954 6716 12954 0 net11
rlabel metal1 6716 20910 6716 20910 0 net110
rlabel metal1 5060 13702 5060 13702 0 net111
rlabel metal2 2070 17035 2070 17035 0 net112
rlabel metal1 6348 12614 6348 12614 0 net113
rlabel metal2 7314 17204 7314 17204 0 net114
rlabel metal2 2346 11696 2346 11696 0 net115
rlabel via2 2254 20893 2254 20893 0 net116
rlabel metal1 3680 20434 3680 20434 0 net117
rlabel metal1 1978 21998 1978 21998 0 net118
rlabel metal2 2162 18564 2162 18564 0 net119
rlabel metal4 15180 17136 15180 17136 0 net12
rlabel via1 4094 20893 4094 20893 0 net120
rlabel metal1 3588 12818 3588 12818 0 net121
rlabel metal2 2254 23137 2254 23137 0 net122
rlabel metal1 12926 20400 12926 20400 0 net123
rlabel metal1 12367 13226 12367 13226 0 net124
rlabel metal1 16100 13906 16100 13906 0 net125
rlabel metal2 15870 17034 15870 17034 0 net126
rlabel metal1 19734 21862 19734 21862 0 net127
rlabel metal1 20141 16490 20141 16490 0 net128
rlabel metal3 20332 12920 20332 12920 0 net129
rlabel metal1 14950 13362 14950 13362 0 net13
rlabel via2 19458 15419 19458 15419 0 net130
rlabel metal1 20562 8534 20562 8534 0 net131
rlabel metal3 25507 19380 25507 19380 0 net132
rlabel metal1 12052 7514 12052 7514 0 net133
rlabel via2 18906 12597 18906 12597 0 net134
rlabel metal1 18170 3570 18170 3570 0 net135
rlabel metal1 12926 6256 12926 6256 0 net136
rlabel metal1 18676 11254 18676 11254 0 net137
rlabel metal2 2622 12461 2622 12461 0 net138
rlabel metal1 19458 19686 19458 19686 0 net139
rlabel metal2 15318 21709 15318 21709 0 net14
rlabel metal1 18492 17714 18492 17714 0 net140
rlabel metal2 874 16932 874 16932 0 net141
rlabel metal4 2300 13464 2300 13464 0 net142
rlabel metal2 966 15725 966 15725 0 net143
rlabel metal1 9384 19686 9384 19686 0 net144
rlabel metal1 18538 22610 18538 22610 0 net145
rlabel metal3 9936 19652 9936 19652 0 net146
rlabel metal1 11868 20502 11868 20502 0 net147
rlabel metal1 2208 12206 2208 12206 0 net148
rlabel metal1 14168 19686 14168 19686 0 net149
rlabel metal1 17986 21998 17986 21998 0 net15
rlabel metal1 2116 8602 2116 8602 0 net150
rlabel metal2 11178 16337 11178 16337 0 net151
rlabel metal2 12742 14824 12742 14824 0 net152
rlabel metal1 14628 16082 14628 16082 0 net153
rlabel metal1 13846 17578 13846 17578 0 net154
rlabel via2 1794 24021 1794 24021 0 net155
rlabel metal4 2484 18224 2484 18224 0 net156
rlabel via2 19366 20213 19366 20213 0 net157
rlabel metal1 23782 17578 23782 17578 0 net158
rlabel metal1 16836 1870 16836 1870 0 net159
rlabel metal3 16192 15028 16192 15028 0 net16
rlabel metal2 12926 6511 12926 6511 0 net160
rlabel metal2 16422 4658 16422 4658 0 net161
rlabel metal1 13156 5542 13156 5542 0 net162
rlabel metal1 19688 13158 19688 13158 0 net163
rlabel metal1 20332 13838 20332 13838 0 net164
rlabel metal1 20792 15470 20792 15470 0 net165
rlabel metal2 7406 3468 7406 3468 0 net166
rlabel metal1 9614 6426 9614 6426 0 net167
rlabel metal2 2622 15300 2622 15300 0 net168
rlabel metal1 20240 6766 20240 6766 0 net169
rlabel metal3 19780 16524 19780 16524 0 net17
rlabel metal1 17940 6290 17940 6290 0 net170
rlabel metal2 3818 17476 3818 17476 0 net171
rlabel metal2 12190 12342 12190 12342 0 net172
rlabel metal1 2070 18292 2070 18292 0 net173
rlabel metal1 21068 17306 21068 17306 0 net174
rlabel metal1 25300 12614 25300 12614 0 net175
rlabel metal1 24932 8942 24932 8942 0 net176
rlabel metal2 19182 10846 19182 10846 0 net177
rlabel metal2 10534 16252 10534 16252 0 net178
rlabel metal1 24196 15674 24196 15674 0 net179
rlabel metal3 18331 20332 18331 20332 0 net18
rlabel metal2 14582 8772 14582 8772 0 net180
rlabel metal1 22126 10234 22126 10234 0 net181
rlabel metal1 24932 3502 24932 3502 0 net182
rlabel metal1 15962 8942 15962 8942 0 net183
rlabel metal2 18630 8772 18630 8772 0 net184
rlabel metal2 1702 17850 1702 17850 0 net185
rlabel metal1 2300 18598 2300 18598 0 net186
rlabel metal2 5750 19210 5750 19210 0 net187
rlabel metal2 19274 7599 19274 7599 0 net188
rlabel metal2 13202 14212 13202 14212 0 net189
rlabel metal2 20010 24616 20010 24616 0 net19
rlabel metal1 25208 2618 25208 2618 0 net190
rlabel metal1 4968 17850 4968 17850 0 net191
rlabel metal1 12673 10642 12673 10642 0 net192
rlabel metal1 14490 11866 14490 11866 0 net193
rlabel metal1 4600 16218 4600 16218 0 net194
rlabel metal2 6026 19958 6026 19958 0 net195
rlabel metal1 18538 6970 18538 6970 0 net196
rlabel metal2 20608 12852 20608 12852 0 net197
rlabel metal1 16238 10778 16238 10778 0 net198
rlabel metal1 10258 11730 10258 11730 0 net199
rlabel metal2 19458 3417 19458 3417 0 net2
rlabel via2 16606 15691 16606 15691 0 net20
rlabel metal1 3312 21658 3312 21658 0 net200
rlabel metal1 17158 8058 17158 8058 0 net201
rlabel metal1 18308 10642 18308 10642 0 net202
rlabel metal1 15962 2482 15962 2482 0 net203
rlabel metal1 6210 13838 6210 13838 0 net204
rlabel metal2 10534 15164 10534 15164 0 net205
rlabel metal2 13294 6426 13294 6426 0 net206
rlabel metal2 17986 9350 17986 9350 0 net207
rlabel metal1 13248 23086 13248 23086 0 net208
rlabel metal2 12374 11985 12374 11985 0 net209
rlabel via2 20838 22627 20838 22627 0 net21
rlabel metal1 26082 13498 26082 13498 0 net210
rlabel metal1 5888 17850 5888 17850 0 net211
rlabel metal1 8326 17170 8326 17170 0 net212
rlabel metal1 15686 8500 15686 8500 0 net213
rlabel metal1 6210 13158 6210 13158 0 net214
rlabel metal1 16468 12954 16468 12954 0 net215
rlabel metal1 6670 20434 6670 20434 0 net216
rlabel metal2 2622 21488 2622 21488 0 net217
rlabel metal1 9200 16082 9200 16082 0 net218
rlabel metal1 17848 10030 17848 10030 0 net219
rlabel metal1 18768 19686 18768 19686 0 net22
rlabel metal2 8602 14790 8602 14790 0 net220
rlabel metal2 19274 4862 19274 4862 0 net221
rlabel metal1 7728 19822 7728 19822 0 net222
rlabel metal2 2346 15436 2346 15436 0 net223
rlabel metal2 7682 17476 7682 17476 0 net224
rlabel metal1 20010 4794 20010 4794 0 net225
rlabel metal2 20102 8262 20102 8262 0 net226
rlabel metal1 6624 14586 6624 14586 0 net227
rlabel metal1 24840 4590 24840 4590 0 net228
rlabel metal1 20838 6800 20838 6800 0 net229
rlabel metal3 13961 22644 13961 22644 0 net23
rlabel metal2 10258 8976 10258 8976 0 net230
rlabel metal1 3864 15878 3864 15878 0 net231
rlabel metal1 9338 13838 9338 13838 0 net232
rlabel metal2 10902 21964 10902 21964 0 net233
rlabel metal1 6348 16558 6348 16558 0 net234
rlabel metal1 11914 17714 11914 17714 0 net235
rlabel metal2 2714 19907 2714 19907 0 net236
rlabel metal3 17940 20468 17940 20468 0 net237
rlabel metal2 13892 13532 13892 13532 0 net238
rlabel metal2 8510 3196 8510 3196 0 net239
rlabel metal2 15502 8075 15502 8075 0 net24
rlabel metal1 7406 2380 7406 2380 0 net240
rlabel metal1 8648 4794 8648 4794 0 net241
rlabel metal1 10442 8058 10442 8058 0 net242
rlabel metal1 4278 14926 4278 14926 0 net243
rlabel metal3 13340 22712 13340 22712 0 net244
rlabel metal1 19872 7378 19872 7378 0 net245
rlabel metal2 20378 9248 20378 9248 0 net246
rlabel metal1 12834 11696 12834 11696 0 net247
rlabel metal1 13202 12886 13202 12886 0 net248
rlabel metal1 20148 5202 20148 5202 0 net249
rlabel metal2 15640 14994 15640 14994 0 net25
rlabel via2 12742 9333 12742 9333 0 net250
rlabel metal2 4278 19244 4278 19244 0 net251
rlabel metal1 10258 18156 10258 18156 0 net252
rlabel metal1 21068 10778 21068 10778 0 net253
rlabel metal1 20562 9146 20562 9146 0 net254
rlabel metal2 15594 16218 15594 16218 0 net255
rlabel metal1 15272 17714 15272 17714 0 net256
rlabel metal3 13524 7208 13524 7208 0 net257
rlabel via2 21022 17595 21022 17595 0 net258
rlabel metal2 24610 11594 24610 11594 0 net259
rlabel metal1 19228 16218 19228 16218 0 net26
rlabel metal2 19734 16320 19734 16320 0 net260
rlabel metal1 21850 11118 21850 11118 0 net261
rlabel metal2 17250 11152 17250 11152 0 net262
rlabel metal2 9706 16626 9706 16626 0 net263
rlabel metal1 11730 16218 11730 16218 0 net264
rlabel metal2 5658 14654 5658 14654 0 net265
rlabel metal1 16008 8602 16008 8602 0 net266
rlabel metal2 20470 9860 20470 9860 0 net267
rlabel metal1 19642 15096 19642 15096 0 net268
rlabel metal1 21758 5678 21758 5678 0 net269
rlabel metal1 18676 14586 18676 14586 0 net27
rlabel metal2 25668 15164 25668 15164 0 net270
rlabel metal1 23690 15470 23690 15470 0 net271
rlabel via2 17250 15555 17250 15555 0 net272
rlabel metal1 15272 10234 15272 10234 0 net273
rlabel metal2 16882 10064 16882 10064 0 net274
rlabel metal1 18216 8058 18216 8058 0 net275
rlabel metal1 17434 12750 17434 12750 0 net276
rlabel metal1 20102 6222 20102 6222 0 net277
rlabel metal2 20470 19465 20470 19465 0 net278
rlabel metal2 1702 18564 1702 18564 0 net279
rlabel metal1 14674 14586 14674 14586 0 net28
rlabel metal2 10258 18224 10258 18224 0 net280
rlabel metal1 13754 12342 13754 12342 0 net281
rlabel metal1 14168 14314 14168 14314 0 net282
rlabel metal1 8924 15470 8924 15470 0 net283
rlabel metal2 11178 15538 11178 15538 0 net284
rlabel metal1 7820 13498 7820 13498 0 net285
rlabel metal1 8786 20366 8786 20366 0 net286
rlabel metal1 6440 15470 6440 15470 0 net287
rlabel metal3 17825 20876 17825 20876 0 net288
rlabel metal2 5382 19516 5382 19516 0 net289
rlabel metal2 15962 23324 15962 23324 0 net29
rlabel metal2 6026 20672 6026 20672 0 net290
rlabel metal1 20976 1938 20976 1938 0 net291
rlabel metal1 20470 3706 20470 3706 0 net292
rlabel metal1 7084 19482 7084 19482 0 net293
rlabel metal2 17434 19397 17434 19397 0 net294
rlabel metal1 4646 17680 4646 17680 0 net295
rlabel metal1 7268 18326 7268 18326 0 net296
rlabel metal1 5658 16218 5658 16218 0 net297
rlabel metal2 18630 21641 18630 21641 0 net298
rlabel metal1 16698 7820 16698 7820 0 net299
rlabel metal2 19366 23817 19366 23817 0 net3
rlabel metal1 21712 16422 21712 16422 0 net30
rlabel metal2 18630 9214 18630 9214 0 net300
rlabel metal2 9982 18496 9982 18496 0 net301
rlabel metal2 21344 12988 21344 12988 0 net302
rlabel metal2 1702 21964 1702 21964 0 net303
rlabel metal2 13754 22542 13754 22542 0 net304
rlabel metal2 13938 11900 13938 11900 0 net305
rlabel metal1 14950 13498 14950 13498 0 net306
rlabel metal3 18975 12852 18975 12852 0 net307
rlabel metal1 17296 14246 17296 14246 0 net308
rlabel metal1 11678 11730 11678 11730 0 net309
rlabel metal2 12558 16320 12558 16320 0 net31
rlabel metal2 11178 13090 11178 13090 0 net310
rlabel metal2 15134 10846 15134 10846 0 net311
rlabel metal1 14529 13702 14529 13702 0 net312
rlabel metal2 17342 9146 17342 9146 0 net313
rlabel metal1 18262 9622 18262 9622 0 net314
rlabel metal1 17756 6766 17756 6766 0 net315
rlabel metal1 22908 13362 22908 13362 0 net316
rlabel metal1 7130 14858 7130 14858 0 net317
rlabel metal1 19826 2618 19826 2618 0 net318
rlabel metal2 7590 14450 7590 14450 0 net319
rlabel metal1 17986 20978 17986 20978 0 net32
rlabel metal1 9752 22542 9752 22542 0 net320
rlabel metal2 15318 24038 15318 24038 0 net321
rlabel metal2 12834 21182 12834 21182 0 net322
rlabel metal1 7360 16218 7360 16218 0 net323
rlabel metal1 9729 17578 9729 17578 0 net324
rlabel metal1 17158 6800 17158 6800 0 net325
rlabel metal1 21850 13838 21850 13838 0 net326
rlabel via2 15134 7973 15134 7973 0 net327
rlabel via2 13846 15691 13846 15691 0 net328
rlabel metal1 15226 9656 15226 9656 0 net329
rlabel metal2 2438 7922 2438 7922 0 net33
rlabel metal2 21206 19363 21206 19363 0 net330
rlabel metal2 21574 6222 21574 6222 0 net331
rlabel metal2 13754 25211 13754 25211 0 net332
rlabel metal2 7866 18428 7866 18428 0 net333
rlabel metal1 10810 17272 10810 17272 0 net334
rlabel metal1 16008 12818 16008 12818 0 net335
rlabel metal1 16054 14042 16054 14042 0 net336
rlabel metal1 6670 21114 6670 21114 0 net337
rlabel metal1 13938 20536 13938 20536 0 net338
rlabel metal2 16974 10234 16974 10234 0 net339
rlabel metal1 25576 13838 25576 13838 0 net34
rlabel metal1 16100 13226 16100 13226 0 net340
rlabel metal1 8142 14382 8142 14382 0 net341
rlabel metal1 10810 14450 10810 14450 0 net342
rlabel metal1 24794 13294 24794 13294 0 net343
rlabel metal1 16100 18802 16100 18802 0 net344
rlabel metal2 8326 16252 8326 16252 0 net345
rlabel metal1 10524 15674 10524 15674 0 net346
rlabel metal2 6762 21148 6762 21148 0 net347
rlabel metal1 10212 19754 10212 19754 0 net348
rlabel metal1 2392 13498 2392 13498 0 net349
rlabel via2 13570 5355 13570 5355 0 net35
rlabel metal1 6870 23800 6870 23800 0 net350
rlabel metal1 18308 5202 18308 5202 0 net351
rlabel metal1 2162 22066 2162 22066 0 net352
rlabel metal2 19458 8058 19458 8058 0 net353
rlabel metal1 20930 8602 20930 8602 0 net354
rlabel metal1 20102 4590 20102 4590 0 net355
rlabel metal1 19044 6358 19044 6358 0 net356
rlabel metal2 7038 17884 7038 17884 0 net357
rlabel metal1 8510 17238 8510 17238 0 net358
rlabel metal2 2714 16354 2714 16354 0 net359
rlabel metal1 20976 19482 20976 19482 0 net36
rlabel metal2 14122 14654 14122 14654 0 net360
rlabel metal1 24932 6766 24932 6766 0 net361
rlabel metal1 24005 13702 24005 13702 0 net362
rlabel metal1 18446 5610 18446 5610 0 net363
rlabel metal1 21022 12104 21022 12104 0 net364
rlabel metal1 6854 14450 6854 14450 0 net365
rlabel metal1 6992 15674 6992 15674 0 net366
rlabel metal1 22540 6426 22540 6426 0 net367
rlabel metal1 20746 6630 20746 6630 0 net368
rlabel metal2 16238 7480 16238 7480 0 net369
rlabel metal1 20884 20570 20884 20570 0 net37
rlabel metal2 20010 19159 20010 19159 0 net370
rlabel metal1 8970 12954 8970 12954 0 net371
rlabel metal1 7084 19278 7084 19278 0 net372
rlabel metal1 8786 13906 8786 13906 0 net373
rlabel metal1 6854 18258 6854 18258 0 net374
rlabel metal1 25392 18394 25392 18394 0 net375
rlabel metal1 2070 17136 2070 17136 0 net376
rlabel via2 18906 5627 18906 5627 0 net377
rlabel metal2 12006 11764 12006 11764 0 net378
rlabel metal1 8142 3434 8142 3434 0 net379
rlabel metal2 21482 15113 21482 15113 0 net38
rlabel metal2 9154 3638 9154 3638 0 net380
rlabel metal1 5382 2482 5382 2482 0 net381
rlabel metal1 6946 2448 6946 2448 0 net382
rlabel metal1 8050 3706 8050 3706 0 net383
rlabel metal2 12466 16048 12466 16048 0 net39
rlabel metal2 15502 15215 15502 15215 0 net4
rlabel via2 1886 11611 1886 11611 0 net40
rlabel via2 19366 10251 19366 10251 0 net41
rlabel metal1 2254 9146 2254 9146 0 net42
rlabel metal1 20654 8874 20654 8874 0 net43
rlabel metal2 19642 18785 19642 18785 0 net44
rlabel metal1 13570 13940 13570 13940 0 net45
rlabel metal1 21850 12954 21850 12954 0 net46
rlabel metal2 20378 16915 20378 16915 0 net47
rlabel metal2 17250 17340 17250 17340 0 net48
rlabel metal1 24380 23290 24380 23290 0 net49
rlabel metal2 12650 15844 12650 15844 0 net5
rlabel via2 2438 11067 2438 11067 0 net50
rlabel via2 17434 24259 17434 24259 0 net51
rlabel via2 20470 14229 20470 14229 0 net52
rlabel metal1 14766 12682 14766 12682 0 net53
rlabel metal1 21620 11118 21620 11118 0 net54
rlabel metal2 16146 15113 16146 15113 0 net55
rlabel metal2 18078 9146 18078 9146 0 net56
rlabel metal1 19734 16082 19734 16082 0 net57
rlabel metal1 21022 18258 21022 18258 0 net58
rlabel via3 18515 18020 18515 18020 0 net59
rlabel via2 17618 19669 17618 19669 0 net6
rlabel metal1 17020 18190 17020 18190 0 net60
rlabel metal1 16100 1802 16100 1802 0 net61
rlabel metal1 18630 17102 18630 17102 0 net62
rlabel metal1 20102 2380 20102 2380 0 net63
rlabel metal1 21068 3026 21068 3026 0 net64
rlabel metal1 25162 14790 25162 14790 0 net65
rlabel metal1 25300 18870 25300 18870 0 net66
rlabel metal1 21413 5542 21413 5542 0 net67
rlabel metal2 23506 5236 23506 5236 0 net68
rlabel metal2 16790 6256 16790 6256 0 net69
rlabel metal2 15134 19091 15134 19091 0 net7
rlabel metal2 18078 7140 18078 7140 0 net70
rlabel metal1 12834 6188 12834 6188 0 net71
rlabel via2 22862 7837 22862 7837 0 net72
rlabel metal4 12604 10472 12604 10472 0 net73
rlabel via3 19757 18020 19757 18020 0 net74
rlabel metal1 21482 3502 21482 3502 0 net75
rlabel metal2 19642 8772 19642 8772 0 net76
rlabel metal1 17250 7956 17250 7956 0 net77
rlabel metal2 10442 8721 10442 8721 0 net78
rlabel metal2 21758 10234 21758 10234 0 net79
rlabel metal1 19228 21930 19228 21930 0 net8
rlabel metal2 10902 9809 10902 9809 0 net80
rlabel metal1 20930 7854 20930 7854 0 net81
rlabel metal1 17158 7276 17158 7276 0 net82
rlabel metal1 20930 9554 20930 9554 0 net83
rlabel via2 10626 9571 10626 9571 0 net84
rlabel metal2 13294 8806 13294 8806 0 net85
rlabel metal1 16422 14858 16422 14858 0 net86
rlabel metal1 18446 2992 18446 2992 0 net87
rlabel metal2 22678 2244 22678 2244 0 net88
rlabel metal1 22080 2618 22080 2618 0 net89
rlabel metal2 3358 20417 3358 20417 0 net9
rlabel metal1 20470 4488 20470 4488 0 net90
rlabel metal2 17802 4828 17802 4828 0 net91
rlabel metal1 21022 4624 21022 4624 0 net92
rlabel metal1 22402 14858 22402 14858 0 net93
rlabel metal2 1978 21199 1978 21199 0 net94
rlabel metal3 16284 23800 16284 23800 0 net95
rlabel metal4 12788 23528 12788 23528 0 net96
rlabel metal2 5474 20009 5474 20009 0 net97
rlabel metal1 2300 24174 2300 24174 0 net98
rlabel metal2 4278 14450 4278 14450 0 net99
rlabel metal1 18078 16082 18078 16082 0 prog_clk
rlabel metal1 12742 15028 12742 15028 0 prog_reset
rlabel metal1 16734 18258 16734 18258 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 18446 18462 18446 18462 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 19596 15164 19596 15164 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 15272 12614 15272 12614 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 14858 14994 14858 14994 0 sb_0__0_.mem_right_track_0.ccff_head
rlabel metal1 17940 19142 17940 19142 0 sb_0__0_.mem_right_track_0.ccff_tail
rlabel metal1 18262 21012 18262 21012 0 sb_0__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 25162 18751 25162 18751 0 sb_0__0_.mem_right_track_10.ccff_head
rlabel metal1 23552 17102 23552 17102 0 sb_0__0_.mem_right_track_10.ccff_tail
rlabel metal2 18998 10319 18998 10319 0 sb_0__0_.mem_right_track_10.mem_out\[0\]
rlabel metal2 21206 14892 21206 14892 0 sb_0__0_.mem_right_track_12.ccff_tail
rlabel metal1 21390 12954 21390 12954 0 sb_0__0_.mem_right_track_12.mem_out\[0\]
rlabel metal1 16882 8398 16882 8398 0 sb_0__0_.mem_right_track_14.ccff_tail
rlabel metal1 16606 17578 16606 17578 0 sb_0__0_.mem_right_track_14.mem_out\[0\]
rlabel metal2 19274 10506 19274 10506 0 sb_0__0_.mem_right_track_16.ccff_tail
rlabel metal1 24472 14926 24472 14926 0 sb_0__0_.mem_right_track_16.mem_out\[0\]
rlabel metal2 14858 10132 14858 10132 0 sb_0__0_.mem_right_track_18.ccff_tail
rlabel metal1 19044 10098 19044 10098 0 sb_0__0_.mem_right_track_18.mem_out\[0\]
rlabel metal1 19734 5236 19734 5236 0 sb_0__0_.mem_right_track_2.ccff_tail
rlabel metal1 16560 19142 16560 19142 0 sb_0__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 20332 9554 20332 9554 0 sb_0__0_.mem_right_track_28.ccff_tail
rlabel metal1 23598 6324 23598 6324 0 sb_0__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 21390 15504 21390 15504 0 sb_0__0_.mem_right_track_30.ccff_tail
rlabel metal1 21597 14858 21597 14858 0 sb_0__0_.mem_right_track_30.mem_out\[0\]
rlabel metal1 20194 15572 20194 15572 0 sb_0__0_.mem_right_track_32.ccff_tail
rlabel metal1 4278 21964 4278 21964 0 sb_0__0_.mem_right_track_32.mem_out\[0\]
rlabel metal1 21068 14450 21068 14450 0 sb_0__0_.mem_right_track_34.ccff_tail
rlabel metal2 21482 15606 21482 15606 0 sb_0__0_.mem_right_track_34.mem_out\[0\]
rlabel metal2 18998 13056 18998 13056 0 sb_0__0_.mem_right_track_4.ccff_tail
rlabel metal1 23690 19924 23690 19924 0 sb_0__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 17066 13158 17066 13158 0 sb_0__0_.mem_right_track_44.ccff_tail
rlabel metal1 18032 14586 18032 14586 0 sb_0__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 18906 12750 18906 12750 0 sb_0__0_.mem_right_track_46.ccff_tail
rlabel metal1 18078 18802 18078 18802 0 sb_0__0_.mem_right_track_46.mem_out\[0\]
rlabel metal1 21068 12750 21068 12750 0 sb_0__0_.mem_right_track_48.ccff_tail
rlabel metal2 19228 15062 19228 15062 0 sb_0__0_.mem_right_track_48.mem_out\[0\]
rlabel metal2 21114 8364 21114 8364 0 sb_0__0_.mem_right_track_50.mem_out\[0\]
rlabel metal1 16100 14450 16100 14450 0 sb_0__0_.mem_right_track_6.ccff_tail
rlabel metal1 18124 11050 18124 11050 0 sb_0__0_.mem_right_track_6.mem_out\[0\]
rlabel metal3 15732 13872 15732 13872 0 sb_0__0_.mem_right_track_8.mem_out\[0\]
rlabel metal2 16054 16932 16054 16932 0 sb_0__0_.mem_top_track_0.ccff_tail
rlabel metal1 19550 19890 19550 19890 0 sb_0__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 1702 22644 1702 22644 0 sb_0__0_.mem_top_track_10.ccff_head
rlabel via2 7866 20451 7866 20451 0 sb_0__0_.mem_top_track_10.ccff_tail
rlabel metal2 9614 21148 9614 21148 0 sb_0__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 13386 19958 13386 19958 0 sb_0__0_.mem_top_track_12.ccff_tail
rlabel metal1 14398 19142 14398 19142 0 sb_0__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 4554 20774 4554 20774 0 sb_0__0_.mem_top_track_14.ccff_tail
rlabel metal2 8878 20247 8878 20247 0 sb_0__0_.mem_top_track_14.mem_out\[0\]
rlabel metal2 10626 18972 10626 18972 0 sb_0__0_.mem_top_track_16.ccff_tail
rlabel metal2 12650 21216 12650 21216 0 sb_0__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 9706 19856 9706 19856 0 sb_0__0_.mem_top_track_18.ccff_tail
rlabel metal2 15594 19703 15594 19703 0 sb_0__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 18722 20230 18722 20230 0 sb_0__0_.mem_top_track_2.ccff_tail
rlabel metal1 17480 18870 17480 18870 0 sb_0__0_.mem_top_track_2.mem_out\[0\]
rlabel metal2 10994 16558 10994 16558 0 sb_0__0_.mem_top_track_28.ccff_tail
rlabel metal2 14122 18836 14122 18836 0 sb_0__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 12650 20281 12650 20281 0 sb_0__0_.mem_top_track_30.ccff_tail
rlabel via2 18354 19907 18354 19907 0 sb_0__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 12282 18190 12282 18190 0 sb_0__0_.mem_top_track_32.ccff_tail
rlabel metal2 9476 17102 9476 17102 0 sb_0__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 9982 15470 9982 15470 0 sb_0__0_.mem_top_track_34.ccff_tail
rlabel metal2 13478 16660 13478 16660 0 sb_0__0_.mem_top_track_34.mem_out\[0\]
rlabel metal2 1794 21301 1794 21301 0 sb_0__0_.mem_top_track_4.ccff_tail
rlabel metal2 20102 21505 20102 21505 0 sb_0__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 11224 14042 11224 14042 0 sb_0__0_.mem_top_track_44.ccff_tail
rlabel metal2 15962 15657 15962 15657 0 sb_0__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 13524 15538 13524 15538 0 sb_0__0_.mem_top_track_46.ccff_tail
rlabel metal1 14306 13430 14306 13430 0 sb_0__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 15272 13838 15272 13838 0 sb_0__0_.mem_top_track_48.ccff_tail
rlabel metal2 15042 13124 15042 13124 0 sb_0__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16422 14586 16422 14586 0 sb_0__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 1794 20468 1794 20468 0 sb_0__0_.mem_top_track_6.ccff_tail
rlabel metal2 17434 21709 17434 21709 0 sb_0__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 1518 13294 1518 13294 0 sb_0__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 11730 6188 11730 6188 0 sb_0__0_.mux_right_track_0.out
rlabel metal1 19228 19414 19228 19414 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19642 19856 19642 19856 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 18975 15164 18975 15164 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 9706 9894 9706 9894 0 sb_0__0_.mux_right_track_10.out
rlabel metal1 24150 17646 24150 17646 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18078 4828 18078 4828 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15870 3910 15870 3910 0 sb_0__0_.mux_right_track_12.out
rlabel metal2 21574 19006 21574 19006 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 21459 15708 21459 15708 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18078 3400 18078 3400 0 sb_0__0_.mux_right_track_14.out
rlabel metal1 23690 16218 23690 16218 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal4 21988 7616 21988 7616 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10994 5372 10994 5372 0 sb_0__0_.mux_right_track_16.out
rlabel metal1 25254 14382 25254 14382 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17802 3094 17802 3094 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15594 5644 15594 5644 0 sb_0__0_.mux_right_track_18.out
rlabel metal1 23460 14450 23460 14450 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13892 7854 13892 7854 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10810 7140 10810 7140 0 sb_0__0_.mux_right_track_2.out
rlabel metal2 18722 21597 18722 21597 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 4590 16284 4590 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18538 3910 18538 3910 0 sb_0__0_.mux_right_track_28.out
rlabel metal1 21298 13974 21298 13974 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19366 6256 19366 6256 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10764 7514 10764 7514 0 sb_0__0_.mux_right_track_30.out
rlabel metal2 21298 17884 21298 17884 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13984 13396 13984 13396 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19228 3706 19228 3706 0 sb_0__0_.mux_right_track_32.out
rlabel metal2 20102 17884 20102 17884 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 20171 15300 20171 15300 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20930 5508 20930 5508 0 sb_0__0_.mux_right_track_34.out
rlabel metal1 20194 14382 20194 14382 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 13770 17158 13770 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14490 17238 14490 17238 0 sb_0__0_.mux_right_track_4.out
rlabel metal1 24104 19754 24104 19754 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15502 18547 15502 18547 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17250 5338 17250 5338 0 sb_0__0_.mux_right_track_44.out
rlabel metal1 18492 13226 18492 13226 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18400 13430 18400 13430 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 18722 4352 18722 4352 0 sb_0__0_.mux_right_track_46.out
rlabel metal1 19550 12818 19550 12818 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14950 12648 14950 12648 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21206 2414 21206 2414 0 sb_0__0_.mux_right_track_48.out
rlabel metal1 20700 12954 20700 12954 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20148 2278 20148 2278 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17526 2618 17526 2618 0 sb_0__0_.mux_right_track_50.out
rlabel metal1 22218 15912 22218 15912 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21850 2006 21850 2006 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16790 4794 16790 4794 0 sb_0__0_.mux_right_track_6.out
rlabel metal1 24518 20842 24518 20842 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24610 21386 24610 21386 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 16514 5083 16514 5083 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19458 2142 19458 2142 0 sb_0__0_.mux_right_track_8.out
rlabel metal1 24840 24310 24840 24310 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19642 2465 19642 2465 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4278 9996 4278 9996 0 sb_0__0_.mux_top_track_0.out
rlabel metal1 14352 18938 14352 18938 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15318 19890 15318 19890 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 13432 15980 13432 15980 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7774 11322 7774 11322 0 sb_0__0_.mux_top_track_10.out
rlabel metal1 17986 21896 17986 21896 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 2714 11764 2714 11764 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2070 8058 2070 8058 0 sb_0__0_.mux_top_track_12.out
rlabel metal1 14628 21046 14628 21046 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 2622 7973 2622 7973 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5014 10098 5014 10098 0 sb_0__0_.mux_top_track_14.out
rlabel metal1 13478 21862 13478 21862 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12558 11288 12558 11288 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 1610 14076 1610 14076 0 sb_0__0_.mux_top_track_16.out
rlabel metal1 10442 21012 10442 21012 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 2162 14484 2162 14484 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6072 9418 6072 9418 0 sb_0__0_.mux_top_track_18.out
rlabel metal1 9798 19686 9798 19686 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8786 19686 8786 19686 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 7705 9588 7705 9588 0 sb_0__0_.mux_top_track_2.out
rlabel metal1 19504 22746 19504 22746 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18262 22746 18262 22746 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 2714 13141 2714 13141 0 sb_0__0_.mux_top_track_28.out
rlabel metal2 14766 19652 14766 19652 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel via3 10373 19516 10373 19516 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 2162 11390 2162 11390 0 sb_0__0_.mux_top_track_30.out
rlabel metal1 17480 20026 17480 20026 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 2346 9503 2346 9503 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5290 13838 5290 13838 0 sb_0__0_.mux_top_track_32.out
rlabel metal1 12282 18156 12282 18156 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11822 15237 11822 15237 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6256 11730 6256 11730 0 sb_0__0_.mux_top_track_34.out
rlabel metal1 15042 16966 15042 16966 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 4692 12852 4692 12852 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8556 8602 8556 8602 0 sb_0__0_.mux_top_track_4.out
rlabel metal1 19504 23834 19504 23834 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18170 24599 18170 24599 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3036 12750 3036 12750 0 sb_0__0_.mux_top_track_44.out
rlabel metal1 14582 16218 14582 16218 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4462 13498 4462 13498 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7728 10778 7728 10778 0 sb_0__0_.mux_top_track_46.out
rlabel metal1 13754 15402 13754 15402 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 14110 12466 14110 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 1518 12818 1518 12818 0 sb_0__0_.mux_top_track_48.out
rlabel metal1 17802 15946 17802 15946 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13800 13668 13800 13668 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6256 9350 6256 9350 0 sb_0__0_.mux_top_track_50.out
rlabel metal1 17066 17850 17066 17850 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7268 12818 7268 12818 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 1978 12750 1978 12750 0 sb_0__0_.mux_top_track_6.out
rlabel metal1 17296 21658 17296 21658 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18308 23086 18308 23086 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14122 16133 14122 16133 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 3542 10710 3542 10710 0 sb_0__0_.mux_top_track_8.out
rlabel metal1 18722 22406 18722 22406 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 14122 23579 14122 23579 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15226 21658 15226 21658 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 17204 17102 17204 17102 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 15732 18394 15732 18394 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 16698 18666 16698 18666 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 27000
<< end >>
