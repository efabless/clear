* NGSPICE file created from right_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

.subckt right_tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ ccff_head_0_0 ccff_head_1 ccff_head_2 ccff_tail ccff_tail_0 ccff_tail_1 chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23]
+ chanx_left_in[24] chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28]
+ chanx_left_in[29] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23]
+ chanx_left_out[24] chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28]
+ chanx_left_out[29] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21]
+ chany_bottom_in[22] chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25]
+ chany_bottom_in[26] chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29]
+ chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6]
+ chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10]
+ chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14]
+ chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18]
+ chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21]
+ chany_bottom_out[22] chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25]
+ chany_bottom_out[26] chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9]
+ chany_top_in_0[0] chany_top_in_0[10] chany_top_in_0[11] chany_top_in_0[12] chany_top_in_0[13]
+ chany_top_in_0[14] chany_top_in_0[15] chany_top_in_0[16] chany_top_in_0[17] chany_top_in_0[18]
+ chany_top_in_0[19] chany_top_in_0[1] chany_top_in_0[20] chany_top_in_0[21] chany_top_in_0[22]
+ chany_top_in_0[23] chany_top_in_0[24] chany_top_in_0[25] chany_top_in_0[26] chany_top_in_0[27]
+ chany_top_in_0[28] chany_top_in_0[29] chany_top_in_0[2] chany_top_in_0[3] chany_top_in_0[4]
+ chany_top_in_0[5] chany_top_in_0[6] chany_top_in_0[7] chany_top_in_0[8] chany_top_in_0[9]
+ chany_top_out_0[0] chany_top_out_0[10] chany_top_out_0[11] chany_top_out_0[12] chany_top_out_0[13]
+ chany_top_out_0[14] chany_top_out_0[15] chany_top_out_0[16] chany_top_out_0[17]
+ chany_top_out_0[18] chany_top_out_0[19] chany_top_out_0[1] chany_top_out_0[20] chany_top_out_0[21]
+ chany_top_out_0[22] chany_top_out_0[23] chany_top_out_0[24] chany_top_out_0[25]
+ chany_top_out_0[26] chany_top_out_0[27] chany_top_out_0[28] chany_top_out_0[29]
+ chany_top_out_0[2] chany_top_out_0[3] chany_top_out_0[4] chany_top_out_0[5] chany_top_out_0[6]
+ chany_top_out_0[7] chany_top_out_0[8] chany_top_out_0[9] clk0 gfpga_pad_io_soc_dir[0]
+ gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0]
+ gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0]
+ gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n left_width_0_height_0_subtile_0__pin_inpad_0_
+ left_width_0_height_0_subtile_1__pin_inpad_0_ left_width_0_height_0_subtile_2__pin_inpad_0_
+ left_width_0_height_0_subtile_3__pin_inpad_0_ prog_clk prog_reset reset right_width_0_height_0_subtile_0__pin_O_10_
+ right_width_0_height_0_subtile_0__pin_O_11_ right_width_0_height_0_subtile_0__pin_O_12_
+ right_width_0_height_0_subtile_0__pin_O_13_ right_width_0_height_0_subtile_0__pin_O_14_
+ right_width_0_height_0_subtile_0__pin_O_15_ right_width_0_height_0_subtile_0__pin_O_8_
+ right_width_0_height_0_subtile_0__pin_O_9_ sc_in sc_out test_enable top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ top_width_0_height_0_subtile_0__pin_O_0_
+ top_width_0_height_0_subtile_0__pin_O_1_ top_width_0_height_0_subtile_0__pin_O_2_
+ top_width_0_height_0_subtile_0__pin_O_3_ top_width_0_height_0_subtile_0__pin_O_4_
+ top_width_0_height_0_subtile_0__pin_O_5_ top_width_0_height_0_subtile_0__pin_O_6_
+ top_width_0_height_0_subtile_0__pin_O_7_ top_width_0_height_0_subtile_0__pin_cin_0_
+ top_width_0_height_0_subtile_0__pin_reg_in_0_
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk net542 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk
+ net818 net232 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_2__A0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk net765 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xhold351 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold340 sb_8__1_.mem_top_track_36.ccff_tail VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold362 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold373 sb_8__1_.mem_left_track_41.ccff_tail VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold395 sb_8__1_.mem_left_track_33.ccff_tail VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold384 sb_8__1_.mem_bottom_track_11.ccff_tail VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_leaf_53_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_2__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net286 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_2.mux_l2_in_3_ net350 net32 sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_23_prog_clk net825
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input92_A chany_top_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_294_ sb_8__1_.mux_left_track_3.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3_A reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__304__A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_2_ net7 net19 sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_59_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_17.mux_l1_in_0__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net290 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk net823
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_23.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold170 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net536
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_38_prog_clk net654 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold192 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold181 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk net687 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_33_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_346_ net47 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
Xsb_8__1_.mux_left_track_1.mux_l2_in_1__320 VGND VGND VPWR VPWR net320 sb_8__1_.mux_left_track_1.mux_l2_in_1__320/LO
+ sky130_fd_sc_hd__conb_1
X_277_ sb_8__1_.mux_left_track_37.out VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_23_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_39_prog_clk net463 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__A1 net429 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net231
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk net793
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput220 net220 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2__S cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_0__A0 sb_8__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_44_prog_clk
+ net862 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_8.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold504_A sb_8__1_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_29.mux_l1_in_1__330 VGND VGND VPWR VPWR net330 sb_8__1_.mux_left_track_29.mux_l1_in_1__330/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk net648 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input55_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_329_ sb_8__1_.mux_top_track_52.out VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__268
+ VGND VGND VPWR VPWR net268 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__268/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2_ net78 net47 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_2.mux_l4_in_0_ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X
+ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sb_8__1_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_5.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_2_ sb_8__1_.mux_left_track_21.out net14 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net391 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_0__A0 sb_8__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_0__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk net865
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_15.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
Xsb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_45_prog_clk sb_8__1_.mem_bottom_track_7.mem_out\[2\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold63_A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__312__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_45.mux_l1_in_0_ net221 net92 sb_8__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk
+ net858 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold41 cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X VGND VGND
+ VPWR VPWR net407 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold63 net86 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold52 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold74 chany_bottom_in[0] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_57.mux_l2_in_0_ net344 sb_8__1_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_0_X
+ cbx_8__1_.ccff_head VGND VGND VPWR VPWR sb_8__1_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold85 cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X VGND VGND
+ VPWR VPWR net451 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold96 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_input18_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_0__S sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_2__A0 sb_8__1_.mux_left_track_13.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_2.mux_l3_in_1_ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 net649 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__A0 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_0__S sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2__A0 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__307__A sb_8__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold511 cbx_8__1_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold500 sb_8__1_.mem_top_track_12.mem_out\[0\] VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold522 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR net888
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net458 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_13.mux_l2_in_0_ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_1_ net9 cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_25.mux_l1_in_0__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold26_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net532 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk
+ net852 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_36.mux_l2_in_1__353 VGND VGND VPWR VPWR net353 sb_8__1_.mux_top_track_36.mux_l2_in_1__353/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_2__A1 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk net556 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold341 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold352 cbx_8__1_.mem_top_ipin_11.ccff_tail VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xhold330 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold385 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold374 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold363 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR net729
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold396 sb_8__1_.mem_left_track_3.ccff_tail VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net97 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_26_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_2.mux_l2_in_2_ net14 net63 sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_26_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net379 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_8__1_.mem_top_track_2.mem_out\[1\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_293_ sb_8__1_.mux_left_track_5.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input85_A chany_top_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_13_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_29.mux_l2_in_1__313 VGND VGND VPWR VPWR net313 sb_8__1_.mux_bottom_track_29.mux_l2_in_1__313/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_52_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_1_ net212 left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_15.mux_l1_in_2_ sb_8__1_.mux_left_track_13.out net19 cbx_8__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA__320__A sb_8__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_17.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk net651
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_2__A0 net212 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold171 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold160 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold182 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold193 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_38_prog_clk net622 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_73_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_345_ sb_8__1_.mux_top_track_20.out VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_14_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_276_ net226 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_2__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_40_prog_clk net582 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_36.mem_out\[0\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__315__A sb_8__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.out sky130_fd_sc_hd__clkbuf_2
Xoutput210 net210 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ net403 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xoutput221 net221 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_44_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_1__S sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input48_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_3__S sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
X_328_ net57 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_46_prog_clk net583 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l1_in_1__A0 sb_8__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_3__238 VGND VGND VPWR VPWR net238 cbx_8__1_.mux_top_ipin_7.mux_l2_in_3__238/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_87_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input102_A net378 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2__A1 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__291
+ VGND VGND VPWR VPWR net291 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__291/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_2__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk net700
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_45_prog_clk sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_15.mux_l2_in_1__A1 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_45_prog_clk
+ net667 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_65_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__270
+ VGND VGND VPWR VPWR net270 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__270/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold31 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold20 chanx_left_in[10] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold64 cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X VGND VGND
+ VPWR VPWR net430 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold42 cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net408 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold53 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold97 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold75 cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X VGND VGND
+ VPWR VPWR net441 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_33.mux_l1_in_0__A0 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_2.mux_l3_in_0_ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_6 cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net270 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__mux2_8
Xsb_8__1_.mux_top_track_28.mux_l1_in_3__352 VGND VGND VPWR VPWR net352 sb_8__1_.mux_top_track_28.mux_l1_in_3__352/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__A1 net63 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2__A1 net68 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold501 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold512 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR net878
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__323__A sb_8__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold523 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[2\] VGND VGND VPWR VPWR net889
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_16_prog_clk net560
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_41.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_82_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ net424 VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_30_prog_clk net504 net233 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR
+ VPWR net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input30_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_13.mux_l2_in_1__322 VGND VGND VPWR VPWR net322 sb_8__1_.mux_left_track_13.mux_l2_in_1__322/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output117_A net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_3__359 VGND VGND VPWR VPWR net359 cbx_8__1_.mux_top_ipin_1.mux_l2_in_3__359/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_42_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3_ net255 sb_8__1_.mux_bottom_track_53.out
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_25.mux_l1_in_0__A1 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l2_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_0__A0 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ net790 net229 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_2__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__318__A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_15.mux_l3_in_0_ sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_15.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_57.mux_l1_in_0_ net227 net83 sb_8__1_.mem_left_track_57.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xhold320 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold331 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold353 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xhold342 cby_8__1_.cby_8__8_.mem_right_ipin_2.ccff_tail VGND VGND VPWR VPWR net708
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold386 sb_8__1_.mem_left_track_37.ccff_tail VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold364 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold375 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold397 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_2.mux_l2_in_1_ net49 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__1_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__A1 sb_8__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l2_in_3__A1 sb_8__1_.mux_left_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk net805
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_13_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net304 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_292_ sb_8__1_.mux_left_track_7.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input78_A chany_top_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_1__S sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_33.mux_l1_in_1__333 VGND VGND VPWR VPWR net333 sb_8__1_.mux_left_track_33.mux_l1_in_1__333/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_0_ net87 net73 sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_15.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_82_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_2__A0 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_20.mux_l1_in_3_ net351 net26 sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk net715
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_2__A1 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold150 cbx_8__1_.mem_top_ipin_2.ccff_tail VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__300
+ VGND VGND VPWR VPWR net300 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__300/LO
+ sky130_fd_sc_hd__conb_1
Xhold161 sb_8__1_.mem_bottom_track_53.ccff_tail VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold194 sb_8__1_.mem_left_track_41.mem_out\[0\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold183 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_38_prog_clk net609 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold172 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail
+ VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_92_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4_ net65 net63 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_344_ net44 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_275_ sb_8__1_.mux_left_track_41.out VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_2__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_41.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_41.out sky130_fd_sc_hd__buf_4
Xsb_8__1_.mux_bottom_track_37.mux_l3_in_0_ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_39_prog_clk net462 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_15.mux_l2_in_1_ net323 net222 sb_8__1_.mem_left_track_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2__A0 net74 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk net699
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput200 net200 VGND VGND VPWR VPWR chany_top_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
Xoutput211 net211 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
XFILLER_87_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__331__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_44_prog_clk
+ net851 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_25_prog_clk net627 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_23.mux_l2_in_1__A1 net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_327_ net56 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net723 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__326__A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_41.mux_l1_in_0__A0 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_35.out sky130_fd_sc_hd__clkbuf_1
XFILLER_55_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net271 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_37.mux_l2_in_1_ net315 net33 sb_8__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3_ net260 net429 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input60_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_1__A0 net63 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_78_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_20.mux_l3_in_0_ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_43_prog_clk net461 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net99 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net798 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_65_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold10 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold32 chany_bottom_in[5] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 net5 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold65 cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net431 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold43 cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold54 chanx_left_in[14] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold98 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_56_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold87 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold76 cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X VGND VGND
+ VPWR VPWR net442 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_33.mux_l1_in_0__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_30_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold502 cbx_8__1_.mem_top_ipin_5.mem_out\[2\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold524 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR net890
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold513 sb_8__1_.mem_left_track_15.mem_out\[1\] VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk net752
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_41.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_20.mux_l2_in_1_ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__D cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput111 net381 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput100 net370 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input23_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net299 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__mux2_4
XFILLER_44_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_3_ net359 sb_8__1_.mux_left_track_51.out cbx_8__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_71_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_2_ net57 cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__263
+ VGND VGND VPWR VPWR net263 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__263/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_0__S sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l4_in_0_ net430 cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_head VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__334__A net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold310 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold343 cbx_8__1_.mem_top_ipin_6.mem_out\[2\] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold332 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold321 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold365 sb_8__1_.mem_left_track_49.mem_out\[0\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold387 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold354 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold376 sb_8__1_.mem_bottom_track_3.ccff_tail VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold398 cby_8__1_.cby_8__8_.mem_left_ipin_3.ccff_tail VGND VGND VPWR VPWR net764
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_2.mux_l2_in_0_ net108 sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk net475
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ sb_8__1_.mux_left_track_9.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk net879
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_19.mux_l2_in_0__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_5.mux_l3_in_0_ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_output227_A net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk net857
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_15.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_2__A1 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_20.mux_l1_in_2_ net8 net20 sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk net784
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold151 sb_8__1_.mem_left_track_35.ccff_tail VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold162 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold140 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold184 sb_8__1_.mem_top_track_10.ccff_head VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold195 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold173 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_38_prog_clk net459 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_49.mux_l2_in_0__339 VGND VGND VPWR VPWR net339 sb_8__1_.mux_left_track_49.mux_l2_in_0__339/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3_ sb_8__1_.mux_bottom_track_29.out
+ net40 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3__A0 net73 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_343_ net43 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input90_A chany_top_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_274_ net88 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk net705
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_47.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1_A net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_40_prog_clk net664 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__244 VGND VGND VPWR VPWR net244 cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__244/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_15.mux_l2_in_0_ net40 sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_15.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2__A1 net43 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold79_A net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput201 net201 VGND VGND VPWR VPWR chany_top_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_2_3__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput212 net212 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk net512 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_1.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ net395 cbx_8__1_.mem_top_ipin_1.ccff_tail VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net787 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_2__S sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk
+ net574 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_5.mux_l2_in_1_ net340 net226 sb_8__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_25_prog_clk net611 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_326_ net45 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk net501 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_2__A0 net399 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l2_in_2__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__342__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk net717 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_3_ net237 sb_8__1_.mux_left_track_49.out cbx_8__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.out sky130_fd_sc_hd__buf_4
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_37.mux_l2_in_0_ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2_ net45 net66 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input53_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net117 net98 VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
Xsb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_44_prog_clk net533
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_44_prog_clk net624 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_309_ net69 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mux_top_ipin_1.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_6_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_3__S sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_3__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_2__S sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold11 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold22 cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X VGND VGND VPWR VPWR
+ net388 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 net59 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold44 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold55 net9 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold66 cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold88 chanx_left_in[23] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold77 cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net443 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold99 sb_8__1_.mem_left_track_11.ccff_head VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_57.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_57.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net99
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_8 net769 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__277
+ VGND VGND VPWR VPWR net277 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__277/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold525 sc_in VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold514 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold503 cbx_8__1_.mem_top_ipin_13.mem_out\[2\] VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_4_ sb_8__1_.mux_left_track_37.out net6 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_37.mux_l1_in_1_ net16 net215 sb_8__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_65_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_20.mux_l2_in_0_ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_1_prog_clk net860
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 net892 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput112 net374 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input16_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_2_ net28 sb_8__1_.mux_left_track_33.out cbx_8__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_8__1_.mux_top_ipin_6.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold311 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold300 cbx_8__1_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold333 sb_8__1_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold322 sb_8__1_.mem_top_track_12.ccff_tail VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold344 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold366 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold355 sb_8__1_.mem_top_track_4.ccff_tail VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold377 sb_8__1_.mem_bottom_track_29.ccff_tail VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold399 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold388 cby_8__1_.cby_8__8_.mem_left_ipin_1.ccff_tail VGND VGND VPWR VPWR net754
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk net561 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_290_ sb_8__1_.mux_left_track_11.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk net656
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net434 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk net846
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ net431 VGND VGND VPWR
+ VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__A1 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_20.mux_l1_in_1_ net56 net42 sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk net838
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold130 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold152 sb_8__1_.mem_bottom_track_21.ccff_tail VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold141 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold174 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold163 cbx_8__1_.mem_top_ipin_12.ccff_tail VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold185 sb_8__1_.mem_bottom_track_37.mem_out\[0\] VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk net634 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold196 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2_ net78 net47 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_1__S sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_342_ net42 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_273_ sb_8__1_.mux_left_track_45.out VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input83_A chany_top_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk net786
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_47.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_6.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_38_prog_clk net589 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk net525 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_top_track_2.mux_l1_in_0_ net105 net110 sb_8__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[2\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3_ net248 net93 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xoutput202 net202 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput224 net224 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
Xoutput213 net213 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk net749 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk
+ net819 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_5.mux_l2_in_0_ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_51_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_25_prog_clk net489 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_325_ sb_8__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_80_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net693 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__A1 net89 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk net847
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk net882 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_2_ net29 cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_0__S sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_1_ net35 cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_15.mux_l1_in_0_ net41 net70 sb_8__1_.mem_left_track_15.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_59_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk net704
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input46_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_44_prog_clk net792 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_27.mux_l1_in_1__A1 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_5.mux_l1_in_1__A0 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_308_ net68 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mux_top_ipin_1.mux_l3_in_0_ net394 cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mem_top_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_27.mux_l2_in_0_ sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_27.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_5.mux_l1_in_1_ net223 net48 sb_8__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold12 net380 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_1
Xhold23 cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X VGND VGND VPWR VPWR
+ net389 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X VGND VGND VPWR VPWR net422
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold45 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold34 cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X VGND VGND
+ VPWR VPWR net400 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold89 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold67 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold78 chanx_left_in[24] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input100_A net370 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net379 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_3_ net317 net28 sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_2_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_1__A0 sb_8__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net307 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold526 net372 VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold504 sb_8__1_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold515 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[2\] VGND VGND VPWR VPWR net881
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_hold54_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_3_ sb_8__1_.mux_left_track_25.out net12 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_2__S sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_37.mux_l1_in_0_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ net69 sb_8__1_.mem_bottom_track_37.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2_ net72 net41 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail net98 VGND
+ VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XANTENNA__348__A net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_4.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_88_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput102 net378 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_6
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_1_ net393 cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_27.mux_l1_in_1_ net329 net228 sb_8__1_.mem_left_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4__A0 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold301 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR net667
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold323 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold312 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold334 sb_8__1_.mem_left_track_27.ccff_tail VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold356 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold367 sb_8__1_.mem_left_track_7.ccff_tail VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold378 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold345 cbx_8__1_.mem_top_ipin_1.ccff_tail VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold389 sb_8__1_.mem_left_track_53.mem_out\[0\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk
+ net575 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk net526 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net281 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__mux2_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__251 VGND VGND VPWR VPWR net251
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__251/LO sky130_fd_sc_hd__conb_1
XFILLER_53_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net770
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk net564 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ net453 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_40_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__261
+ VGND VGND VPWR VPWR net261 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__261/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output115_A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk net490
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_32_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__284
+ VGND VGND VPWR VPWR net284 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__284/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_20.mux_l1_in_0_ net108 net110 sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_5.mux_l4_in_0_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_31_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk net811
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold142 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold131 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold153 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold120 sb_8__1_.mem_bottom_track_45.ccff_tail VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_1.mux_l1_in_2_ sb_8__1_.mux_left_track_15.out net18 cbx_8__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold186 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold175 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk net686 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold164 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold197 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_0__S sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk net803
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_3__S sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold525_A sc_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_341_ sb_8__1_.mux_top_track_28.out VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2__A0 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_272_ sb_8__1_.mux_left_track_47.out VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l2_in_2__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input76_A chany_top_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__271__A sb_8__1_.mux_left_track_49.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_6.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_44.mux_l3_in_0_ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.out sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net867 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ net822 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2_ net62 net70 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xoutput203 net203 VGND VGND VPWR VPWR chany_top_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput225 net225 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
Xoutput214 net214 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__356__A cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_TE_B
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_35.mux_l1_in_1__A1 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold475_A sb_8__1_.mem_top_track_52.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_26_prog_clk net584 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__266__A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_324_ sb_8__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__258 VGND VGND VPWR VPWR net258
+ cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__258/LO sky130_fd_sc_hd__conb_1
XFILLER_6_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_5.mux_l3_in_1_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold84_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3_ net244 net87 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk net778
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__248 VGND VGND VPWR VPWR net248
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__248/LO sky130_fd_sc_hd__conb_1
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_2_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_3_ net361 sb_8__1_.mux_left_track_53.out cbx_8__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk cbx_8__1_.mem_top_ipin_7.mem_out\[1\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_44.mux_l2_in_1_ net355 sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_top_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_44_prog_clk net779 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input39_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l2_in_3__A1 sb_8__1_.mux_left_track_49.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_5.mux_l1_in_1__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_307_ sb_8__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_load_slew229_A net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_5.mux_l1_in_0_ net54 net78 sb_8__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_80_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_0__A0 sb_8__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 net102 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_8
Xhold24 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold46 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold35 cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X VGND VGND
+ VPWR VPWR net401 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold57 cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X VGND VGND VPWR VPWR net423
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold68 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold79 net20 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2__A1 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_2_ net10 net22 sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4_ net93 net62 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold516 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold505 cbx_8__1_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_hold47_A chany_top_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_2_ sb_8__1_.mux_left_track_13.out net19 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net701 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_2__A0 sb_8__1_.mux_left_track_13.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_44.mux_l1_in_2_ net29 net11 sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA__364__A net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__273
+ VGND VGND VPWR VPWR net273 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__273/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_3__S sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput103 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_left_track_27.mux_l1_in_0_ net61 net91 sb_8__1_.mem_left_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_left_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__274__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4__A1 net63 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_3__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_11.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold302 cbx_8__1_.ccff_head VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold324 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold335 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold313 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_clkbuf_leaf_31_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold357 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold346 sb_8__1_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold379 sb_8__1_.mem_left_track_55.ccff_tail VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_4__A0 sb_8__1_.mux_left_track_45.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_41.mux_l2_in_0_ net336 sb_8__1_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_41.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk net806 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input21_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__269__A sb_8__1_.mux_left_track_53.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net396 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk net703
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold110 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold121 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold143 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold132 cbx_8__1_.mem_top_ipin_13.ccff_tail VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_1.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xhold154 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold176 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold165 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR net531
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold187 sb_8__1_.mem_top_track_2.ccff_tail VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold198 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__A1 sb_8__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_28.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_340_ net40 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2__A1 net72 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_271_ sb_8__1_.mux_left_track_49.out VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input69_A chany_top_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net230
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output225_A net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_1_ net39 cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput204 net204 VGND VGND VPWR VPWR chany_top_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput226 net226 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_3__364 VGND VGND VPWR VPWR net364 cbx_8__1_.mux_top_ipin_14.mux_l2_in_3__364/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ net746 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_11_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_2_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__301
+ VGND VGND VPWR VPWR net301 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__301/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk net753 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_19_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_0.mux_l2_in_3__347 VGND VGND VPWR VPWR net347 sb_8__1_.mux_top_track_0.mux_l2_in_3__347/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_26_prog_clk net596 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_2__S sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_323_ sb_8__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_5.mux_l3_in_0_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_77_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_0__S sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net267 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_2_ net56 cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_3__236 VGND VGND VPWR VPWR net236 cbx_8__1_.mux_top_ipin_5.mux_l2_in_3__236/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk net733
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ net402 VGND VGND VPWR
+ VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_24_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net296 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_2_ net27 sb_8__1_.mux_left_track_35.out cbx_8__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk net836
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_8__1_.mux_top_track_44.mux_l2_in_0_ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_44_prog_clk net552 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__277__A sb_8__1_.mux_left_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_306_ net66 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk net734 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__285
+ VGND VGND VPWR VPWR net285 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__285/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net379 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold14 test_enable VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold47 chany_top_in_0[7] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold25 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X VGND VGND
+ VPWR VPWR net402 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold58 cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR VPWR net424
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__1_.mux_top_track_2.mux_l1_in_0__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold69 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_1_ net217 net214 sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_hold500_A sb_8__1_.mem_top_track_12.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk net863
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_33.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_0__S sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3_ net70 net39 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_30_prog_clk net658 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_21_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold506 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net872
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold517 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net883
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net815 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_44.mux_l1_in_1_ net23 net38 sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_0__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk net661
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput104 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_39_prog_clk net535 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input99_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__290__A sb_8__1_.mux_left_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_left_track_51.mux_l1_in_1__A1 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold303 cbx_8__1_.mem_top_ipin_8.ccff_tail VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold314 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold325 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold369 sb_8__1_.mem_left_track_49.ccff_tail VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold347 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold358 cby_8__1_.cby_8__8_.mem_right_ipin_14.ccff_tail VGND VGND VPWR VPWR net724
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ net812 net232 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold336 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_0__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_4__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_83_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input14_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__285__A sb_8__1_.mux_left_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l1_in_1__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net263 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__mux2_8
XFILLER_67_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_3__S sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_2_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_1.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xhold111 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold144 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold133 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold122 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_3_ net312 net4 sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xhold155 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold177 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_1__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold166 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold199 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold188 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input6_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk net474
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_270_ sb_8__1_.mux_left_track_51.out VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_2__A0 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output218_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.out cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_9_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ net601 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__299
+ VGND VGND VPWR VPWR net299 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__299/LO
+ sky130_fd_sc_hd__conb_1
Xoutput205 net205 VGND VGND VPWR VPWR chany_top_out_0[7] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput216 net216 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_1_prog_clk net855
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput227 net227 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
XFILLER_95_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l2_in_3__A1 sb_8__1_.mux_left_track_57.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_41.mux_l1_in_0_ net227 net64 sb_8__1_.mem_left_track_41.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk net763 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3__A0 net73 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_26_prog_clk net500 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l1_in_0__A0 sb_8__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2__A0 net74 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_2__A0 sb_8__1_.mux_left_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ sb_8__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
Xsb_8__1_.mux_left_track_53.mux_l2_in_0_ net342 sb_8__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_53.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input81_A chany_top_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_3__S sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__297
+ VGND VGND VPWR VPWR net297 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__297/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__S
+ net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_1_ net7 cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_12_prog_clk net802
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_1_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_43_prog_clk net677 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__293__A sb_8__1_.mux_left_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_305_ net65 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk net577 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_2__A0 sb_8__1_.mux_left_track_15.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_11_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_4__A0 sb_8__1_.mux_left_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_21.mux_l3_in_0_ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_6_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_47.mux_l1_in_0__A0 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_2__A0 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l1_in_0__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_50_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold15 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold26 chanx_left_in[13] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold37 cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold59 cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND
+ VPWR VPWR net425 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_68_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold48 net91 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_0_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk net515
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_33.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input44_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__288__A sb_8__1_.mux_left_track_15.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_30_prog_clk net591 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2_ net77 net46 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold518 cbx_8__1_.mem_top_ipin_15.mem_out\[2\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold507 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[2\] VGND VGND VPWR VPWR net873
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net409 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_11.mux_l1_in_2_ sb_8__1_.mux_left_track_23.out net13 cbx_8__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_80_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_44.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ net105 sb_8__1_.mem_top_track_44.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_2__S cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput105 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_42_prog_clk net496 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_21.mux_l2_in_1_ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_left_track_11.mux_l2_in_1__321 VGND VGND VPWR VPWR net321 sb_8__1_.mux_left_track_11.mux_l2_in_1__321/LO
+ sky130_fd_sc_hd__conb_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_0__S sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold326 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold315 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold304 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold348 sb_8__1_.mem_left_track_55.mem_out\[0\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold359 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold337 cbx_8__1_.mem_top_ipin_0.ccff_tail VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk
+ net724 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xcbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_1_prog_clk net869
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_5.mux_l1_in_1_ net219 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_0__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk net758 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l1_in_1__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_31.mux_l1_in_1__332 VGND VGND VPWR VPWR net332 sb_8__1_.mux_left_track_31.mux_l1_in_1__332/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold101 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold123 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold134 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold112 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_2_ net6 net18 sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xhold156 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_1__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold145 cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_tail VGND VGND VPWR VPWR net511
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold167 sb_8__1_.mem_bottom_track_5.ccff_tail VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold178 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold189 cbx_8__1_.mem_top_ipin_7.ccff_tail VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_2__A1 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__296__A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__242 VGND VGND VPWR VPWR net242 cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__242/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_2__S sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput206 net206 VGND VGND VPWR VPWR chany_top_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput217 net217 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_10.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xoutput228 net228 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold15_A top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_1__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_25_prog_clk net477 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2__A1 net43 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input109_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_321_ net82 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input74_A chany_top_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_55.mux_l1_in_0__A0 net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l1_in_0__A0 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net233 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net285 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk net785 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.out cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__ebufn_8
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_0_ net446 cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ cbx_8__1_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_43_prog_clk net797 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_304_ net93 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_4__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_7_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3_ net245 net86 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_1__S sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold82_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk net710 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_11.mux_l3_in_0_ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xhold16 net111 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_8__1_.mux_left_track_53.mux_l1_in_0_ net225 net80 sb_8__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xhold38 chany_bottom_in[12] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold27 net8 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold49 cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X VGND VGND
+ VPWR VPWR net415 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_13.mux_l1_in_0__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_30_prog_clk net594 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_43_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
+ net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold508 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net874
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold519 sb_8__1_.mem_top_track_44.mem_out\[1\] VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_11.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net445 cbx_8__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput106 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net106 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_41_prog_clk net602 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l2_in_3__A1 sb_8__1_.mux_left_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_21.mux_l2_in_0_ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4_ sb_8__1_.mux_bottom_track_45.out
+ net61 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net277 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__299__A sb_8__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l1_in_0__A0 sb_8__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ net417 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_11.mux_l2_in_1_ net321 net226 sb_8__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold316 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold305 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold327 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold338 cbx_8__1_.mem_top_ipin_7.mem_out\[2\] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold349 sb_8__1_.mem_bottom_track_1.ccff_head VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__clkdlybuf4s25_1
Xload_slew230 net99 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_16
Xcbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_13.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_5.mux_l1_in_0_ net91 net78 sb_8__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_31.out sky130_fd_sc_hd__clkbuf_1
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk net722 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_1__A0 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold135 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold124 sb_8__1_.mem_left_track_1.ccff_tail VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_1_ net213 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xhold113 sb_8__1_.mem_left_track_25.ccff_tail VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold102 sb_8__1_.mem_left_track_5.ccff_tail VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold146 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold168 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold157 cby_8__1_.cby_8__8_.ccff_tail VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold179 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_47.mux_l2_in_0__338 VGND VGND VPWR VPWR net338 sb_8__1_.mux_left_track_47.mux_l2_in_0__338/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_0__A0 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3_ net256 net90 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_30_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_25.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_25.out sky130_fd_sc_hd__clkbuf_2
Xoutput207 net207 VGND VGND VPWR VPWR chany_top_out_0[9] sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput218 net218 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0__S cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_1__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__288
+ VGND VGND VPWR VPWR net288 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__288/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_26_prog_clk net614 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_320_ sb_8__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk net799
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_51.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input67_A chany_top_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output223_A net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_52.mux_l2_in_1__356 VGND VGND VPWR VPWR net356 sb_8__1_.mux_top_track_52.mux_l2_in_1__356/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net390 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk net543 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_21.mux_l1_in_0__A0 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_0__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.out sky130_fd_sc_hd__clkbuf_2
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_bottom_track_45.mux_l2_in_1__316 VGND VGND VPWR VPWR net316 sb_8__1_.mux_bottom_track_45.mux_l2_in_1__316/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_46_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l1_in_0__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_303_ sb_8__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_2_ net45 cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_0__A0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk net643 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xhold17 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in VGND VGND
+ VPWR VPWR net383 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold28 cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X VGND VGND VPWR VPWR net394
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold39 net37 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_13.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_30_prog_clk net633 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ net425 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_74_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_left_track_1.mux_l3_in_0_ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2__A0 net77 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold509 sb_8__1_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_11.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput107 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net107 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_41_prog_clk net670 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3_ net69 net38 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_1__A0 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__245 VGND VGND VPWR VPWR net245
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__245/LO sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_11.mux_l2_in_0_ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3__S cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold317 cbx_8__1_.mem_top_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold306 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold339 sb_8__1_.mem_left_track_47.mem_out\[0\] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold328 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk net831
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__A0 net66 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold38_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xload_slew231 net232 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_23.mux_l3_in_0_ sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_23.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l1_in_1__A0 sb_8__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_1__A0 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_1.mux_l2_in_1_ net320 sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input97_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_1__S sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold8_A top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_79_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_1__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold114 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold125 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold103 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_0_ net86 net72 sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xhold158 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold136 sb_8__1_.mem_bottom_track_11.ccff_head VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold147 sb_8__1_.mem_bottom_track_1.ccff_tail VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold169 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_11.mux_l2_in_1__A1 net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_53.out sky130_fd_sc_hd__buf_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net300 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__mux2_4
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_3_ net366 sb_8__1_.mux_left_track_53.out cbx_8__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_0__A1 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2_ net399 net70 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_11.mux_l1_in_1_ net223 net43 sb_8__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input12_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk net612
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xoutput208 net208 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xoutput219 net219 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_bottom_track_45.mux_l3_in_0_ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_23.mux_l2_in_1_ net327 net226 sb_8__1_.mem_left_track_23.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2__A0 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_1.mux_l1_in_2_ net227 net224 sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net379 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_86_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk net635 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk net735
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_51.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__256 VGND VGND VPWR VPWR net256
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__256/LO sky130_fd_sc_hd__conb_1
XFILLER_89_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output216_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net303 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__271
+ VGND VGND VPWR VPWR net271 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__271/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold20_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_47.out sky130_fd_sc_hd__clkbuf_1
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_2__S sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_4_ sb_8__1_.mux_left_track_41.out net33 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_21.mux_l1_in_0__A1 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_0__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_302_ net91 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_45.mux_l2_in_1_ net316 net32 sb_8__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__A1 net86 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net266 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_2.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xhold18 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold29 cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X VGND VGND VPWR VPWR net395
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net274 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_1__A0 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_0_prog_clk
+ net874 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_30_prog_clk net626 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_55_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_52_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk net782
+ net232 VGND VGND VPWR VPWR cbx_8__1_.ccff_head sky130_fd_sc_hd__dfrtp_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_2__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_3_ net238 sb_8__1_.mux_left_track_45.out cbx_8__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xinput108 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net108 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_41_prog_clk net665 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_10_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2_ sb_8__1_.mux_bottom_track_21.out
+ net44 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input42_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_2.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_46_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__267
+ VGND VGND VPWR VPWR net267 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__267/LO
+ sky130_fd_sc_hd__conb_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold307 cby_8__1_.cby_8__8_.mem_right_ipin_5.ccff_tail VGND VGND VPWR VPWR net673
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold318 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold329 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_load_slew232_A net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk net529
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xload_slew232 net233 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__buf_12
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_1__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 chany_top_in_0[6] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_1__A1 net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_1.mux_l2_in_0_ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_41_prog_clk net768 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 sb_8__1_.mem_left_track_45.mem_out\[0\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold104 sb_8__1_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold126 sb_8__1_.mem_bottom_track_53.mem_out\[1\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold159 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold137 sb_8__1_.mem_left_track_17.mem_out\[0\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold148 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_2_ net27 cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__266
+ VGND VGND VPWR VPWR net266 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__266/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_1_ net39 cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_11.mux_l1_in_0_ net50 net73 sb_8__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_3__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__A1 net89 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net382 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xoutput209 net209 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_3__362 VGND VGND VPWR VPWR net362 cbx_8__1_.mux_top_ipin_12.mux_l2_in_3__362/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_23.mux_l2_in_0_ net34 sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_23.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2__A1 net66 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_1.mux_l1_in_1_ net221 net52 sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk net546 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ net881 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_3_ net309 net30 sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xhold490 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR net856
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ net800 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_3__234 VGND VGND VPWR VPWR net234 cbx_8__1_.mux_top_ipin_3.mux_l2_in_3__234/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_3_ sb_8__1_.mux_left_track_29.out net10 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l2_in_2__A1 sb_8__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2_ net77 net46 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk net540 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_39_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input107_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_301_ net90 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xsb_8__1_.mux_bottom_track_45.mux_l2_in_0_ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk net538 net233 VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input72_A chany_top_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3_ net249 net86 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk sb_8__1_.mem_left_track_25.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_25.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_18_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_3.mem_out\[2\]
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_left_track_15.mux_l2_in_0__A0 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__302__A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold19 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_1__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk
+ net872 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__279
+ VGND VGND VPWR VPWR net279 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__279/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_30_prog_clk net641 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_1__A0 sb_8__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk net745
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_57.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_1.mux_l4_in_0_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_2_ net31 sb_8__1_.mux_left_track_27.out cbx_8__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput109 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR
+ VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_41_prog_clk net748 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_45.mux_l1_in_1_ net14 net216 sb_8__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0__S cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_6_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4_ sb_8__1_.mux_bottom_track_45.out
+ net61 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_2.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold308 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold319 sb_8__1_.mem_bottom_track_13.ccff_tail VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew233 net99 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_16
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_2__A0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_1__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput80 chany_top_in_0[24] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
Xinput91 net413 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
Xcbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_2__S sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_41_prog_clk net680 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ net636 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_7.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_1.mux_l3_in_1_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold105 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold116 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold149 sb_8__1_.mem_left_track_31.ccff_tail VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold138 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail
+ VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold127 sb_8__1_.mem_left_track_27.mem_out\[0\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__310__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_9.mux_l2_in_1__346 VGND VGND VPWR VPWR net346 sb_8__1_.mux_left_track_9.mux_l2_in_1__346/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_1__A0 net212 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net231
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_1__A0 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_91_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_1__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net379 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_1.mux_l1_in_0_ net82 net85 sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_3__309 VGND VGND VPWR VPWR net309 sb_8__1_.mux_bottom_track_1.mux_l2_in_3__309/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net282 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__mux2_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__305__A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_3__A0 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_3__366 VGND VGND VPWR VPWR net366 cbx_8__1_.mux_top_ipin_2.mux_l2_in_3__366/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk
+ net820 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_2_ net12 net24 sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xhold480 sb_8__1_.mem_left_track_3.mem_out\[0\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold491 sb_8__1_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.out sky130_fd_sc_hd__clkbuf_2
XFILLER_54_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_8__1_.mem_bottom_track_11.mem_out\[1\] net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l1_in_0__A0 sb_8__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_23_prog_clk net813
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_2_ sb_8__1_.mux_left_track_17.out net17 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ net453 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3__S cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_300_ net89 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_23.mux_l1_in_0_ net35 net65 sb_8__1_.mem_left_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input65_A chany_top_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output221_A net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_2_ net45 cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk net807
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_25.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_35.mux_l2_in_0_ sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_35.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 ccff_head_0_0 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_71_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net292 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_2__A0 sb_8__1_.mux_left_track_15.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_2__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ net840 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk net549 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_30_prog_clk net471 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_32_prog_clk net480 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net433 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__313__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_1_ net11 cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_41_prog_clk net713 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_45.mux_l1_in_0_ net218 net68 sb_8__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_3_ net362 sb_8__1_.mux_left_track_49.out cbx_8__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net302 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3_ net69 net38 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xoutput190 net190 VGND VGND VPWR VPWR chany_top_out_0[20] sky130_fd_sc_hd__buf_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input28_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_29_prog_clk net659 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_35.mux_l1_in_1_ net334 net224 sb_8__1_.mem_left_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_1__S sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold309 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l2_in_1__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_1__S sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_1__A0 net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_2__A1 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__308__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 chany_top_in_0[15] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
Xinput81 chany_top_in_0[25] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
Xinput92 chany_top_in_0[8] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__A1 net93 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__293
+ VGND VGND VPWR VPWR net293 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__293/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_41_prog_clk net744 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_1.mux_l3_in_0_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_90_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_7.mux_l1_in_2_ sb_8__1_.mux_left_track_15.out net18 cbx_8__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_90_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_4_ sb_8__1_.mux_left_track_37.out net6 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold106 cby_8__1_.cby_8__8_.mem_right_ipin_8.ccff_tail VGND VGND VPWR VPWR net472
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold117 cbx_8__1_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold128 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold139 sb_8__1_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_1__A0 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_1__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_1__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input95_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk net737 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_52.mux_l3_in_0_ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_bottom_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__321__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_3__A1 net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_1_ net215 net212 sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xhold470 cbx_8__1_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold481 sb_8__1_.mem_left_track_9.mem_out\[1\] VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold492 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR net858
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input10_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk
+ sb_8__1_.mem_bottom_track_11.mem_out\[0\] net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_5_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_3__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_8__1_.mem_top_track_4.mem_out\[1\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__316__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input2_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_2__S sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_12.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input58_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_52.mux_l2_in_1_ net356 sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output214_A net214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk net887
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_359_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_2__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk net751 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xinput2 ccff_head_1 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_2__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk
+ net829 net229 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk net719 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_31_prog_clk net499 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_29_prog_clk net613 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_19.mux_l1_in_0__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_2_ net29 cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_52.mux_l1_in_2_ net30 net12 sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2_ sb_8__1_.mux_bottom_track_21.out
+ net44 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput180 net180 VGND VGND VPWR VPWR chany_top_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput191 net191 VGND VGND VPWR VPWR chany_top_out_0[21] sky130_fd_sc_hd__buf_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_29_prog_clk net570 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_left_track_35.mux_l1_in_0_ net56 net86 sb_8__1_.mem_left_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_31.mux_l1_in_1__A1 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_1__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_47.mux_l2_in_0_ net338 sb_8__1_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_47.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__324__A sb_8__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput82 chany_top_in_0[26] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_4
Xinput71 chany_top_in_0[16] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
Xinput60 chany_bottom_in[6] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
Xinput93 chany_top_in_0[9] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_41_prog_clk net767 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ net856 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk net848
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_7.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_73_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_3_ sb_8__1_.mux_left_track_25.out net12 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xhold107 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_load_slew230_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold118 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold129 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_10.mux_l2_in_3_ net348 net4 sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l2_in_3__A1 net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net435 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__A0 net73 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_1__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__319__A sb_8__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_2__A0 sb_8__1_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_10.mux_l2_in_3__348 VGND VGND VPWR VPWR net348 sb_8__1_.mux_top_track_10.mux_l2_in_3__348/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input88_A chany_top_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk net559 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_2__S sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ net810 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_0_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xhold460 cbx_8__1_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold471 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net837
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold493 sb_8__1_.mem_top_track_0.mem_out\[1\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold482 sb_8__1_.mem_left_track_11.mem_out\[1\] VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_2__A0 sb_8__1_.mux_left_track_17.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net264 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__mux2_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_2__A0 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_44_prog_clk
+ net502 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_79_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_23_prog_clk net616
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net233
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l2_in_1__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__332__A net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_12.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_10.mux_l4_in_0_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X sb_8__1_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_52.mux_l2_in_0_ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold290 sb_8__1_.mem_left_track_15.mem_out\[0\] VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_27.mux_l1_in_0__A0 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_3__312 VGND VGND VPWR VPWR net312 sb_8__1_.mux_bottom_track_21.mux_l1_in_3__312/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk net513
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_358_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_4__A0 sb_8__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_289_ sb_8__1_.mux_left_track_13.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk net695 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_68_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 ccff_head_2 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_top_track_4.mux_l2_in_3_ net354 net33 sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_1.mux_l1_in_1_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__327__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_29_prog_clk net478 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_29_prog_clk net598 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input70_A chany_top_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_19.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_10.mux_l3_in_1_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_52.mux_l1_in_1_ net24 net36 sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_0__S sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput170 net170 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chany_top_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chany_top_out_0[22] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk net683
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_46_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_29_prog_clk net597 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_49_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput72 chany_top_in_0[17] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
Xinput50 chany_bottom_in[24] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
Xinput61 chany_bottom_in[7] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
Xinput83 chany_top_in_0[27] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
Xinput94 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XANTENNA__340__A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_41_prog_clk net740 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_top_track_4.mux_l4_in_0_ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X
+ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sb_8__1_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ net809 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__282
+ VGND VGND VPWR VPWR net282 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__282/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input33_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk
+ net845 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__1_.mem_left_track_11.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_7.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold108 sb_8__1_.mem_top_track_20.ccff_tail VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_2_ sb_8__1_.mux_left_track_13.out net19 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold119 cbx_8__1_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_10.mux_l2_in_2_ net6 net18 sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_1__S sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_45.mux_l2_in_0__337 VGND VGND VPWR VPWR net337 sb_8__1_.mux_left_track_45.mux_l2_in_0__337/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__335__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_0__S sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net283 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk net537 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_47.mux_l1_in_0_ net222 net67 sb_8__1_.mem_left_track_47.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_17.mux_l2_in_1__A1 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__289
+ VGND VGND VPWR VPWR net289 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__289/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_4.mux_l3_in_1_ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xhold461 sb_8__1_.mem_top_track_0.mem_out\[0\] VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold450 sb_8__1_.mem_left_track_21.mem_out\[0\] VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold472 cbx_8__1_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold483 cbx_8__1_.mem_top_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold494 cbx_8__1_.mem_top_ipin_4.mem_out\[2\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_35.mux_l1_in_0__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__254 VGND VGND VPWR VPWR net254
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__254/LO sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_10.mux_l1_in_3_ net59 net44 sb_8__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_2__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2__A1 net66 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk net553
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_17.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk net505
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net293 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__mux2_4
Xhold280 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold291 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l2_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_left_track_27.mux_l1_in_0__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk net839
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
X_357_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_5.mux_l1_in_0__A0 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_4__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_288_ sb_8__1_.mux_left_track_15.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR_A
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_4.mux_l2_in_2_ net16 net61 sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 chanx_left_in[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_bottom_track_1.mux_l1_in_0_ net65 net82 sb_8__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk net731
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_49.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA__343__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__A1 net429 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk net563 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l2_in_3__A1 sb_8__1_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_29_prog_clk net460 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold512_A cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input63_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_0__A0 sb_8__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk
+ net536 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_2__A0 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_52_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__338__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_10.mux_l3_in_0_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_52.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ net106 sb_8__1_.mem_top_track_52.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_3__S sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput160 net160 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net99 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput182 net182 VGND VGND VPWR VPWR chany_top_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR chany_top_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l2_in_3__A1 sb_8__1_.mux_left_track_49.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_15_prog_clk cbx_8__1_.mem_top_ipin_0.mem_out\[1\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_29_prog_clk net508 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3_ net246 net75 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net379 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2__A0 net79 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_2__A0 sb_8__1_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold71_A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput40 chany_bottom_in[15] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_4
Xinput73 chany_top_in_0[18] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_4
Xinput51 chany_bottom_in[25] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
Xinput62 chany_bottom_in[8] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
Xinput84 net447 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
Xinput95 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.out sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk net521 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ net889 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_41_prog_clk net678 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk
+ net828 net232 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input26_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net465
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold109 sb_8__1_.mem_top_track_0.ccff_tail VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__1_.mux_top_track_10.mux_l2_in_1_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__351__A net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_1__A0 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk net726 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_3__360 VGND VGND VPWR VPWR net360 cbx_8__1_.mux_top_ipin_10.mux_l2_in_3__360/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk net709
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_0__S sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_3__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l4_in_0_ net442 cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_1.ccff_tail VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__275
+ VGND VGND VPWR VPWR net275 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__275/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__346__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_4.mux_l3_in_0_ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold451 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold462 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR net828
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold440 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold495 sb_8__1_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold473 cbx_8__1_.mem_top_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold484 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net850
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_35.mux_l1_in_0__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_2__S sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_10.mux_l1_in_2_ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ sb_8__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input93_A chany_top_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0__A cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net503
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_17.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk net875
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3_ net257 net429 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_29_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold270 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[2\] VGND VGND VPWR VPWR net636
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold281 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold292 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_2__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk net826
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xsb_8__1_.mux_left_track_17.mux_l3_in_0_ sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_17.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_356_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__1_.mux_left_track_5.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_287_ sb_8__1_.mux_left_track_17.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ net441 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_4.mux_l2_in_1_ net48 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__1_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xinput5 net386 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk net771
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_49.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk net684 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__296
+ VGND VGND VPWR VPWR net296 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__296/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_28_prog_clk net569 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk
+ net639 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_1__S sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk net732 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input56_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output212_A net212 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk
+ net531 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk net547 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
X_339_ net39 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__A0 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_2__A1 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4_ sb_8__1_.mux_bottom_track_45.out
+ net61 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_1__A0 sb_8__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__305
+ VGND VGND VPWR VPWR net305 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__305/LO
+ sky130_fd_sc_hd__conb_1
Xoutput161 net161 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput150 net150 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput194 net194 VGND VGND VPWR VPWR chany_top_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_top_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_left_track_17.mux_l2_in_1_ net324 net223 sb_8__1_.mem_left_track_17.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_30_prog_clk net497 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input110_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2_ net34 net65 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_3__239 VGND VGND VPWR VPWR net239 cbx_8__1_.mux_top_ipin_8.mux_l2_in_3__239/LO
+ sky130_fd_sc_hd__conb_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_2__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l4_in_0_ net439 cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_6.ccff_tail VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_12.mux_l1_in_3__349 VGND VGND VPWR VPWR net349 sb_8__1_.mux_top_track_12.mux_l1_in_3__349/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_left_track_51.mux_l1_in_0__A0 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput30 chanx_left_in[6] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_13_prog_clk net843
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xinput41 chany_bottom_in[16] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xinput52 chany_bottom_in[26] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_4
Xinput63 chany_bottom_in[9] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
Xinput85 chany_top_in_0[29] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
Xinput74 chany_top_in_0[19] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net272 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xinput96 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_3__S sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk net756 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_18_prog_clk net655 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_41_prog_clk net662 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ net443 VGND VGND VPWR
+ VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_10.mux_l2_in_0_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net419 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_37.out sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ net438 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[2\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_33_prog_clk net603 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_13_prog_clk net871
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_27.mux_l1_in_1__329 VGND VGND VPWR VPWR net329 sb_8__1_.mux_left_track_27.mux_l1_in_1__329/LO
+ sky130_fd_sc_hd__conb_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_19_prog_clk net487 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold27_A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l2_in_2__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold441 sb_8__1_.mem_left_track_23.ccff_tail VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold463 cby_8__1_.cby_8__8_.mem_right_ipin_0.ccff_tail VGND VGND VPWR VPWR net829
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold430 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold452 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net818
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold485 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR net851
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold496 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[2\] VGND VGND VPWR VPWR net862
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold474 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR net840
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_1__S sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_10.mux_l1_in_1_ net108 net106 sb_8__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__A1 net75 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk net774
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_3_ net234 sb_8__1_.mux_left_track_55.out cbx_8__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_82_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk net762
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_2_ net437 cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__D cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold271 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold260 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net730 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xhold293 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold282 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_8__1_.mem_top_ipin_3.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__267__A sb_8__1_.mux_left_track_57.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
X_355_ sb_8__1_.mux_top_track_0.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_286_ sb_8__1_.mux_left_track_19.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_4.mux_l2_in_0_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xinput6 chanx_left_in[11] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XFILLER_49_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net880 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net275 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__mux2_8
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_7.mux_l3_in_0_ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_left_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_59_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_29_prog_clk net623 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_45_prog_clk
+ net890 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk net557 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input49_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ net38 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk net696 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
X_269_ sb_8__1_.mux_left_track_53.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__A1 net63 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3_ net69 net38 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput151 net151 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput140 net140 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chany_top_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chany_top_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput173 net173 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
XFILLER_87_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_17.mux_l2_in_0_ net37 sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_17.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk net668
+ net231 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_29_prog_clk net572 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_1_ net63 cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net379 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input103_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l1_in_1__A0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_57.mux_l2_in_0__344 VGND VGND VPWR VPWR net344 sb_8__1_.mux_left_track_57.mux_l2_in_0__344/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_0__S sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_3.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_78_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_7.mux_l2_in_1_ net345 sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.out sky130_fd_sc_hd__buf_4
Xinput31 chanx_left_in[7] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xinput20 net444 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
Xinput64 chany_top_in_0[0] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_13_prog_clk cbx_8__1_.mem_top_ipin_9.mem_out\[1\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xinput53 chany_bottom_in[27] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
Xinput42 chany_bottom_in[17] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xinput86 net428 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xinput75 chany_top_in_0[1] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_4
Xinput97 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_18_prog_clk net630 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_41_prog_clk net488 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_3__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_40_prog_clk
+ net1 net233 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_87_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__A1 sb_8__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__275__A sb_8__1_.mux_left_track_41.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l1_in_0__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_3_ net239 sb_8__1_.mux_left_track_53.out cbx_8__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net231
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__304
+ VGND VGND VPWR VPWR net304 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__304/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_7.mux_l2_in_1__345 VGND VGND VPWR VPWR net345 sb_8__1_.mux_left_track_7.mux_l2_in_1__345/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2_ net74 net43 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_48_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_3.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_21_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_29.mux_l1_in_1__A1 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_7.mux_l1_in_2_ net227 net224 sb_8__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input31_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_1__A0 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_33_prog_clk net660 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output118_A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_53.mux_l3_in_0_ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_bottom_track_53.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk net725 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold420 sb_8__1_.mem_left_track_45.ccff_tail VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold442 sb_8__1_.mem_left_track_37.mem_out\[0\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold431 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold453 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net819
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold475 sb_8__1_.mem_top_track_52.mem_out\[0\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold486 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR net852
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xclkbuf_leaf_3_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold464 cbx_8__1_.mem_top_ipin_14.ccff_tail VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold497 sb_8__1_.mem_left_track_33.mem_out\[0\] VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__264
+ VGND VGND VPWR VPWR net264 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__264/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_10.mux_l1_in_0_ net104 net110 sb_8__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_1__A0 sb_8__1_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input79_A chany_top_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_4_ sb_8__1_.mux_left_track_41.out net33 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_2_ net26 sb_8__1_.mux_left_track_37.out cbx_8__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold261 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold250 sb_8__1_.mem_top_track_4.mem_out\[0\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net539 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold272 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold283 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_49_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold294 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_8.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk net516
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_bottom_track_53.mux_l2_in_1_ net318 sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_bottom_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_354_ sb_8__1_.mux_top_track_2.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_285_ sb_8__1_.mux_left_track_21.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 chanx_left_in[12] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__308
+ VGND VGND VPWR VPWR net308 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__308/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_1__S sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_29_prog_clk net587 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_44_prog_clk
+ net878 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk sb_8__1_.mem_top_track_10.mem_out\[2\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ net766 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ sb_8__1_.mux_top_track_36.out VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_268_ sb_8__1_.mux_left_track_55.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2_ sb_8__1_.mux_bottom_track_21.out
+ net44 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk net672 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_8.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xoutput130 net130 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput152 net152 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_top_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chany_top_out_0[26] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_bottom_track_53.mux_l1_in_2_ net31 net13 sb_8__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2__A0 net399 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_29_prog_clk net491 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l2_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_0.mux_l1_in_1__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_4.mux_l1_in_0_ net106 net103 sb_8__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3_ net250 net414 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input61_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xload_slew229 net230 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_12
XFILLER_78_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_1__S sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.out sky130_fd_sc_hd__buf_4
XFILLER_93_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_7.mux_l2_in_0_ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 chanx_left_in[15] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput21 chanx_left_in[25] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
Xcbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_13_prog_clk cbx_8__1_.mem_top_ipin_9.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xinput32 chanx_left_in[8] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput54 chany_bottom_in[28] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
Xinput43 chany_bottom_in[18] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput76 chany_top_in_0[20] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xinput87 chany_top_in_0[3] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xinput65 chany_top_in_0[10] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
Xinput98 isol_n VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_18_prog_clk net625 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net511 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_38_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_37.mux_l1_in_1__A1 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net642 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net273 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA__291__A sb_8__1_.mux_left_track_9.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_2_ net27 cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk net835
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_35.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_15_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_3_ net310 net26 sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_17.mux_l1_in_0_ net39 net69 sb_8__1_.mem_left_track_17.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk net492
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_53.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_3.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net308 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ net115 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_29.mux_l2_in_0_ sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_88_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_1__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_7.mux_l1_in_1_ net221 net47 sb_8__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input24_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_33_prog_clk net644 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk net578
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_31.mux_l2_in_0_ sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_31.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_3_ net319 net27 sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_50_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l4_in_0_ net415 cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.ccff_tail VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xhold410 sb_8__1_.mem_left_track_31.mem_out\[0\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold421 cby_8__1_.cby_8__8_.mem_right_ipin_7.ccff_tail VGND VGND VPWR VPWR net787
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold454 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR net820
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold432 cby_8__1_.cby_8__8_.mem_right_ipin_4.ccff_tail VGND VGND VPWR VPWR net798
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold443 cby_8__1_.cby_8__8_.mem_right_ipin_6.ccff_tail VGND VGND VPWR VPWR net809
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold476 cbx_8__1_.mem_top_ipin_12.mem_out\[2\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold487 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[2\] VGND VGND VPWR VPWR net853
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold465 cbx_8__1_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold498 sb_8__1_.mem_top_track_20.mem_out\[1\] VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_0__S cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_3_ sb_8__1_.mux_left_track_29.out net10 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_output228_A net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.out sky130_fd_sc_hd__clkbuf_2
XFILLER_48_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3_ net241 net90 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold32_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_1_ net6 cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_2__A0 sb_8__1_.mux_left_track_17.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_left_track_29.mux_l1_in_1_ net330 net221 sb_8__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_82_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold240 sb_8__1_.mem_top_track_44.ccff_tail VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold262 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold251 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold284 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold273 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[2\] VGND VGND VPWR VPWR net639
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold295 cbx_8__1_.mem_top_ipin_3.ccff_tail VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_11.mux_l4_in_0_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X sb_8__1_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_53.mux_l2_in_0_ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_353_ sb_8__1_.mux_top_track_4.out VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_284_ sb_8__1_.mux_left_track_23.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_31.mux_l1_in_1_ net332 net222 sb_8__1_.mem_left_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_3__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput8 net392 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_4__A0 sb_8__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net652 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk net842
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_11_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_8__1_.mem_top_track_10.mem_out\[1\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4_ sb_8__1_.mux_bottom_track_37.out
+ net36 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l4_in_0_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X sb_8__1_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_61_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__294__A sb_8__1_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_336_ net36 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_267_ sb_8__1_.mux_left_track_57.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
Xcbx_8__1_.mux_top_ipin_3.mux_l1_in_2_ sb_8__1_.mux_left_track_19.out net16 cbx_8__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_0__S sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk net691 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_19.mux_l2_in_1__325 VGND VGND VPWR VPWR net325 sb_8__1_.mux_left_track_19.mux_l2_in_1__325/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_64_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_8.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__A1 net86 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput131 net131 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chany_top_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_bottom_track_11.mux_l3_in_1_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xoutput197 net197 VGND VGND VPWR VPWR chany_top_out_0[27] sky130_fd_sc_hd__buf_12
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_53.mux_l1_in_1_ net25 net217 sb_8__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2__A1 net70 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_32_prog_clk net628 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_left_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2_ net60 net68 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input54_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__289__A sb_8__1_.mux_left_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_11.mux_l1_in_1__A0 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_319_ sb_8__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_left_in[16] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 chanx_left_in[26] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XFILLER_52_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk net669
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xinput33 chanx_left_in[9] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
Xinput55 chany_bottom_in[29] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput44 chany_bottom_in[19] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
Xinput77 chany_top_in_0[21] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
Xinput66 chany_top_in_0[11] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
Xinput88 chany_top_in_0[4] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput99 prog_reset VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_18_prog_clk net455 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk net886
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_3__S cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net757 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_7.mux_l3_in_1_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_1__S sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_74_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk net761
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_35.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_2_ net8 net20 sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_3_ net363 sb_8__1_.mux_left_track_57.out cbx_8__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_hold62_A chany_top_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__1_.mem_bottom_track_53.mem_out\[0\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_5.mux_l2_in_1__340 VGND VGND VPWR VPWR net340 sb_8__1_.mux_left_track_5.mux_l2_in_1__340/LO
+ sky130_fd_sc_hd__conb_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_7.mux_l1_in_0_ net53 net77 sb_8__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_33_prog_clk net473 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_6.mux_l2_in_3__357 VGND VGND VPWR VPWR net357 sb_8__1_.mux_top_track_6.mux_l2_in_3__357/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_2_ net9 net21 sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3__A0 net69 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold400 cby_8__1_.cby_8__8_.mem_left_ipin_2.ccff_tail VGND VGND VPWR VPWR net766
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold411 cbx_8__1_.mem_top_ipin_4.ccff_tail VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold433 sb_8__1_.mem_left_track_51.mem_out\[0\] VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold422 cby_8__1_.cby_8__8_.mem_right_ipin_12.ccff_tail VGND VGND VPWR VPWR net788
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold444 cby_8__1_.cby_8__8_.mem_right_ipin_3.ccff_tail VGND VGND VPWR VPWR net810
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold477 cbx_8__1_.mem_top_ipin_9.mem_out\[2\] VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold455 sb_8__1_.mem_left_track_23.mem_out\[0\] VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold466 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR net832
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold488 cbx_8__1_.mem_top_ipin_8.mem_out\[2\] VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold499 sb_8__1_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_13_prog_clk net884
+ net229 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_2_ sb_8__1_.mux_left_track_17.out net17 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_11.mux_l1_in_3_ net217 net215 sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__297__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_2_ net59 cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_3__S sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__252 VGND VGND VPWR VPWR net252
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__252/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_11_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_94_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_29.mux_l1_in_0_ net60 net90 sb_8__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_54_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold230 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold241 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold252 sb_8__1_.mem_bottom_track_5.mem_out\[2\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold296 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold263 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold274 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold285 sb_8__1_.mem_bottom_track_1.mem_out\[0\] VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_23.mux_l2_in_1__327 VGND VGND VPWR VPWR net327 sb_8__1_.mux_left_track_23.mux_l2_in_1__327/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_352_ sb_8__1_.mux_top_track_6.out VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mux_top_ipin_13.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ net389 cbx_8__1_.mem_top_ipin_13.ccff_tail VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
X_283_ sb_8__1_.mux_left_track_25.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xsb_8__1_.mux_left_track_31.mux_l1_in_0_ net59 net89 sb_8__1_.mem_left_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l1_in_3_ net216 net214 sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_2__A0 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xinput9 net420 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_18_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_4__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk cbx_8__1_.mem_top_ipin_12.mem_out\[1\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_2__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_8__1_.mem_top_track_10.mem_out\[0\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3_ net73 net42 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_335_ net35 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
X_266_ net84 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l1_in_1__A0 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_3.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_2__S sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_1__A0 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput132 net132 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput143 net143 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__259 VGND VGND VPWR VPWR net259
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__259/LO sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_bottom_track_11.mux_l3_in_0_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xoutput198 net198 VGND VGND VPWR VPWR chany_top_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chany_top_out_0[18] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_bottom_track_53.mux_l1_in_0_ net219 net66 sb_8__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_13.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk net620 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_1_ net405 cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_2__A0 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input47_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_11.mux_l1_in_1__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_318_ net79 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[17] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput34 net440 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 net436 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
Xinput23 chanx_left_in[27] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
Xinput67 chany_top_in_0[12] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
Xinput78 chany_top_in_0[22] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
Xinput89 chany_top_in_0[5] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput56 chany_bottom_in[2] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__249 VGND VGND VPWR VPWR net249
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__249/LO sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l2_in_3__A1 sb_8__1_.mux_left_track_49.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3__A0 net72 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_25_prog_clk net581 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l3_in_0_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l1_in_0__A0 sb_8__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2__A0 net72 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net291 net411 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_0__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_74_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_1_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_2_ net15 net226 cbx_8__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold55_A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net486
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2_ net78 net47 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_32_prog_clk net599 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_2__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_4__A0 sb_8__1_.mux_left_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_49.mux_l1_in_0__A0 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk net494 net231 VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net262 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1 net369 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_15_prog_clk net522 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_1__A0 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_1_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_0.mux_l2_in_3_ net347 net31 sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_30_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold401 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_8__1_.mux_top_track_4.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold412 sb_8__1_.mem_left_track_9.mem_out\[0\] VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold434 sb_8__1_.mem_bottom_track_11.mem_out\[2\] VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold423 sb_8__1_.mem_left_track_11.ccff_tail VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold445 cbx_8__1_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold478 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR net844
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold456 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR net822
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold467 sb_8__1_.mem_left_track_19.mem_out\[0\] VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold489 cbx_8__1_.mem_top_ipin_10.mem_out\[2\] VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_13_prog_clk cbx_8__1_.mem_top_ipin_15.mem_out\[1\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_bottom_track_11.mux_l1_in_2_ net213 net219 sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_3__240 VGND VGND VPWR VPWR net240 cbx_8__1_.mux_top_ipin_9.mux_l2_in_3__240/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1__S cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_47_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l2_in_1__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold220 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold253 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold231 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold242 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold264 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold275 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold286 cby_8__1_.cby_8__8_.mem_right_ipin_13.ccff_tail VGND VGND VPWR VPWR net652
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold297 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_351_ net52 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net379 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_282_ sb_8__1_.mux_left_track_27.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input77_A chany_top_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_7.mux_l1_in_2_ net212 net218 sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net289 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_43_prog_clk net791 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_21.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_3_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_13_prog_clk net877
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk net550
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_3__365 VGND VGND VPWR VPWR net365 cbx_8__1_.mux_top_ipin_15.mux_l2_in_3__365/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_46_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_0.mux_l4_in_0_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ net63 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l1_in_1__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_3.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk net755
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_53.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_1__A1 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk net524 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xoutput133 net133 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput177 net177 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chany_top_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chany_top_out_0[19] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk net707 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_13.mux_l3_in_0_ net388 cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mem_top_ipin_13.mem_out\[2\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk net523 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_2__A1 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_3__237 VGND VGND VPWR VPWR net237 cbx_8__1_.mux_top_ipin_6.mux_l2_in_3__237/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_78_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_317_ net78 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
Xinput13 chanx_left_in[18] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
Xinput35 chany_bottom_in[10] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xinput46 chany_bottom_in[20] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput24 chanx_left_in[28] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
Xinput68 chany_top_in_0[13] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_4
Xinput79 chany_top_in_0[23] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput57 net450 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk net519 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ net685 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_25_prog_clk net580 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_55.mux_l2_in_0_ net343 sb_8__1_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_55.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_0__S sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__283
+ VGND VGND VPWR VPWR net283 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__283/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_3__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_0.mux_l3_in_1_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_57.mux_l1_in_0__A0 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_0_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4__S cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_1_ net387 cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail net98 VGND
+ VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XANTENNA_hold48_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_32_prog_clk net469 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_2__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_4__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_2__S sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_37_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 net371 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__buf_8
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_14_prog_clk net637 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_0_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_62_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_0.mux_l2_in_2_ net13 net25 sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xhold402 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold435 sb_8__1_.mem_top_track_0.mem_out\[2\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold413 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold424 cby_8__1_.cby_8__8_.mem_right_ipin_1.ccff_tail VGND VGND VPWR VPWR net790
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold457 sb_8__1_.mem_left_track_21.ccff_tail VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold468 sb_8__1_.mem_bottom_track_45.mem_out\[1\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold446 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR net812
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold479 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net845
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_3__358 VGND VGND VPWR VPWR net358 cbx_8__1_.mux_top_ipin_0.mux_l2_in_3__358/LO
+ sky130_fd_sc_hd__conb_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_15.mux_l1_in_0__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_13_prog_clk cbx_8__1_.mem_top_ipin_15.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_11.mux_l1_in_1_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ left_width_0_height_0_subtile_1__pin_inpad_0_ sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_48_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input22_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_13.mux_l1_in_2_ sb_8__1_.mux_left_track_27.out net11 cbx_8__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_5_prog_clk
+ net850 net229 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_90_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__A1 sb_8__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold210 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l2_in_3__A1 sb_8__1_.mux_left_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold221 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold232 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold243 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold254 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold287 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold276 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold265 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold298 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net466 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_350_ sb_8__1_.mux_top_track_10.out VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_281_ sb_8__1_.mux_left_track_29.out VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net111 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_7.mux_l1_in_1_ left_width_0_height_0_subtile_2__pin_inpad_0_
+ left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_43_prog_clk net671 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output226_A net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk net548 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net816
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_3__S sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk net718
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l2_in_3__A1 sb_8__1_.mux_left_track_51.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ sb_8__1_.mux_top_track_44.out VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l2_in_1__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__278
+ VGND VGND VPWR VPWR net278 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__278/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_41_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_0__A0 sb_8__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l1_in_2__A0 sb_8__1_.mux_left_track_23.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk net772
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold78_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk net675 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xoutput134 net134 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput167 net167 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chany_top_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput189 net189 VGND VGND VPWR VPWR chany_top_out_0[1] sky130_fd_sc_hd__buf_12
XFILLER_87_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net817 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net294 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__mux2_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_316_ net77 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chany_bottom_in[11] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_4
Xinput14 chanx_left_in[19] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput25 chanx_left_in[29] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xinput69 chany_top_in_0[14] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
Xinput47 chany_bottom_in[21] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xinput58 chany_bottom_in[4] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk net698 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_25_prog_clk net562 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_1__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_0.mux_l3_in_0_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2__A0 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_57.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l2_in_1__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input52_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk
+ net571 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__300__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_23.mux_l1_in_0__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_3__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_0__A0 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3_ net253 net90 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_0__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_31_prog_clk net520 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net427 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ net385 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_13.mux_l3_in_0_ sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_55.mux_l1_in_0_ net226 net81 sb_8__1_.mem_left_track_55.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3 reset VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_94_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_14_prog_clk net579 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net280 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_25.mux_l1_in_1__328 VGND VGND VPWR VPWR net328 sb_8__1_.mux_left_track_25.mux_l1_in_1__328/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_0.mux_l2_in_1_ net35 net52 sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_90_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold436 cbx_8__1_.mem_top_ipin_6.ccff_tail VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold403 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold425 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold414 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net780
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold447 sb_8__1_.mem_top_track_4.mem_out\[2\] VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold469 sb_8__1_.mem_left_track_35.mem_out\[0\] VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold458 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net278 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_15.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__290
+ VGND VGND VPWR VPWR net290 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__290/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk net514 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk net830
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_2__A0 net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail net98 VGND
+ VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
Xsb_8__1_.mux_bottom_track_11.mux_l1_in_0_ net89 net74 sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_13.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input15_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk
+ net729 net229 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ net432 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4_ sb_8__1_.mux_bottom_track_37.out
+ net36 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net379 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk net801
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xhold200 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold211 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold244 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold233 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold222 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold266 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold277 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold255 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold299 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold288 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input7_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk net681 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l2_in_1__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_13.mux_l2_in_1_ net322 net221 sb_8__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_280_ sb_8__1_.mux_left_track_31.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_0__S sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_7.mux_l1_in_0_ net90 net77 sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_43_prog_clk net674 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk net824 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output219_A net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4__A0 net93 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l4_in_0_ net401 cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_2.ccff_tail VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk net804
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_44.mux_l2_in_1__355 VGND VGND VPWR VPWR net355 sb_8__1_.mux_top_track_44.mux_l2_in_1__355/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_1__A0 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__243 VGND VGND VPWR VPWR net243 cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__243/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_33.out sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ net61 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_bottom_track_37.mux_l2_in_1__315 VGND VGND VPWR VPWR net315 sb_8__1_.mux_bottom_track_37.mux_l2_in_1__315/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input82_A chany_top_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 net377 net368 net373 net379 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_50_prog_clk
+ net773 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput124 net124 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3_ net258 sb_8__1_.mux_bottom_track_53.out
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput135 net135 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
XANTENNA__303__A sb_8__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput157 net157 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput179 net179 VGND VGND VPWR VPWR chany_top_out_0[10] sky130_fd_sc_hd__buf_12
XFILLER_87_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_13.mux_l2_in_1__A1 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_55.mux_l2_in_0__343 VGND VGND VPWR VPWR net343 sb_8__1_.mux_left_track_55.mux_l2_in_0__343/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ net400 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_315_ sb_8__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput26 chanx_left_in[2] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_left_in[1] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput37 net404 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput48 chany_bottom_in[22] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
Xinput59 net398 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
XANTENNA_sb_8__1_.mux_left_track_31.mux_l1_in_0__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk net796 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_27.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_27.out sky130_fd_sc_hd__clkbuf_2
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_0__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4__A1 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_1__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2__A1 net70 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk net493
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_27.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_45_prog_clk net618
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1__S cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk net834
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk net728 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_left_track_23.mux_l1_in_0__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l2_in_2__A0 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_0__A0 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_2_ net399 cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_32_prog_clk net586 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_3__S sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ net407 cby_8__1_.cby_8__8_.mem_right_ipin_7.ccff_tail VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 net367 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_14_prog_clk net663 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_0.mux_l2_in_0_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_4.mux_l2_in_3__354 VGND VGND VPWR VPWR net354 sb_8__1_.mux_top_track_4.mux_l2_in_3__354/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold426 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold415 sb_8__1_.mem_left_track_17.ccff_tail VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold404 sb_8__1_.mem_left_track_13.ccff_tail VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold437 sb_8__1_.mem_top_track_28.mem_out\[1\] VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold459 sb_8__1_.mem_top_track_2.mem_out\[2\] VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold448 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_3.mux_l3_in_0_ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_80_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk net814 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_2__A1 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_13.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_2__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3_ net73 net42 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk net859
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__306__A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold201 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold212 cbx_8__1_.mem_top_ipin_5.ccff_tail VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold223 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold234 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold245 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold267 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[2\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
Xhold256 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xhold278 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold289 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_13.mux_l2_in_0_ net42 sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_0.mux_l1_in_1_ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ net107 sb_8__1_.mem_top_track_0.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_43_prog_clk net747 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output114_A net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_21.mux_l2_in_1__A1 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_3.mux_l2_in_1_ net331 sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_1__A0 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_1__A1 net214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_28.mux_l1_in_3_ net352 net27 sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_76_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4__S cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_331_ net60 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_46_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input75_A chany_top_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_3_ net235 sb_8__1_.mux_left_track_57.out cbx_8__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk
+ net832 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput125 net125 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput114 net114 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2_ net57 net68 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xoutput136 net136 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
XFILLER_87_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_3__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_8__1_.mem_bottom_track_13.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__A1 net87 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_22_prog_clk sb_8__1_.mem_top_track_6.mem_out\[2\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_55.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_55.out sky130_fd_sc_hd__clkbuf_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_2_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_3.mux_l1_in_2_ net228 net225 sb_8__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_314_ net74 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 chanx_left_in[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
Xinput16 chanx_left_in[20] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xinput49 chany_bottom_in[23] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_4
Xinput38 chany_bottom_in[13] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_31.mux_l1_in_0__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk net507 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net276 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__mux2_8
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__314__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net479
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_27.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ net738 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_0__S sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input38_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_4_ sb_8__1_.mux_left_track_45.out net31 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_2__S sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__1_.mux_top_track_28.mux_l3_in_0_ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_2__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_2__S sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk net794 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l2_in_2__A1 sb_8__1_.mux_left_track_41.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_0__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__309__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_49.out sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk net647 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_1__A0 sb_8__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_4.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__buf_4
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_14_prog_clk net566 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold5 net100 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net298 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ net408 VGND VGND VPWR
+ VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold405 sb_8__1_.mem_left_track_47.ccff_tail VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold416 sb_8__1_.mem_left_track_57.mem_out\[0\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold427 sb_8__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold449 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold438 sb_8__1_.mem_left_track_19.ccff_tail VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__302
+ VGND VGND VPWR VPWR net302 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__302/LO
+ sky130_fd_sc_hd__conb_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__260 VGND VGND VPWR VPWR net260
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__260/LO sky130_fd_sc_hd__conb_1
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__246 VGND VGND VPWR VPWR net246
+ cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__246/LO sky130_fd_sc_hd__conb_1
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_28.mux_l2_in_1_ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk
+ net764 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_1__A0 sb_8__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3__A0 net69 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_3_ net240 sb_8__1_.mux_left_track_49.out cbx_8__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_1__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__250 VGND VGND VPWR VPWR net250
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__250/LO sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_1__A0 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk net827
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold202 sb_8__1_.mem_bottom_track_37.ccff_tail VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold224 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold213 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ net844 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold235 cby_8__1_.cby_8__8_.mem_right_ipin_11.ccff_tail VGND VGND VPWR VPWR net601
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold246 cbx_8__1_.mem_top_ipin_10.ccff_head VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold257 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__322__A sb_8__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold268 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold279 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_4.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l3_in_0_ net406 cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[2\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_36_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_0.mux_l1_in_0_ net104 net109 sb_8__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_43_prog_clk net769 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_22_prog_clk net509 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_3.mux_l2_in_0_ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_4_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_1__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__317__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_28.mux_l1_in_2_ net9 net21 sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_2__A0 net437 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l2_in_2__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_330_ net59 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_3__S sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input68_A chany_top_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output224_A net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_0__S sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_17.mux_l2_in_1__324 VGND VGND VPWR VPWR net324 sb_8__1_.mux_left_track_17.mux_l2_in_1__324/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_2_ net15 cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ net410 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xoutput115 net115 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_1_ net405 cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xoutput137 net137 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.out cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__ebufn_8
Xsb_8__1_.mux_left_track_13.mux_l1_in_0_ net46 net72 sb_8__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_3__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__257 VGND VGND VPWR VPWR net257
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__257/LO sky130_fd_sc_hd__conb_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_9.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ net423 cbx_8__1_.mem_top_ipin_10.ccff_head VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net418 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_8__1_.mem_top_track_6.mem_out\[1\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_25.mux_l2_in_0_ sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_25.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l2_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_3.mux_l1_in_1_ net222 net49 sb_8__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_313_ net73 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 chanx_left_in[4] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
Xinput17 chanx_left_in[21] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput39 chany_bottom_in[14] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__247 VGND VGND VPWR VPWR net247
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__247/LO sky130_fd_sc_hd__conb_1
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_3_ net314 net29 sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk net645 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__330__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ net416 VGND VGND
+ VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_37.mux_l1_in_1__335 VGND VGND VPWR VPWR net335 sb_8__1_.mux_left_track_37.mux_l1_in_1__335/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_5.mem_out\[0\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ net568 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_3__A0 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_3__310 VGND VGND VPWR VPWR net310 sb_8__1_.mux_bottom_track_11.mux_l2_in_3__310/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_3_ sb_8__1_.mux_left_track_33.out net8 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2_ net74 net43 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ net708 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_8_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net305 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__mux2_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_9.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__280
+ VGND VGND VPWR VPWR net280 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__280/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_25.mux_l1_in_1_ net328 net227 sb_8__1_.mem_left_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA__325__A sb_8__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2__A1 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk net554 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3_ net251 net90 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_3__319 VGND VGND VPWR VPWR net319 sb_8__1_.mux_bottom_track_7.mux_l2_in_3__319/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input50_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold6 net891 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_14_prog_clk net590 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold417 sb_8__1_.mem_left_track_53.ccff_tail VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold406 sb_8__1_.mem_left_track_51.ccff_tail VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold439 sb_8__1_.mem_top_track_2.mem_out\[0\] VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold428 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_28.mux_l2_in_0_ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input98_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_3.mux_l4_in_0_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_2_ net29 sb_8__1_.mux_left_track_31.out cbx_8__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_1__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk net876
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_5_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_3__S sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_28_prog_clk net3
+ net233 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4_ sb_8__1_.mux_bottom_track_37.out
+ net36 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xhold214 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold203 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold225 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ net888 net229 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold269 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold247 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold236 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold258 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_4.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk sb_8__1_.mem_left_track_13.mem_out\[1\]
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold128_A cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk net470
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_21.mux_l2_in_1__326 VGND VGND VPWR VPWR net326 sb_8__1_.mux_left_track_21.mux_l2_in_1__326/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_43_prog_clk net649 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_35_prog_clk net495 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_33_prog_clk net588 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input13_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_3__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__A1 net414 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_28.mux_l1_in_1_ net45 net40 sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk net481
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l2_in_2__A1 net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_3.mux_l3_in_1_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_3__363 VGND VGND VPWR VPWR net363 cbx_8__1_.mux_top_ipin_13.mux_l2_in_3__363/LO
+ sky130_fd_sc_hd__conb_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3_ net242 net89 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output217_A net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk
+ net673 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_cbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_left_track_25.mux_l1_in_1__A1 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput116 net116 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xoutput138 net138 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_1__A0 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput149 net149 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_48_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold21_A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__328__A net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ net750 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_11_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_23_prog_clk sb_8__1_.mem_top_track_6.mem_out\[0\]
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_86_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_3__235 VGND VGND VPWR VPWR net235 cbx_8__1_.mux_top_ipin_4.mux_l2_in_3__235/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_left_track_3.mux_l1_in_0_ net55 net79 sb_8__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_312_ net72 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input80_A chany_top_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_left_in[22] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput29 chanx_left_in[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__292
+ VGND VGND VPWR VPWR net292 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__292/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_2_ net11 net23 sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk net608 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk net467 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk net742
+ net99 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_3__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4_ net66 net35 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_1__S sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_3__A1 net214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.out cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__ebufn_8
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_2_ sb_8__1_.mux_left_track_21.out net14 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_3__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_9.mux_l3_in_0_ net422 cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mem_top_ipin_9.mem_out\[2\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_16_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_left_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_25.mux_l1_in_0_ net63 net93 sb_8__1_.mem_left_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net379 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_88_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_2_ net59 cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_37.mux_l2_in_0_ sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk net864
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input43_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_14_prog_clk net592 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold7 net101 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_load_slew233_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold407 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[2\] VGND VGND VPWR VPWR net773
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold418 cbx_8__1_.mem_top_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold429 sb_8__1_.mem_bottom_track_29.mem_out\[1\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__1_.mux_top_track_2.mux_l2_in_3__350 VGND VGND VPWR VPWR net350 sb_8__1_.mux_top_track_2.mux_l2_in_3__350/LO
+ sky130_fd_sc_hd__conb_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_2__S sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk net849
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_2__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__336__A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_1__S sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_8_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_1_ net421 cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk net841
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_3_ net364 sb_8__1_.mux_left_track_53.out cbx_8__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3_ net73 net42 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xhold215 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold226 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold204 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net472 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold259 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold248 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold237 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_50_prog_clk
+ net780 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk net712
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_left_track_37.mux_l1_in_1_ net335 net225 sb_8__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk net870
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_43_prog_clk net653 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk net456 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_33_prog_clk net600 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_33.mux_l1_in_1__A1 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_28.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ net103 sb_8__1_.mem_top_track_28.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk net739
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_3.mux_l3_in_0_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_9.mux_l1_in_2_ sb_8__1_.mux_left_track_19.out net16 cbx_8__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_4_ sb_8__1_.mux_left_track_41.out net33 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_2_ net58 cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_52_prog_clk
+ net853 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_14_prog_clk net619 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l2_in_3__A1 sb_8__1_.mux_left_track_45.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput117 net117 VGND VGND VPWR VPWR ccff_tail_1 sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_1__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold14_A test_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__344__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_0__A0 sb_8__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk net721
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_14.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input108_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_0__S sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_311_ sb_8__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_19.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_19.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_42_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 net454 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input73_A chany_top_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk net861
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net295 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_1_ net216 net213 sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk net558 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk net868
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_56_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__339__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3_ net72 net41 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_2__A0 sb_8__1_.mux_left_track_21.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__265
+ VGND VGND VPWR VPWR net265 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__265/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_41.mux_l2_in_0__336 VGND VGND VPWR VPWR net336 sb_8__1_.mux_left_track_41.mux_l2_in_0__336/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_14.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_hold81_A chany_top_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net287 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__mux2_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk sb_8__1_.mem_top_track_20.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_left_track_29.mux_l1_in_0__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input36_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_4__A0 sb_8__1_.mux_left_track_41.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold408 sb_8__1_.mem_left_track_15.ccff_tail VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold419 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk net485
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk net606
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2__A1 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_2_ net27 cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[2\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__294
+ VGND VGND VPWR VPWR net294 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__294/LO
+ sky130_fd_sc_hd__conb_1
Xhold216 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold205 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net571
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold249 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold227 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold238 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk
+ net837 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_1__S sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net789
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_left_track_37.mux_l1_in_0_ net45 net75 sb_8__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__347__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk net527
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_43_prog_clk net484 net230 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_3__S sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_33_prog_clk net605 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_49.mux_l2_in_0_ net339 sb_8__1_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_49.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__303
+ VGND VGND VPWR VPWR net303 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__303/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_82_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_51.mux_l2_in_0_ sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_51.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__241 VGND VGND VPWR VPWR net241 cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__241/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_20.mux_l1_in_3__351 VGND VGND VPWR VPWR net351 sb_8__1_.mux_top_track_20.mux_l1_in_3__351/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__1_.mux_top_ipin_9.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk net854
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_54_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_3_ sb_8__1_.mux_left_track_29.out net10 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_14_prog_clk net638 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_3__311 VGND VGND VPWR VPWR net311 sb_8__1_.mux_bottom_track_13.mux_l1_in_3__311/LO
+ sky130_fd_sc_hd__conb_1
Xoutput118 net118 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_leaf_35_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net232
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ net70 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_2__S sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net833
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_19.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input66_A chany_top_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__270__A sb_8__1_.mux_left_track_51.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk
+ net595 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_left_track_19.mux_l2_in_1__A1 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk sb_8__1_.mem_left_track_7.mem_out\[0\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output222_A net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_51.mux_l1_in_1_ net341 net228 sb_8__1_.mem_left_track_51.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_0_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_5.mem_out\[1\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2_ net79 net48 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_37.mux_l1_in_0__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_2__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4__A1 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net379 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_88_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net720 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_3.mux_l2_in_1__331 VGND VGND VPWR VPWR net331 sb_8__1_.mux_left_track_3.mux_l2_in_1__331/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0__A1
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xcbx_8__1_.mux_top_ipin_14.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold74_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net412 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk net688
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mux_left_track_29.mux_l1_in_0__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_6.mux_l2_in_3_ net357 net5 sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xhold9 net112 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_0__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_3.mux_l1_in_1_ net218 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_4__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold409 cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_head VGND VGND VPWR VPWR net775
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l2_in_3__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net379 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_0__A0 sb_8__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__272
+ VGND VGND VPWR VPWR net272 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__272/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold206 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold217 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold228 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold239 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l2_in_3__A1 sb_8__1_.mux_left_track_53.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net541 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_2__S sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_33_prog_clk net567 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3__A0 net69 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input96_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__273__A sb_8__1_.mux_left_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2__A0 net77 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_2__A0 sb_8__1_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_25_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_6.mux_l4_in_0_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X
+ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X sb_8__1_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net284 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_9.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_66_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk cbx_8__1_.mem_top_ipin_8.mem_out\[1\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net261 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_2_ sb_8__1_.mux_left_track_17.out net17 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__287
+ VGND VGND VPWR VPWR net287 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__287/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_14_prog_clk net510 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input11_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput119 net119 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_4__A0 sb_8__1_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_45.mux_l1_in_0__A0 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_2__A0 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_49.mux_l1_in_0_ net223 net71 sb_8__1_.mem_left_track_49.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input3_A ccff_head_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_53.mux_l2_in_0__342 VGND VGND VPWR VPWR net342 sb_8__1_.mux_left_track_53.mux_l2_in_0__342/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_1__A0 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_31_prog_clk net573 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk net781
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_45_prog_clk
+ net551 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk net468
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_left_track_51.mux_l1_in_0_ net224 net76 sb_8__1_.mem_left_track_51.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_output215_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_6.mux_l3_in_1_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sb_8__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk net666
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_12.mux_l1_in_3_ net349 net15 sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_37.mux_l1_in_0__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_1__S sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net482 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_29.mux_l3_in_0_ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk net776
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_6.mux_l2_in_2_ net17 net60 sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_3.mux_l1_in_0_ net93 net79 sb_8__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__276__A net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk net711
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net269 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__mux2_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_29.mux_l2_in_1_ net313 sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_bottom_track_29.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_15_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input41_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_12.mux_l3_in_0_ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_23.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.out sky130_fd_sc_hd__clkbuf_2
XFILLER_62_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__262
+ VGND VGND VPWR VPWR net262 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__262/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold207 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold218 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold229 sb_8__1_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ net754 net232 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_load_slew231_A net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3_ net254 sb_8__1_.mux_bottom_track_45.out
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_1__A0 sb_8__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk net679 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.out sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_33_prog_clk net617 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input89_A chany_top_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk net689 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_53.mux_l1_in_0__A0 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold90 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_29.mux_l1_in_2_ net5 net17 sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_10_prog_clk cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_81_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.out sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_12.mux_l2_in_1_ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_5.mux_l2_in_1__A1 net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ net775 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_17_prog_clk net565 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__284__A sb_8__1_.mux_left_track_23.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_4__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_2__S sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__255 VGND VGND VPWR VPWR net255
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__255/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_31_prog_clk net528 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ net743 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xhold390 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_11.mux_l1_in_0__A0 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_6.mux_l3_in_0_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_52_prog_clk net2 net230 VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_299_ sb_8__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XFILLER_87_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l2_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk net777
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_12.mux_l1_in_2_ net7 net19 sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input106_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__A1 sb_8__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l2_in_3__A1 sb_8__1_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input71_A chany_top_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_2__S sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3_ net259 net90 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk net760
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_31.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_19.mux_l3_in_0_ sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_19.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_6.mux_l2_in_1_ net47 sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk net534 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_3__317 VGND VGND VPWR VPWR net317 sb_8__1_.mux_bottom_track_5.mux_l2_in_3__317/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__274
+ VGND VGND VPWR VPWR net274 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__274/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__292__A sb_8__1_.mux_left_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_21.mux_l3_in_0_ sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net379 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk net885
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_65_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_51.out sky130_fd_sc_hd__clkbuf_2
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_29.mux_l2_in_0_ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4_ sb_8__1_.mux_bottom_track_37.out
+ net36 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ net788 net230 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk cbx_8__1_.mem_top_ipin_11.mem_out\[2\]
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__287__A sb_8__1_.mux_left_track_17.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_0_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold208 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net574
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold219 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_3_ net358 sb_8__1_.mux_left_track_49.out cbx_8__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_3_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_left_track_19.mux_l2_in_1_ net325 net224 sb_8__1_.mem_left_track_19.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2_ net61 net72 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_top_track_6.mux_l1_in_2_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_1__S cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_33_prog_clk net585 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_15_prog_clk net808
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_21.mux_l2_in_1_ net326 net225 sb_8__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk net697 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_53.mux_l1_in_0__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold91 cbx_8__1_.mem_top_ipin_14.mem_out\[2\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold80 cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X VGND VGND VPWR VPWR
+ net446 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_2
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_29.mux_l1_in_1_ net214 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk net555
+ net229 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_3__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_1__A0 net214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net279 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_12.mux_l2_in_0_ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_3__361 VGND VGND VPWR VPWR net361 cbx_8__1_.mux_top_ipin_11.mux_l2_in_3__361/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_17_prog_clk net632 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_4_ sb_8__1_.mux_left_track_37.out net6 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l1_in_0__A0 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__276
+ VGND VGND VPWR VPWR net276 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__276/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_15.mux_l2_in_1__323 VGND VGND VPWR VPWR net323 sb_8__1_.mux_left_track_15.mux_l2_in_1__323/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_0__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_30_prog_clk net464 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_1__A0 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_0.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold380 cby_8__1_.cby_8__8_.mem_left_ipin_0.ccff_tail VGND VGND VPWR VPWR net746
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold391 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_11.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__295__A sb_8__1_.mux_left_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_1__S sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_298_ net87 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2__A0 net79 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_12.mux_l1_in_1_ net57 net43 sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_35.mux_l1_in_1__334 VGND VGND VPWR VPWR net334 sb_8__1_.mux_left_track_35.mux_l1_in_1__334/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_32_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__286
+ VGND VGND VPWR VPWR net286 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__286/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net265 net376 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_34_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input64_A chany_top_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_3_ net236 net448 cbx_8__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_77_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_38_prog_clk net650 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_2_ net399 cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk net457
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_12.mem_out\[1\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_21_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk net676 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_4__S cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_53.mux_l2_in_1__318 VGND VGND VPWR VPWR net318 sb_8__1_.mux_bottom_track_53.mux_l2_in_1__318/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_50_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_top_track_6.mux_l2_in_0_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net506 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l1_in_1__A0 sb_8__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_1__A0 net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_2__S sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net426 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_left_track_9.mux_l3_in_0_ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_8__1_.mem_top_track_44.mem_out\[0\]
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__306
+ VGND VGND VPWR VPWR net306 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__306/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_0__S sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2__A1 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3_ net73 net42 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input27_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk net483
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold209 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[2\] VGND VGND VPWR VPWR net575
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_2_ net29 cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_19.mux_l2_in_0_ net62 sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_19.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_1_ net41 cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l1_in_1__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_6.mux_l1_in_1_ net107 net105 sb_8__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_5.mux_l4_in_0_ net449 cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ cbx_8__1_.mem_top_ipin_5.ccff_tail VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_12_prog_clk net517
+ net229 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_21.mux_l2_in_0_ net58 sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_9.mux_l2_in_1_ net346 sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_left_track_9.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__298__A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold81 chany_top_in_0[28] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold92 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold70 chany_bottom_in[1] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__mux2_1
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_29.mux_l1_in_0_ net75 net70 sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_1__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_17_prog_clk net576 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_3_ sb_8__1_.mux_left_track_25.out net12 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input94_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_prog_clk clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2_ net79 net48 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__298
+ VGND VGND VPWR VPWR net298 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__298/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_5.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0_clk0_A clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net397 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_9.mux_l1_in_2_ net228 net225 sb_8__1_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_31_prog_clk net530 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_24_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3_ net247 sb_8__1_.mux_bottom_track_53.out
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold493_A sb_8__1_.mem_top_track_0.mem_out\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold381 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold370 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold392 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_297_ net86 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_12.mux_l1_in_0_ net107 net109 sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_3__S sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_2__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__269
+ VGND VGND VPWR VPWR net269 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__269/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input1_A ccff_head_0_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_2_ net4 sb_8__1_.mux_left_track_41.out cbx_8__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_38_prog_clk net640 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output213_A net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk cbx_8__1_.mem_top_ipin_14.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk net866
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_36.mux_l3_in_0_ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
X_349_ sb_8__1_.mux_top_track_12.out VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk net759 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4_ net65 net63 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_0.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4__A1 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_1__A1 net212 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l1_in_1__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk net706
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net375 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_4__A0 sb_8__1_.mux_left_track_41.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_36.mux_l2_in_1_ net353 sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net306 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__mux2_4
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk cbx_8__1_.mem_top_ipin_11.mem_out\[0\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l1_in_1__A1 net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_6.mux_l1_in_0_ net103 net109 sb_8__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3_ net252 net89 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_51.mux_l1_in_1__341 VGND VGND VPWR VPWR net341 sb_8__1_.mux_left_track_51.mux_l1_in_1__341/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_29_prog_clk clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2__A1 net68 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_9.mux_l2_in_0_ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__295
+ VGND VGND VPWR VPWR net295 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__295/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk net545 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ net451 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[2\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold82 net84 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold60 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold71 net45 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold93 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2__S cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_14_prog_clk_A clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_36.mux_l1_in_2_ net28 net10 sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net297 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_53_prog_clk_A clknet_2_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_17_prog_clk net607 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_2_ sb_8__1_.mux_left_track_13.out net19 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_19.mux_l1_in_0_ net38 net68 sb_8__1_.mem_left_track_19.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input87_A chany_top_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_0__S sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__A0 sb_8__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net232 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l1_in_1__A0 sb_8__1_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk
+ net795 net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_5.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_21.mux_l1_in_0_ net36 net66 sb_8__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_9.mux_l1_in_1_ net222 net44 sb_8__1_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_86_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_13.mux_l2_in_0__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_30_prog_clk net621 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_2_ net57 cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.out sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_44_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold360 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold371 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__1_.mux_left_track_33.mux_l2_in_0_ sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_33.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xhold382 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_hold486_A cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold393 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net268 net384 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_296_ net75 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3__A0 net73 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_0__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_1__A0 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3_ net243 sb_8__1_.mux_bottom_track_53.out
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk net682 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_23.mem_out\[1\]
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_23.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_1__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_1_ net33 cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xhold190 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_38_prog_clk net646 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_3_ net360 sb_8__1_.mux_left_track_57.out cbx_8__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk net716
+ net231 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_348_ net49 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_279_ sb_8__1_.mux_left_track_33.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3_ sb_8__1_.mux_bottom_track_29.out
+ net40 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_39_prog_clk net629 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_2__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_1__S sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_52_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_33.mux_l1_in_1_ net333 net223 sb_8__1_.mem_left_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk net714
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_55.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input104_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_2__A0 net399 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_30_prog_clk net476 net233 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l1_in_1__A1 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net301 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4_ net65 net63 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk net692 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_4__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_5.mux_l1_in_2_ sb_8__1_.mux_left_track_23.out net13 cbx_8__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_1__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_4_ sb_8__1_.mux_left_track_45.out net31 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_36.mux_l2_in_0_ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk net727
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l1_in_1__A0 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_left_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_1__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2_ net58 net66 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_prog_clk_A clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_10.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk net690 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input32_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold50 cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net416 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold61 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold83 cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X VGND VGND VPWR VPWR net449
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold72 cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X VGND VGND
+ VPWR VPWR net438 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold94 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l2_in_3__A1 sb_8__1_.mux_left_track_53.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3__A0 net70 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_3 cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_21.mux_l2_in_0__A0 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_36.mux_l1_in_1_ net22 net39 sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net114 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold520 sb_8__1_.mem_bottom_track_21.mem_out\[1\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net379 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__sdfrtp_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_17_prog_clk net615 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_3_ net365 net88 cbx_8__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ sb_8__1_.mem_bottom_track_29.mem_out\[0\] net230 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_29.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_10.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_9.mux_l1_in_0_ net51 net74 sb_8__1_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk
+ net883 net231 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_30_prog_clk net593 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_prog_clk clknet_2_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l1_in_2__A0 sb_8__1_.mux_left_track_23.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold350 sb_8__1_.mem_top_track_10.ccff_tail VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold361 cbx_8__1_.mem_top_ipin_10.ccff_tail VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_2__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold383 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xhold372 sb_8__1_.mem_bottom_track_45.mem_out\[0\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold394 sb_8__1_.mem_left_track_29.ccff_tail VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_364_ net114 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_1
X_295_ sb_8__1_.mux_left_track_1.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net229 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net231 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_2__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net368 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net379 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold88_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_3_ net311 net15 sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_59_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_2_ net57 cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk net694 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net821
+ net230 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_23.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net230 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_1.mem_out\[2\]
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_1__A1 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold180 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold191 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_38_prog_clk net657 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk net498
+ net230 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk net736 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_2_ net15 cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_347_ net48 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
X_278_ sb_8__1_.mux_left_track_35.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2_ net78 net47 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_39_prog_clk net631 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l2_in_1__A0 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_15.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X net116 VGND VGND VPWR VPWR
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_33.mux_l1_in_0_ net57 net87 sb_8__1_.mem_left_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ net383 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk net783
+ net232 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_55.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_3__314 VGND VGND VPWR VPWR net314 sb_8__1_.mux_bottom_track_3.mux_l2_in_3__314/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_45.mux_l2_in_0_ net337 sb_8__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_45.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input62_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk net741 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk net702 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3_ sb_8__1_.mux_bottom_track_29.out
+ net40 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk net544 net231 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_33_prog_clk_A clknet_2_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__301__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_5.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_1__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_3_ sb_8__1_.mux_left_track_33.out net8 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l1_in_1__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0__A1
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_13.mux_l3_in_0_ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_15.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_1__A1 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_1_ net35 cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold70_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__281
+ VGND VGND VPWR VPWR net281 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__281/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net288 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__mux2_4
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__307
+ VGND VGND VPWR VPWR net307 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__307/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_38_prog_clk clknet_2_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk
+ net873 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_2__A0 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold40 cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X VGND VGND
+ VPWR VPWR net406 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold62 chany_top_in_0[2] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold51 cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold73 cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X VGND VGND
+ VPWR VPWR net439 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input25_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold95 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold84 chany_bottom_in[3] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_90_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_4 net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_0__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_3__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_36.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ net104 sb_8__1_.mem_top_track_36.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xhold510 sb_8__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold521 sb_8__1_.mem_bottom_track_3.mem_out\[0\] VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk net610 net232 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_13.mux_l2_in_1_ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_2_ net32 sb_8__1_.mux_left_track_31.out cbx_8__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_13_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_2__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_1__S sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2_ sb_8__1_.mux_bottom_track_21.out
+ net44 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ net518 net229 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_10.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__253 VGND VGND VPWR VPWR net253
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__253/LO sky130_fd_sc_hd__conb_1
XANTENNA_hold33_A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_30_prog_clk net604 net233 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
.ends

