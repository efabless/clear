magic
tech sky130A
magscale 1 2
timestamp 1679318170
<< viali >>
rect 33517 54281 33551 54315
rect 36277 54213 36311 54247
rect 46857 54213 46891 54247
rect 1777 54145 1811 54179
rect 4353 54145 4387 54179
rect 6929 54145 6963 54179
rect 9597 54145 9631 54179
rect 12265 54145 12299 54179
rect 15025 54145 15059 54179
rect 17693 54145 17727 54179
rect 20269 54145 20303 54179
rect 22845 54145 22879 54179
rect 25697 54145 25731 54179
rect 28365 54145 28399 54179
rect 31033 54145 31067 54179
rect 33701 54145 33735 54179
rect 38853 54145 38887 54179
rect 41521 54145 41555 54179
rect 44189 54145 44223 54179
rect 48329 54145 48363 54179
rect 49065 54145 49099 54179
rect 2053 54077 2087 54111
rect 4629 54077 4663 54111
rect 7297 54077 7331 54111
rect 9965 54077 9999 54111
rect 12633 54077 12667 54111
rect 15301 54077 15335 54111
rect 17969 54077 18003 54111
rect 20545 54077 20579 54111
rect 23121 54077 23155 54111
rect 36461 54009 36495 54043
rect 25513 53941 25547 53975
rect 28181 53941 28215 53975
rect 30849 53941 30883 53975
rect 39037 53941 39071 53975
rect 41705 53941 41739 53975
rect 44373 53941 44407 53975
rect 46949 53941 46983 53975
rect 48513 53941 48547 53975
rect 49249 53941 49283 53975
rect 47869 53533 47903 53567
rect 48329 53533 48363 53567
rect 49065 53533 49099 53567
rect 47685 53397 47719 53431
rect 48513 53397 48547 53431
rect 49249 53397 49283 53431
rect 9873 53193 9907 53227
rect 9781 53057 9815 53091
rect 49065 53057 49099 53091
rect 49249 52853 49283 52887
rect 49341 52445 49375 52479
rect 48973 52377 49007 52411
rect 12817 52105 12851 52139
rect 12725 51969 12759 52003
rect 16313 51561 16347 51595
rect 17325 51493 17359 51527
rect 14933 51357 14967 51391
rect 16497 51357 16531 51391
rect 17141 51289 17175 51323
rect 48973 51289 49007 51323
rect 49341 51289 49375 51323
rect 15025 51221 15059 51255
rect 48973 50881 49007 50915
rect 49065 50677 49099 50711
rect 15301 50473 15335 50507
rect 19625 50473 19659 50507
rect 15669 50405 15703 50439
rect 15209 50269 15243 50303
rect 19533 50201 19567 50235
rect 49157 49793 49191 49827
rect 49341 49725 49375 49759
rect 21005 49385 21039 49419
rect 23029 49385 23063 49419
rect 20913 49113 20947 49147
rect 22937 49113 22971 49147
rect 49157 49113 49191 49147
rect 49341 49113 49375 49147
rect 16129 48229 16163 48263
rect 14381 48161 14415 48195
rect 14657 48025 14691 48059
rect 49157 48025 49191 48059
rect 49249 47957 49283 47991
rect 19809 47753 19843 47787
rect 19349 47617 19383 47651
rect 20304 47617 20338 47651
rect 49341 47617 49375 47651
rect 19533 47413 19567 47447
rect 20407 47413 20441 47447
rect 49157 47413 49191 47447
rect 25697 47073 25731 47107
rect 22328 47005 22362 47039
rect 22431 46937 22465 46971
rect 25881 46937 25915 46971
rect 27537 46937 27571 46971
rect 23213 46529 23247 46563
rect 49341 46529 49375 46563
rect 23397 46461 23431 46495
rect 24777 46461 24811 46495
rect 49157 46325 49191 46359
rect 17509 46121 17543 46155
rect 21465 46121 21499 46155
rect 21649 46121 21683 46155
rect 17325 45985 17359 46019
rect 27353 45985 27387 46019
rect 28917 45985 28951 46019
rect 17141 45917 17175 45951
rect 21189 45917 21223 45951
rect 24628 45917 24662 45951
rect 49341 45917 49375 45951
rect 24731 45849 24765 45883
rect 27537 45849 27571 45883
rect 49157 45781 49191 45815
rect 25916 45441 25950 45475
rect 29561 45441 29595 45475
rect 29745 45373 29779 45407
rect 31401 45373 31435 45407
rect 26019 45237 26053 45271
rect 21189 45033 21223 45067
rect 19717 44897 19751 44931
rect 19441 44829 19475 44863
rect 49341 44829 49375 44863
rect 49157 44693 49191 44727
rect 20637 44489 20671 44523
rect 22937 44489 22971 44523
rect 20177 44353 20211 44387
rect 22477 44353 22511 44387
rect 49157 44353 49191 44387
rect 19993 44285 20027 44319
rect 49341 44217 49375 44251
rect 22569 44149 22603 44183
rect 41797 43809 41831 43843
rect 41521 43741 41555 43775
rect 43269 43605 43303 43639
rect 49157 43265 49191 43299
rect 49341 43129 49375 43163
rect 49157 42585 49191 42619
rect 49249 42517 49283 42551
rect 21465 42313 21499 42347
rect 23029 42313 23063 42347
rect 21005 42177 21039 42211
rect 22385 42177 22419 42211
rect 20821 42109 20855 42143
rect 22569 42109 22603 42143
rect 23305 41769 23339 41803
rect 21557 41633 21591 41667
rect 21833 41497 21867 41531
rect 49157 41497 49191 41531
rect 49249 41429 49283 41463
rect 49341 41089 49375 41123
rect 49157 40885 49191 40919
rect 49157 40137 49191 40171
rect 49341 40001 49375 40035
rect 49341 39389 49375 39423
rect 49157 39253 49191 39287
rect 49341 38301 49375 38335
rect 49157 38165 49191 38199
rect 49157 37825 49191 37859
rect 49341 37689 49375 37723
rect 20453 37213 20487 37247
rect 20269 37077 20303 37111
rect 49157 36737 49191 36771
rect 49249 36533 49283 36567
rect 49341 36125 49375 36159
rect 49157 35989 49191 36023
rect 49341 35037 49375 35071
rect 49157 34901 49191 34935
rect 24685 34697 24719 34731
rect 49157 34697 49191 34731
rect 49341 34561 49375 34595
rect 22937 34493 22971 34527
rect 23200 34357 23234 34391
rect 22845 34153 22879 34187
rect 42165 34085 42199 34119
rect 41429 34017 41463 34051
rect 41521 34017 41555 34051
rect 42717 34017 42751 34051
rect 23029 33949 23063 33983
rect 42533 33949 42567 33983
rect 41337 33881 41371 33915
rect 40417 33813 40451 33847
rect 40969 33813 41003 33847
rect 42625 33813 42659 33847
rect 43453 33813 43487 33847
rect 43085 33609 43119 33643
rect 42993 33473 43027 33507
rect 49341 33473 49375 33507
rect 43269 33405 43303 33439
rect 42625 33269 42659 33303
rect 43821 33269 43855 33303
rect 49157 33269 49191 33303
rect 49341 32861 49375 32895
rect 49157 32725 49191 32759
rect 38485 32317 38519 32351
rect 38761 32317 38795 32351
rect 40233 32181 40267 32215
rect 42809 31977 42843 32011
rect 41797 31909 41831 31943
rect 43269 31909 43303 31943
rect 49157 31909 49191 31943
rect 40325 31841 40359 31875
rect 43821 31841 43855 31875
rect 40049 31773 40083 31807
rect 43637 31773 43671 31807
rect 43729 31773 43763 31807
rect 49341 31773 49375 31807
rect 43729 31433 43763 31467
rect 43821 31433 43855 31467
rect 33977 31297 34011 31331
rect 34805 31297 34839 31331
rect 34897 31297 34931 31331
rect 37933 31297 37967 31331
rect 40325 31297 40359 31331
rect 49341 31297 49375 31331
rect 35081 31229 35115 31263
rect 38209 31229 38243 31263
rect 40601 31229 40635 31263
rect 43913 31229 43947 31263
rect 34437 31161 34471 31195
rect 39681 31093 39715 31127
rect 42073 31093 42107 31127
rect 43361 31093 43395 31127
rect 49157 31093 49191 31127
rect 22293 30889 22327 30923
rect 22937 30889 22971 30923
rect 43177 30889 43211 30923
rect 40785 30753 40819 30787
rect 41429 30753 41463 30787
rect 22477 30685 22511 30719
rect 23121 30685 23155 30719
rect 40601 30685 40635 30719
rect 32781 30617 32815 30651
rect 33517 30617 33551 30651
rect 35449 30617 35483 30651
rect 36277 30617 36311 30651
rect 41705 30617 41739 30651
rect 40233 30549 40267 30583
rect 40693 30549 40727 30583
rect 34621 30277 34655 30311
rect 35449 30277 35483 30311
rect 41153 30277 41187 30311
rect 35541 30209 35575 30243
rect 38117 30209 38151 30243
rect 42625 30209 42659 30243
rect 49341 30209 49375 30243
rect 35633 30141 35667 30175
rect 38393 30141 38427 30175
rect 41245 30141 41279 30175
rect 41337 30141 41371 30175
rect 42901 30141 42935 30175
rect 35081 30005 35115 30039
rect 39865 30005 39899 30039
rect 40785 30005 40819 30039
rect 44373 30005 44407 30039
rect 49157 30005 49191 30039
rect 31572 29801 31606 29835
rect 35541 29665 35575 29699
rect 43545 29665 43579 29699
rect 31309 29597 31343 29631
rect 35357 29597 35391 29631
rect 36185 29597 36219 29631
rect 49341 29597 49375 29631
rect 34069 29529 34103 29563
rect 35265 29529 35299 29563
rect 42809 29529 42843 29563
rect 33057 29461 33091 29495
rect 34897 29461 34931 29495
rect 49157 29461 49191 29495
rect 34253 29257 34287 29291
rect 34621 29257 34655 29291
rect 35541 29257 35575 29291
rect 44373 29257 44407 29291
rect 32965 29189 32999 29223
rect 36093 29189 36127 29223
rect 32873 29121 32907 29155
rect 34713 29121 34747 29155
rect 36001 29121 36035 29155
rect 37473 29121 37507 29155
rect 39681 29121 39715 29155
rect 42625 29121 42659 29155
rect 33149 29053 33183 29087
rect 33793 29053 33827 29087
rect 34805 29053 34839 29087
rect 36185 29053 36219 29087
rect 39221 29053 39255 29087
rect 39957 29053 39991 29087
rect 32505 28985 32539 29019
rect 35633 28985 35667 29019
rect 37736 28917 37770 28951
rect 41429 28917 41463 28951
rect 42882 28917 42916 28951
rect 36185 28713 36219 28747
rect 30297 28577 30331 28611
rect 33241 28577 33275 28611
rect 35449 28577 35483 28611
rect 38761 28577 38795 28611
rect 42257 28577 42291 28611
rect 37013 28509 37047 28543
rect 39405 28509 39439 28543
rect 40049 28509 40083 28543
rect 49341 28509 49375 28543
rect 30573 28441 30607 28475
rect 32505 28441 32539 28475
rect 35265 28441 35299 28475
rect 37289 28441 37323 28475
rect 40325 28441 40359 28475
rect 42533 28441 42567 28475
rect 32045 28373 32079 28407
rect 34897 28373 34931 28407
rect 35357 28373 35391 28407
rect 41797 28373 41831 28407
rect 44005 28373 44039 28407
rect 49157 28373 49191 28407
rect 23673 28169 23707 28203
rect 31493 28169 31527 28203
rect 38393 28169 38427 28203
rect 40233 28169 40267 28203
rect 43913 28169 43947 28203
rect 44005 28169 44039 28203
rect 24041 28101 24075 28135
rect 28825 28101 28859 28135
rect 35437 28101 35471 28135
rect 41797 28101 41831 28135
rect 24133 28033 24167 28067
rect 28549 28033 28583 28067
rect 31401 28033 31435 28067
rect 33241 28033 33275 28067
rect 38485 28033 38519 28067
rect 40141 28033 40175 28067
rect 41705 28033 41739 28067
rect 49341 28033 49375 28067
rect 24225 27965 24259 27999
rect 31585 27965 31619 27999
rect 33517 27965 33551 27999
rect 36185 27965 36219 27999
rect 38577 27965 38611 27999
rect 40325 27965 40359 27999
rect 41889 27965 41923 27999
rect 44097 27965 44131 27999
rect 31033 27897 31067 27931
rect 30297 27829 30331 27863
rect 34989 27829 35023 27863
rect 38025 27829 38059 27863
rect 39773 27829 39807 27863
rect 41337 27829 41371 27863
rect 43545 27829 43579 27863
rect 49157 27829 49191 27863
rect 24856 27625 24890 27659
rect 31020 27625 31054 27659
rect 40417 27625 40451 27659
rect 37289 27557 37323 27591
rect 24593 27489 24627 27523
rect 30757 27489 30791 27523
rect 32505 27489 32539 27523
rect 33517 27489 33551 27523
rect 36093 27489 36127 27523
rect 37933 27489 37967 27523
rect 43913 27489 43947 27523
rect 33333 27421 33367 27455
rect 35909 27421 35943 27455
rect 37657 27421 37691 27455
rect 38669 27421 38703 27455
rect 41521 27421 41555 27455
rect 41981 27421 42015 27455
rect 43729 27421 43763 27455
rect 43821 27421 43855 27455
rect 37749 27353 37783 27387
rect 42717 27353 42751 27387
rect 26341 27285 26375 27319
rect 32965 27285 32999 27319
rect 33425 27285 33459 27319
rect 35541 27285 35575 27319
rect 36001 27285 36035 27319
rect 43361 27285 43395 27319
rect 31401 27081 31435 27115
rect 31493 27081 31527 27115
rect 33149 27081 33183 27115
rect 35265 27081 35299 27115
rect 39497 27081 39531 27115
rect 41705 27081 41739 27115
rect 41797 27081 41831 27115
rect 44649 27081 44683 27115
rect 44741 27081 44775 27115
rect 28733 27013 28767 27047
rect 28457 26945 28491 26979
rect 33241 26945 33275 26979
rect 49341 26945 49375 26979
rect 31585 26877 31619 26911
rect 33333 26877 33367 26911
rect 35357 26877 35391 26911
rect 35449 26877 35483 26911
rect 37749 26877 37783 26911
rect 38025 26877 38059 26911
rect 41889 26877 41923 26911
rect 44925 26877 44959 26911
rect 34897 26809 34931 26843
rect 30205 26741 30239 26775
rect 31033 26741 31067 26775
rect 32781 26741 32815 26775
rect 41337 26741 41371 26775
rect 44281 26741 44315 26775
rect 49157 26741 49191 26775
rect 29193 26537 29227 26571
rect 34897 26537 34931 26571
rect 38209 26469 38243 26503
rect 41889 26469 41923 26503
rect 27445 26401 27479 26435
rect 30573 26401 30607 26435
rect 30849 26401 30883 26435
rect 32321 26401 32355 26435
rect 35357 26401 35391 26435
rect 35449 26401 35483 26435
rect 38669 26401 38703 26435
rect 38853 26401 38887 26435
rect 35265 26333 35299 26367
rect 37749 26333 37783 26367
rect 38577 26333 38611 26367
rect 40141 26333 40175 26367
rect 42533 26333 42567 26367
rect 48053 26333 48087 26367
rect 48513 26333 48547 26367
rect 48789 26333 48823 26367
rect 27721 26265 27755 26299
rect 40417 26265 40451 26299
rect 43545 26265 43579 26299
rect 43729 26265 43763 26299
rect 34897 25993 34931 26027
rect 35725 25993 35759 26027
rect 35817 25993 35851 26027
rect 41705 25993 41739 26027
rect 30481 25925 30515 25959
rect 31401 25925 31435 25959
rect 45109 25925 45143 25959
rect 27169 25857 27203 25891
rect 31309 25857 31343 25891
rect 32505 25857 32539 25891
rect 38485 25857 38519 25891
rect 42625 25857 42659 25891
rect 44833 25857 44867 25891
rect 27445 25789 27479 25823
rect 31493 25789 31527 25823
rect 33149 25789 33183 25823
rect 33425 25789 33459 25823
rect 35909 25789 35943 25823
rect 38761 25789 38795 25823
rect 41797 25789 41831 25823
rect 41981 25789 42015 25823
rect 42901 25789 42935 25823
rect 40233 25721 40267 25755
rect 28917 25653 28951 25687
rect 30941 25653 30975 25687
rect 35357 25653 35391 25687
rect 37933 25653 37967 25687
rect 41337 25653 41371 25687
rect 44373 25653 44407 25687
rect 46581 25653 46615 25687
rect 34897 25449 34931 25483
rect 44005 25449 44039 25483
rect 33609 25381 33643 25415
rect 41797 25381 41831 25415
rect 45201 25381 45235 25415
rect 30665 25313 30699 25347
rect 30757 25313 30791 25347
rect 34069 25313 34103 25347
rect 34161 25313 34195 25347
rect 35449 25313 35483 25347
rect 38025 25313 38059 25347
rect 40325 25313 40359 25347
rect 42257 25313 42291 25347
rect 45661 25313 45695 25347
rect 45845 25313 45879 25347
rect 36921 25245 36955 25279
rect 37749 25245 37783 25279
rect 40049 25245 40083 25279
rect 47961 25245 47995 25279
rect 49157 25245 49191 25279
rect 31401 25177 31435 25211
rect 33977 25177 34011 25211
rect 35265 25177 35299 25211
rect 37841 25177 37875 25211
rect 42533 25177 42567 25211
rect 30205 25109 30239 25143
rect 30573 25109 30607 25143
rect 32873 25109 32907 25143
rect 35357 25109 35391 25143
rect 36737 25109 36771 25143
rect 37381 25109 37415 25143
rect 45569 25109 45603 25143
rect 31401 24905 31435 24939
rect 36553 24905 36587 24939
rect 31493 24769 31527 24803
rect 32689 24769 32723 24803
rect 36645 24769 36679 24803
rect 37749 24769 37783 24803
rect 38577 24769 38611 24803
rect 42993 24769 43027 24803
rect 43085 24769 43119 24803
rect 44189 24769 44223 24803
rect 47961 24769 47995 24803
rect 31585 24701 31619 24735
rect 32781 24701 32815 24735
rect 32965 24701 32999 24735
rect 33609 24701 33643 24735
rect 33885 24701 33919 24735
rect 36737 24701 36771 24735
rect 43177 24701 43211 24735
rect 44465 24701 44499 24735
rect 45937 24701 45971 24735
rect 49157 24701 49191 24735
rect 31033 24565 31067 24599
rect 32321 24565 32355 24599
rect 35357 24565 35391 24599
rect 36185 24565 36219 24599
rect 37841 24565 37875 24599
rect 38393 24565 38427 24599
rect 42625 24565 42659 24599
rect 25973 24361 26007 24395
rect 28457 24361 28491 24395
rect 33701 24293 33735 24327
rect 26617 24225 26651 24259
rect 28917 24225 28951 24259
rect 29009 24225 29043 24259
rect 30021 24225 30055 24259
rect 31953 24225 31987 24259
rect 35357 24225 35391 24259
rect 35449 24225 35483 24259
rect 44097 24225 44131 24259
rect 45753 24225 45787 24259
rect 29745 24157 29779 24191
rect 35265 24157 35299 24191
rect 36277 24157 36311 24191
rect 38945 24157 38979 24191
rect 41705 24157 41739 24191
rect 43913 24157 43947 24191
rect 44005 24157 44039 24191
rect 46581 24157 46615 24191
rect 26341 24089 26375 24123
rect 28825 24089 28859 24123
rect 32229 24089 32263 24123
rect 45569 24089 45603 24123
rect 45661 24089 45695 24123
rect 26433 24021 26467 24055
rect 31493 24021 31527 24055
rect 34897 24021 34931 24055
rect 36093 24021 36127 24055
rect 43545 24021 43579 24055
rect 45201 24021 45235 24055
rect 46397 24021 46431 24055
rect 25605 23817 25639 23851
rect 25973 23817 26007 23851
rect 32597 23749 32631 23783
rect 36553 23749 36587 23783
rect 38669 23749 38703 23783
rect 38761 23749 38795 23783
rect 40325 23749 40359 23783
rect 40417 23749 40451 23783
rect 41153 23749 41187 23783
rect 43269 23749 43303 23783
rect 44097 23749 44131 23783
rect 27169 23681 27203 23715
rect 29469 23681 29503 23715
rect 32321 23681 32355 23715
rect 35357 23681 35391 23715
rect 37841 23681 37875 23715
rect 44649 23681 44683 23715
rect 47961 23681 47995 23715
rect 26065 23613 26099 23647
rect 26157 23613 26191 23647
rect 27445 23613 27479 23647
rect 29745 23613 29779 23647
rect 31217 23613 31251 23647
rect 34069 23613 34103 23647
rect 35449 23613 35483 23647
rect 35541 23613 35575 23647
rect 36645 23613 36679 23647
rect 36829 23613 36863 23647
rect 38945 23613 38979 23647
rect 40601 23613 40635 23647
rect 41889 23613 41923 23647
rect 44925 23613 44959 23647
rect 49157 23613 49191 23647
rect 38301 23545 38335 23579
rect 28917 23477 28951 23511
rect 34989 23477 35023 23511
rect 36185 23477 36219 23511
rect 39957 23477 39991 23511
rect 46397 23477 46431 23511
rect 26341 23273 26375 23307
rect 43453 23273 43487 23307
rect 38117 23205 38151 23239
rect 42257 23205 42291 23239
rect 24869 23137 24903 23171
rect 30297 23137 30331 23171
rect 31401 23137 31435 23171
rect 31493 23137 31527 23171
rect 33425 23137 33459 23171
rect 38761 23137 38795 23171
rect 40509 23137 40543 23171
rect 43913 23137 43947 23171
rect 44097 23137 44131 23171
rect 24593 23069 24627 23103
rect 30113 23069 30147 23103
rect 30205 23069 30239 23103
rect 31309 23069 31343 23103
rect 33241 23069 33275 23103
rect 34253 23069 34287 23103
rect 38485 23069 38519 23103
rect 38577 23069 38611 23103
rect 39497 23069 39531 23103
rect 42901 23069 42935 23103
rect 46121 23069 46155 23103
rect 47961 23069 47995 23103
rect 32413 23001 32447 23035
rect 40785 23001 40819 23035
rect 43821 23001 43855 23035
rect 45293 23001 45327 23035
rect 45477 23001 45511 23035
rect 49157 23001 49191 23035
rect 29745 22933 29779 22967
rect 30941 22933 30975 22967
rect 32873 22933 32907 22967
rect 33333 22933 33367 22967
rect 39313 22933 39347 22967
rect 45937 22933 45971 22967
rect 33885 22729 33919 22763
rect 37841 22729 37875 22763
rect 41613 22729 41647 22763
rect 42993 22729 43027 22763
rect 43085 22729 43119 22763
rect 46673 22729 46707 22763
rect 37933 22661 37967 22695
rect 44005 22661 44039 22695
rect 44189 22661 44223 22695
rect 33793 22593 33827 22627
rect 39037 22593 39071 22627
rect 44925 22593 44959 22627
rect 33977 22525 34011 22559
rect 38025 22525 38059 22559
rect 39313 22525 39347 22559
rect 40785 22525 40819 22559
rect 41705 22525 41739 22559
rect 41797 22525 41831 22559
rect 43269 22525 43303 22559
rect 45201 22525 45235 22559
rect 33425 22457 33459 22491
rect 41245 22457 41279 22491
rect 37473 22389 37507 22423
rect 42625 22389 42659 22423
rect 26052 22185 26086 22219
rect 30192 22185 30226 22219
rect 42612 22185 42646 22219
rect 37565 22117 37599 22151
rect 28457 22049 28491 22083
rect 28549 22049 28583 22083
rect 36829 22049 36863 22083
rect 36921 22049 36955 22083
rect 39221 22049 39255 22083
rect 39405 22049 39439 22083
rect 45477 22049 45511 22083
rect 25789 21981 25823 22015
rect 28365 21981 28399 22015
rect 29929 21981 29963 22015
rect 37749 21981 37783 22015
rect 39129 21981 39163 22015
rect 42349 21981 42383 22015
rect 45201 21981 45235 22015
rect 47961 21981 47995 22015
rect 49157 21981 49191 22015
rect 36737 21913 36771 21947
rect 27537 21845 27571 21879
rect 27997 21845 28031 21879
rect 31677 21845 31711 21879
rect 36369 21845 36403 21879
rect 38761 21845 38795 21879
rect 44097 21845 44131 21879
rect 46949 21845 46983 21879
rect 25513 21641 25547 21675
rect 27169 21641 27203 21675
rect 30665 21641 30699 21675
rect 31125 21641 31159 21675
rect 33057 21641 33091 21675
rect 37933 21641 37967 21675
rect 39037 21641 39071 21675
rect 43177 21641 43211 21675
rect 45753 21641 45787 21675
rect 25973 21573 26007 21607
rect 32965 21573 32999 21607
rect 39129 21573 39163 21607
rect 44281 21573 44315 21607
rect 25881 21505 25915 21539
rect 27537 21505 27571 21539
rect 31033 21505 31067 21539
rect 37841 21505 37875 21539
rect 43269 21505 43303 21539
rect 47961 21505 47995 21539
rect 26157 21437 26191 21471
rect 27629 21437 27663 21471
rect 27721 21437 27755 21471
rect 28457 21437 28491 21471
rect 28733 21437 28767 21471
rect 31217 21437 31251 21471
rect 33149 21437 33183 21471
rect 34805 21437 34839 21471
rect 35081 21437 35115 21471
rect 38117 21437 38151 21471
rect 39221 21437 39255 21471
rect 43361 21437 43395 21471
rect 44005 21437 44039 21471
rect 49157 21437 49191 21471
rect 37473 21369 37507 21403
rect 24961 21301 24995 21335
rect 30205 21301 30239 21335
rect 32597 21301 32631 21335
rect 36553 21301 36587 21335
rect 38669 21301 38703 21335
rect 42809 21301 42843 21335
rect 24593 21097 24627 21131
rect 28825 21097 28859 21131
rect 32505 21097 32539 21131
rect 36737 21097 36771 21131
rect 38025 21097 38059 21131
rect 41981 21097 42015 21131
rect 42901 21029 42935 21063
rect 25237 20961 25271 20995
rect 26433 20961 26467 20995
rect 31033 20961 31067 20995
rect 33517 20961 33551 20995
rect 34989 20961 35023 20995
rect 35265 20961 35299 20995
rect 43453 20961 43487 20995
rect 24961 20893 24995 20927
rect 26157 20893 26191 20927
rect 30757 20893 30791 20927
rect 33425 20893 33459 20927
rect 38853 20893 38887 20927
rect 40233 20893 40267 20927
rect 43269 20893 43303 20927
rect 44281 20893 44315 20927
rect 28181 20825 28215 20859
rect 33333 20825 33367 20859
rect 40509 20825 40543 20859
rect 43361 20825 43395 20859
rect 25053 20757 25087 20791
rect 32965 20757 32999 20791
rect 38669 20757 38703 20791
rect 28917 20553 28951 20587
rect 31769 20553 31803 20587
rect 36185 20553 36219 20587
rect 36645 20553 36679 20587
rect 44373 20553 44407 20587
rect 30297 20485 30331 20519
rect 43085 20485 43119 20519
rect 33977 20417 34011 20451
rect 36553 20417 36587 20451
rect 42901 20417 42935 20451
rect 44281 20417 44315 20451
rect 45293 20417 45327 20451
rect 47961 20417 47995 20451
rect 23765 20349 23799 20383
rect 24041 20349 24075 20383
rect 27169 20349 27203 20383
rect 27445 20349 27479 20383
rect 30021 20349 30055 20383
rect 34253 20349 34287 20383
rect 36737 20349 36771 20383
rect 38393 20349 38427 20383
rect 38669 20349 38703 20383
rect 44557 20349 44591 20383
rect 49157 20349 49191 20383
rect 25513 20213 25547 20247
rect 35725 20213 35759 20247
rect 40141 20213 40175 20247
rect 43913 20213 43947 20247
rect 29193 20009 29227 20043
rect 32860 20009 32894 20043
rect 34897 20009 34931 20043
rect 40306 20009 40340 20043
rect 41797 20009 41831 20043
rect 42520 20009 42554 20043
rect 24593 19873 24627 19907
rect 27445 19873 27479 19907
rect 39129 19873 39163 19907
rect 40049 19873 40083 19907
rect 42257 19873 42291 19907
rect 32597 19805 32631 19839
rect 35081 19805 35115 19839
rect 36645 19805 36679 19839
rect 38853 19805 38887 19839
rect 38945 19805 38979 19839
rect 45385 19805 45419 19839
rect 47961 19805 47995 19839
rect 24869 19737 24903 19771
rect 27721 19737 27755 19771
rect 49157 19737 49191 19771
rect 26341 19669 26375 19703
rect 34345 19669 34379 19703
rect 36461 19669 36495 19703
rect 38485 19669 38519 19703
rect 44005 19669 44039 19703
rect 45201 19669 45235 19703
rect 23581 19465 23615 19499
rect 28825 19465 28859 19499
rect 29285 19465 29319 19499
rect 33885 19465 33919 19499
rect 35081 19465 35115 19499
rect 35173 19465 35207 19499
rect 38853 19465 38887 19499
rect 44925 19465 44959 19499
rect 28089 19397 28123 19431
rect 32505 19397 32539 19431
rect 33977 19397 34011 19431
rect 43913 19397 43947 19431
rect 23949 19329 23983 19363
rect 24041 19329 24075 19363
rect 27353 19329 27387 19363
rect 29193 19329 29227 19363
rect 39037 19329 39071 19363
rect 42993 19329 43027 19363
rect 43085 19329 43119 19363
rect 45109 19329 45143 19363
rect 24133 19261 24167 19295
rect 29377 19261 29411 19295
rect 30021 19261 30055 19295
rect 30297 19261 30331 19295
rect 34069 19261 34103 19295
rect 35357 19261 35391 19295
rect 42073 19261 42107 19295
rect 43269 19261 43303 19295
rect 44097 19261 44131 19295
rect 33517 19193 33551 19227
rect 34713 19193 34747 19227
rect 31769 19125 31803 19159
rect 32597 19125 32631 19159
rect 42625 19125 42659 19159
rect 24593 18921 24627 18955
rect 27169 18921 27203 18955
rect 36737 18853 36771 18887
rect 25237 18785 25271 18819
rect 27721 18785 27755 18819
rect 30665 18785 30699 18819
rect 32597 18785 32631 18819
rect 32873 18785 32907 18819
rect 35357 18785 35391 18819
rect 35449 18785 35483 18819
rect 40969 18785 41003 18819
rect 41061 18785 41095 18819
rect 41705 18785 41739 18819
rect 41981 18785 42015 18819
rect 27629 18717 27663 18751
rect 28733 18717 28767 18751
rect 36277 18717 36311 18751
rect 36921 18717 36955 18751
rect 47961 18717 47995 18751
rect 49157 18717 49191 18751
rect 29929 18649 29963 18683
rect 24961 18581 24995 18615
rect 25053 18581 25087 18615
rect 27537 18581 27571 18615
rect 34345 18581 34379 18615
rect 34897 18581 34931 18615
rect 35265 18581 35299 18615
rect 36093 18581 36127 18615
rect 40509 18581 40543 18615
rect 40877 18581 40911 18615
rect 43453 18581 43487 18615
rect 23397 18377 23431 18411
rect 28641 18377 28675 18411
rect 35541 18377 35575 18411
rect 39681 18377 39715 18411
rect 44373 18377 44407 18411
rect 30297 18309 30331 18343
rect 35449 18309 35483 18343
rect 37749 18309 37783 18343
rect 42901 18309 42935 18343
rect 23765 18241 23799 18275
rect 23857 18241 23891 18275
rect 26617 18241 26651 18275
rect 27721 18241 27755 18275
rect 29009 18241 29043 18275
rect 29101 18241 29135 18275
rect 34437 18241 34471 18275
rect 39865 18241 39899 18275
rect 42625 18241 42659 18275
rect 45201 18241 45235 18275
rect 47961 18241 47995 18275
rect 24041 18173 24075 18207
rect 27813 18173 27847 18207
rect 27997 18173 28031 18207
rect 29193 18173 29227 18207
rect 30021 18173 30055 18207
rect 35633 18173 35667 18207
rect 37473 18173 37507 18207
rect 42073 18173 42107 18207
rect 49157 18173 49191 18207
rect 39221 18105 39255 18139
rect 45017 18105 45051 18139
rect 25605 18037 25639 18071
rect 27353 18037 27387 18071
rect 31769 18037 31803 18071
rect 34529 18037 34563 18071
rect 35081 18037 35115 18071
rect 37197 17833 37231 17867
rect 39221 17833 39255 17867
rect 34161 17765 34195 17799
rect 40325 17765 40359 17799
rect 25421 17697 25455 17731
rect 27445 17697 27479 17731
rect 28549 17697 28583 17731
rect 35449 17697 35483 17731
rect 28273 17629 28307 17663
rect 29929 17629 29963 17663
rect 33701 17629 33735 17663
rect 34345 17629 34379 17663
rect 39405 17629 39439 17663
rect 40509 17629 40543 17663
rect 41245 17629 41279 17663
rect 42901 17629 42935 17663
rect 44189 17629 44223 17663
rect 45293 17629 45327 17663
rect 25697 17561 25731 17595
rect 35725 17561 35759 17595
rect 44373 17561 44407 17595
rect 45477 17561 45511 17595
rect 27905 17493 27939 17527
rect 28365 17493 28399 17527
rect 41061 17493 41095 17527
rect 20361 17289 20395 17323
rect 25053 17289 25087 17323
rect 25421 17289 25455 17323
rect 27905 17289 27939 17323
rect 28273 17289 28307 17323
rect 29469 17289 29503 17323
rect 30389 17289 30423 17323
rect 32505 17289 32539 17323
rect 33057 17289 33091 17323
rect 33425 17289 33459 17323
rect 27445 17221 27479 17255
rect 32413 17221 32447 17255
rect 43085 17221 43119 17255
rect 44281 17221 44315 17255
rect 20729 17153 20763 17187
rect 30849 17153 30883 17187
rect 30941 17153 30975 17187
rect 37473 17153 37507 17187
rect 39681 17153 39715 17187
rect 42073 17153 42107 17187
rect 42993 17153 43027 17187
rect 44005 17153 44039 17187
rect 47961 17153 47995 17187
rect 19901 17085 19935 17119
rect 20821 17085 20855 17119
rect 20913 17085 20947 17119
rect 25513 17085 25547 17119
rect 25697 17085 25731 17119
rect 28365 17085 28399 17119
rect 28549 17085 28583 17119
rect 29561 17085 29595 17119
rect 29653 17085 29687 17119
rect 31033 17085 31067 17119
rect 33517 17085 33551 17119
rect 33609 17085 33643 17119
rect 37749 17085 37783 17119
rect 39221 17085 39255 17119
rect 39957 17085 39991 17119
rect 43269 17085 43303 17119
rect 49157 17085 49191 17119
rect 30481 17017 30515 17051
rect 42625 17017 42659 17051
rect 29101 16949 29135 16983
rect 31769 16949 31803 16983
rect 41429 16949 41463 16983
rect 45753 16949 45787 16983
rect 21005 16745 21039 16779
rect 22556 16745 22590 16779
rect 22293 16609 22327 16643
rect 25605 16609 25639 16643
rect 25697 16609 25731 16643
rect 27169 16609 27203 16643
rect 27353 16609 27387 16643
rect 28641 16609 28675 16643
rect 28825 16609 28859 16643
rect 29745 16609 29779 16643
rect 30021 16609 30055 16643
rect 31953 16609 31987 16643
rect 32229 16609 32263 16643
rect 36553 16609 36587 16643
rect 38485 16609 38519 16643
rect 38669 16609 38703 16643
rect 42717 16609 42751 16643
rect 42901 16609 42935 16643
rect 25513 16541 25547 16575
rect 28549 16541 28583 16575
rect 35541 16541 35575 16575
rect 36369 16541 36403 16575
rect 40233 16541 40267 16575
rect 47961 16541 47995 16575
rect 38393 16473 38427 16507
rect 42625 16473 42659 16507
rect 49157 16473 49191 16507
rect 24041 16405 24075 16439
rect 25145 16405 25179 16439
rect 26709 16405 26743 16439
rect 27077 16405 27111 16439
rect 28181 16405 28215 16439
rect 31493 16405 31527 16439
rect 33701 16405 33735 16439
rect 35357 16405 35391 16439
rect 38025 16405 38059 16439
rect 40049 16405 40083 16439
rect 42257 16405 42291 16439
rect 32689 16201 32723 16235
rect 35265 16201 35299 16235
rect 24777 16133 24811 16167
rect 33517 16065 33551 16099
rect 37657 16065 37691 16099
rect 38945 16065 38979 16099
rect 40785 16065 40819 16099
rect 24501 15997 24535 16031
rect 26525 15997 26559 16031
rect 28089 15997 28123 16031
rect 28365 15997 28399 16031
rect 30113 15997 30147 16031
rect 32781 15997 32815 16031
rect 32965 15997 32999 16031
rect 33793 15997 33827 16031
rect 32321 15861 32355 15895
rect 37473 15861 37507 15895
rect 38761 15861 38795 15895
rect 40601 15861 40635 15895
rect 23305 15657 23339 15691
rect 27813 15657 27847 15691
rect 31125 15657 31159 15691
rect 37381 15657 37415 15691
rect 37841 15589 37875 15623
rect 44465 15589 44499 15623
rect 23857 15521 23891 15555
rect 25237 15521 25271 15555
rect 28365 15521 28399 15555
rect 31677 15521 31711 15555
rect 35633 15521 35667 15555
rect 35909 15521 35943 15555
rect 38393 15521 38427 15555
rect 27261 15453 27295 15487
rect 30665 15453 30699 15487
rect 31493 15453 31527 15487
rect 32505 15453 32539 15487
rect 33609 15453 33643 15487
rect 38301 15453 38335 15487
rect 39129 15453 39163 15487
rect 47961 15453 47995 15487
rect 49157 15453 49191 15487
rect 23765 15385 23799 15419
rect 25513 15385 25547 15419
rect 28181 15385 28215 15419
rect 31585 15385 31619 15419
rect 44281 15385 44315 15419
rect 45569 15385 45603 15419
rect 45753 15385 45787 15419
rect 23673 15317 23707 15351
rect 28273 15317 28307 15351
rect 33701 15317 33735 15351
rect 38209 15317 38243 15351
rect 39221 15317 39255 15351
rect 25145 15113 25179 15147
rect 27813 15113 27847 15147
rect 29193 15113 29227 15147
rect 30481 15113 30515 15147
rect 37657 15113 37691 15147
rect 26433 15045 26467 15079
rect 35633 15045 35667 15079
rect 36369 15045 36403 15079
rect 39037 15045 39071 15079
rect 23397 14977 23431 15011
rect 25697 14977 25731 15011
rect 32321 14977 32355 15011
rect 34897 14977 34931 15011
rect 37841 14977 37875 15011
rect 38761 14977 38795 15011
rect 46029 14977 46063 15011
rect 47961 14977 47995 15011
rect 23673 14909 23707 14943
rect 29285 14909 29319 14943
rect 29377 14909 29411 14943
rect 30573 14909 30607 14943
rect 30757 14909 30791 14943
rect 32597 14909 32631 14943
rect 34069 14909 34103 14943
rect 49157 14909 49191 14943
rect 28825 14841 28859 14875
rect 30113 14841 30147 14875
rect 28273 14773 28307 14807
rect 36461 14773 36495 14807
rect 40509 14773 40543 14807
rect 45845 14773 45879 14807
rect 25605 14569 25639 14603
rect 28457 14569 28491 14603
rect 45661 14569 45695 14603
rect 35173 14501 35207 14535
rect 26157 14433 26191 14467
rect 27169 14433 27203 14467
rect 28181 14433 28215 14467
rect 29009 14433 29043 14467
rect 32137 14433 32171 14467
rect 35725 14433 35759 14467
rect 38117 14433 38151 14467
rect 39221 14433 39255 14467
rect 39405 14433 39439 14467
rect 25145 14365 25179 14399
rect 26985 14365 27019 14399
rect 27445 14365 27479 14399
rect 32045 14365 32079 14399
rect 35541 14365 35575 14399
rect 36553 14365 36587 14399
rect 40601 14365 40635 14399
rect 41245 14365 41279 14399
rect 45845 14365 45879 14399
rect 25973 14297 26007 14331
rect 30573 14297 30607 14331
rect 37289 14297 37323 14331
rect 26065 14229 26099 14263
rect 26617 14229 26651 14263
rect 27077 14229 27111 14263
rect 28825 14229 28859 14263
rect 28917 14229 28951 14263
rect 31033 14229 31067 14263
rect 31585 14229 31619 14263
rect 31953 14229 31987 14263
rect 35633 14229 35667 14263
rect 38761 14229 38795 14263
rect 39129 14229 39163 14263
rect 40417 14229 40451 14263
rect 41061 14229 41095 14263
rect 24593 14025 24627 14059
rect 25881 14025 25915 14059
rect 26249 14025 26283 14059
rect 26341 14025 26375 14059
rect 30297 14025 30331 14059
rect 30665 14025 30699 14059
rect 34621 14025 34655 14059
rect 37841 14025 37875 14059
rect 37933 14025 37967 14059
rect 43453 14025 43487 14059
rect 39313 13957 39347 13991
rect 45753 13957 45787 13991
rect 22845 13889 22879 13923
rect 27728 13889 27762 13923
rect 30757 13889 30791 13923
rect 31769 13889 31803 13923
rect 32873 13889 32907 13923
rect 35449 13889 35483 13923
rect 36461 13889 36495 13923
rect 39037 13889 39071 13923
rect 43361 13889 43395 13923
rect 47961 13889 47995 13923
rect 26525 13821 26559 13855
rect 30849 13821 30883 13855
rect 35541 13821 35575 13855
rect 35633 13821 35667 13855
rect 38117 13821 38151 13855
rect 45937 13821 45971 13855
rect 49157 13821 49191 13855
rect 35081 13753 35115 13787
rect 37473 13753 37507 13787
rect 20269 13685 20303 13719
rect 23108 13685 23142 13719
rect 27984 13685 28018 13719
rect 29469 13685 29503 13719
rect 33130 13685 33164 13719
rect 40785 13685 40819 13719
rect 19717 13481 19751 13515
rect 21005 13481 21039 13515
rect 22201 13481 22235 13515
rect 24961 13481 24995 13515
rect 26617 13481 26651 13515
rect 32781 13481 32815 13515
rect 38209 13481 38243 13515
rect 31769 13413 31803 13447
rect 42257 13413 42291 13447
rect 20361 13345 20395 13379
rect 21465 13345 21499 13379
rect 21649 13345 21683 13379
rect 25513 13345 25547 13379
rect 27169 13345 27203 13379
rect 28825 13345 28859 13379
rect 30849 13345 30883 13379
rect 30941 13345 30975 13379
rect 32413 13345 32447 13379
rect 33333 13345 33367 13379
rect 36461 13345 36495 13379
rect 44465 13345 44499 13379
rect 20085 13277 20119 13311
rect 21373 13277 21407 13311
rect 22569 13277 22603 13311
rect 28549 13277 28583 13311
rect 28641 13277 28675 13311
rect 30757 13277 30791 13311
rect 31585 13277 31619 13311
rect 32137 13277 32171 13311
rect 33149 13277 33183 13311
rect 35725 13277 35759 13311
rect 39497 13277 39531 13311
rect 40233 13277 40267 13311
rect 42441 13277 42475 13311
rect 44281 13277 44315 13311
rect 47961 13277 47995 13311
rect 20177 13209 20211 13243
rect 25329 13209 25363 13243
rect 33241 13209 33275 13243
rect 34989 13209 35023 13243
rect 35909 13209 35943 13243
rect 36737 13209 36771 13243
rect 49157 13209 49191 13243
rect 18613 13141 18647 13175
rect 25421 13141 25455 13175
rect 26985 13141 27019 13175
rect 27077 13141 27111 13175
rect 28181 13141 28215 13175
rect 30389 13141 30423 13175
rect 32229 13141 32263 13175
rect 35081 13141 35115 13175
rect 39313 13141 39347 13175
rect 40049 13141 40083 13175
rect 22937 12937 22971 12971
rect 27445 12937 27479 12971
rect 27813 12937 27847 12971
rect 32781 12937 32815 12971
rect 23305 12869 23339 12903
rect 27905 12869 27939 12903
rect 29193 12869 29227 12903
rect 35357 12869 35391 12903
rect 36093 12869 36127 12903
rect 37565 12869 37599 12903
rect 24133 12801 24167 12835
rect 29285 12801 29319 12835
rect 32689 12801 32723 12835
rect 36921 12801 36955 12835
rect 39221 12801 39255 12835
rect 41705 12801 41739 12835
rect 23397 12733 23431 12767
rect 23489 12733 23523 12767
rect 24409 12733 24443 12767
rect 27997 12733 28031 12767
rect 29377 12733 29411 12767
rect 30021 12733 30055 12767
rect 30297 12733 30331 12767
rect 32965 12733 32999 12767
rect 35541 12733 35575 12767
rect 39497 12733 39531 12767
rect 28825 12665 28859 12699
rect 36277 12665 36311 12699
rect 25881 12597 25915 12631
rect 31769 12597 31803 12631
rect 32321 12597 32355 12631
rect 33701 12597 33735 12631
rect 34805 12597 34839 12631
rect 36737 12597 36771 12631
rect 37657 12597 37691 12631
rect 40969 12597 41003 12631
rect 41521 12597 41555 12631
rect 24593 12393 24627 12427
rect 27261 12393 27295 12427
rect 29745 12393 29779 12427
rect 33149 12393 33183 12427
rect 38025 12393 38059 12427
rect 31953 12325 31987 12359
rect 25053 12257 25087 12291
rect 25145 12257 25179 12291
rect 27905 12257 27939 12291
rect 30297 12257 30331 12291
rect 32413 12257 32447 12291
rect 32505 12257 32539 12291
rect 33793 12257 33827 12291
rect 35357 12257 35391 12291
rect 35541 12257 35575 12291
rect 36277 12257 36311 12291
rect 26709 12189 26743 12223
rect 27629 12189 27663 12223
rect 27721 12189 27755 12223
rect 28641 12189 28675 12223
rect 30113 12189 30147 12223
rect 38669 12189 38703 12223
rect 39313 12189 39347 12223
rect 40233 12189 40267 12223
rect 47961 12189 47995 12223
rect 49157 12189 49191 12223
rect 32321 12121 32355 12155
rect 33517 12121 33551 12155
rect 35265 12121 35299 12155
rect 36553 12121 36587 12155
rect 24961 12053 24995 12087
rect 30205 12053 30239 12087
rect 33609 12053 33643 12087
rect 34897 12053 34931 12087
rect 38485 12053 38519 12087
rect 40049 12053 40083 12087
rect 25513 11849 25547 11883
rect 27169 11849 27203 11883
rect 28365 11849 28399 11883
rect 28733 11849 28767 11883
rect 29929 11849 29963 11883
rect 35265 11849 35299 11883
rect 36093 11849 36127 11883
rect 38209 11849 38243 11883
rect 40601 11849 40635 11883
rect 27537 11781 27571 11815
rect 38301 11781 38335 11815
rect 27629 11713 27663 11747
rect 30297 11713 30331 11747
rect 36277 11713 36311 11747
rect 39129 11713 39163 11747
rect 40509 11713 40543 11747
rect 41521 11713 41555 11747
rect 42809 11713 42843 11747
rect 44741 11713 44775 11747
rect 47961 11713 47995 11747
rect 23765 11645 23799 11679
rect 24041 11645 24075 11679
rect 27721 11645 27755 11679
rect 28825 11645 28859 11679
rect 29009 11645 29043 11679
rect 30389 11645 30423 11679
rect 30573 11645 30607 11679
rect 35357 11645 35391 11679
rect 35541 11645 35575 11679
rect 38485 11645 38519 11679
rect 39313 11645 39347 11679
rect 40693 11645 40727 11679
rect 49157 11645 49191 11679
rect 37841 11577 37875 11611
rect 40141 11577 40175 11611
rect 44557 11577 44591 11611
rect 34897 11509 34931 11543
rect 42625 11509 42659 11543
rect 27077 11305 27111 11339
rect 28181 11305 28215 11339
rect 29745 11305 29779 11339
rect 30941 11305 30975 11339
rect 32137 11305 32171 11339
rect 37657 11305 37691 11339
rect 34897 11237 34931 11271
rect 25329 11169 25363 11203
rect 25605 11169 25639 11203
rect 28733 11169 28767 11203
rect 30205 11169 30239 11203
rect 30297 11169 30331 11203
rect 31585 11169 31619 11203
rect 32781 11169 32815 11203
rect 35449 11169 35483 11203
rect 28549 11101 28583 11135
rect 31309 11101 31343 11135
rect 32505 11101 32539 11135
rect 33425 11101 33459 11135
rect 36277 11101 36311 11135
rect 37841 11101 37875 11135
rect 38669 11101 38703 11135
rect 27629 11033 27663 11067
rect 28641 11033 28675 11067
rect 30113 11033 30147 11067
rect 32597 11033 32631 11067
rect 34161 11033 34195 11067
rect 35265 11033 35299 11067
rect 35357 11033 35391 11067
rect 37013 11033 37047 11067
rect 38853 11033 38887 11067
rect 31401 10965 31435 10999
rect 28365 10761 28399 10795
rect 29561 10761 29595 10795
rect 29929 10761 29963 10795
rect 35633 10761 35667 10795
rect 32413 10693 32447 10727
rect 36093 10693 36127 10727
rect 28733 10625 28767 10659
rect 31125 10625 31159 10659
rect 36001 10625 36035 10659
rect 42809 10625 42843 10659
rect 47961 10625 47995 10659
rect 28825 10557 28859 10591
rect 28917 10557 28951 10591
rect 30021 10557 30055 10591
rect 30113 10557 30147 10591
rect 31217 10557 31251 10591
rect 31309 10557 31343 10591
rect 33149 10557 33183 10591
rect 33425 10557 33459 10591
rect 36277 10557 36311 10591
rect 38945 10557 38979 10591
rect 39221 10557 39255 10591
rect 49157 10557 49191 10591
rect 34897 10489 34931 10523
rect 30757 10421 30791 10455
rect 32505 10421 32539 10455
rect 40693 10421 40727 10455
rect 42625 10421 42659 10455
rect 32413 10217 32447 10251
rect 32873 10217 32907 10251
rect 37105 10217 37139 10251
rect 25789 10081 25823 10115
rect 26065 10081 26099 10115
rect 30665 10081 30699 10115
rect 33425 10081 33459 10115
rect 35357 10013 35391 10047
rect 37749 10013 37783 10047
rect 38761 10013 38795 10047
rect 46857 10013 46891 10047
rect 47961 10013 47995 10047
rect 30941 9945 30975 9979
rect 35633 9945 35667 9979
rect 46121 9945 46155 9979
rect 46305 9945 46339 9979
rect 47041 9945 47075 9979
rect 49157 9945 49191 9979
rect 27537 9877 27571 9911
rect 33241 9877 33275 9911
rect 33333 9877 33367 9911
rect 38577 9877 38611 9911
rect 29653 9605 29687 9639
rect 30849 9605 30883 9639
rect 36185 9605 36219 9639
rect 38761 9605 38795 9639
rect 29745 9537 29779 9571
rect 33149 9537 33183 9571
rect 34989 9537 35023 9571
rect 35081 9537 35115 9571
rect 38485 9537 38519 9571
rect 43729 9537 43763 9571
rect 46489 9537 46523 9571
rect 29929 9469 29963 9503
rect 30941 9469 30975 9503
rect 31033 9469 31067 9503
rect 33241 9469 33275 9503
rect 33425 9469 33459 9503
rect 35265 9469 35299 9503
rect 29285 9401 29319 9435
rect 30481 9401 30515 9435
rect 23305 9333 23339 9367
rect 26433 9333 26467 9367
rect 28825 9333 28859 9367
rect 32781 9333 32815 9367
rect 34621 9333 34655 9367
rect 36277 9333 36311 9367
rect 37657 9333 37691 9367
rect 40233 9333 40267 9367
rect 43545 9333 43579 9367
rect 46305 9333 46339 9367
rect 22753 9129 22787 9163
rect 45385 9129 45419 9163
rect 45937 9129 45971 9163
rect 27077 9061 27111 9095
rect 28457 9061 28491 9095
rect 31953 9061 31987 9095
rect 37105 9061 37139 9095
rect 38301 9061 38335 9095
rect 41245 9061 41279 9095
rect 23397 8993 23431 9027
rect 25605 8993 25639 9027
rect 29009 8993 29043 9027
rect 29745 8993 29779 9027
rect 30021 8993 30055 9027
rect 32413 8993 32447 9027
rect 32597 8993 32631 9027
rect 37565 8993 37599 9027
rect 37657 8993 37691 9027
rect 38853 8993 38887 9027
rect 22293 8925 22327 8959
rect 23213 8925 23247 8959
rect 25329 8925 25363 8959
rect 28825 8925 28859 8959
rect 33241 8925 33275 8959
rect 34897 8925 34931 8959
rect 38669 8925 38703 8959
rect 38761 8925 38795 8959
rect 40233 8925 40267 8959
rect 41429 8925 41463 8959
rect 46121 8925 46155 8959
rect 46857 8925 46891 8959
rect 47961 8925 47995 8959
rect 23121 8857 23155 8891
rect 28917 8857 28951 8891
rect 35173 8857 35207 8891
rect 37473 8857 37507 8891
rect 45293 8857 45327 8891
rect 49157 8857 49191 8891
rect 31493 8789 31527 8823
rect 32321 8789 32355 8823
rect 33333 8789 33367 8823
rect 36645 8789 36679 8823
rect 46673 8789 46707 8823
rect 23489 8585 23523 8619
rect 23949 8585 23983 8619
rect 24685 8585 24719 8619
rect 30941 8585 30975 8619
rect 32321 8585 32355 8619
rect 32689 8585 32723 8619
rect 35817 8585 35851 8619
rect 39497 8585 39531 8619
rect 40325 8585 40359 8619
rect 25053 8517 25087 8551
rect 25145 8517 25179 8551
rect 31401 8517 31435 8551
rect 34345 8517 34379 8551
rect 36737 8517 36771 8551
rect 40417 8517 40451 8551
rect 46673 8517 46707 8551
rect 23029 8449 23063 8483
rect 23857 8449 23891 8483
rect 25881 8449 25915 8483
rect 26433 8449 26467 8483
rect 31309 8449 31343 8483
rect 34069 8449 34103 8483
rect 47961 8449 47995 8483
rect 24133 8381 24167 8415
rect 25329 8381 25363 8415
rect 26525 8381 26559 8415
rect 26709 8381 26743 8415
rect 27636 8381 27670 8415
rect 29377 8381 29411 8415
rect 31493 8381 31527 8415
rect 32781 8381 32815 8415
rect 32873 8381 32907 8415
rect 37749 8381 37783 8415
rect 38025 8381 38059 8415
rect 40509 8381 40543 8415
rect 49157 8381 49191 8415
rect 36921 8313 36955 8347
rect 39957 8313 39991 8347
rect 46857 8313 46891 8347
rect 26065 8245 26099 8279
rect 27886 8245 27920 8279
rect 27813 8041 27847 8075
rect 32321 8041 32355 8075
rect 37565 8041 37599 8075
rect 40049 8041 40083 8075
rect 28273 7973 28307 8007
rect 38393 7973 38427 8007
rect 26065 7905 26099 7939
rect 26341 7905 26375 7939
rect 28733 7905 28767 7939
rect 28917 7905 28951 7939
rect 31585 7905 31619 7939
rect 36093 7905 36127 7939
rect 31309 7837 31343 7871
rect 31401 7837 31435 7871
rect 32965 7837 32999 7871
rect 35265 7837 35299 7871
rect 35817 7837 35851 7871
rect 38577 7837 38611 7871
rect 40233 7837 40267 7871
rect 28641 7701 28675 7735
rect 30941 7701 30975 7735
rect 28641 7429 28675 7463
rect 32505 7429 32539 7463
rect 35725 7429 35759 7463
rect 33149 7361 33183 7395
rect 35817 7361 35851 7395
rect 43269 7361 43303 7395
rect 47133 7361 47167 7395
rect 47961 7361 47995 7395
rect 33425 7293 33459 7327
rect 34897 7293 34931 7327
rect 35909 7293 35943 7327
rect 49157 7293 49191 7327
rect 28825 7225 28859 7259
rect 35357 7225 35391 7259
rect 32597 7157 32631 7191
rect 38485 7157 38519 7191
rect 43085 7157 43119 7191
rect 46949 7157 46983 7191
rect 30008 6953 30042 6987
rect 36718 6953 36752 6987
rect 29745 6817 29779 6851
rect 31953 6817 31987 6851
rect 36461 6817 36495 6851
rect 38209 6817 38243 6851
rect 39221 6817 39255 6851
rect 34989 6749 35023 6783
rect 35173 6749 35207 6783
rect 39037 6749 39071 6783
rect 39129 6749 39163 6783
rect 41705 6749 41739 6783
rect 47961 6749 47995 6783
rect 32229 6681 32263 6715
rect 35817 6681 35851 6715
rect 49157 6681 49191 6715
rect 31493 6613 31527 6647
rect 33701 6613 33735 6647
rect 35909 6613 35943 6647
rect 38669 6613 38703 6647
rect 41521 6613 41555 6647
rect 34069 6409 34103 6443
rect 32597 6341 32631 6375
rect 37565 6341 37599 6375
rect 38301 6341 38335 6375
rect 39497 6341 39531 6375
rect 32321 6273 32355 6307
rect 47961 6273 47995 6307
rect 37749 6205 37783 6239
rect 49157 6205 49191 6239
rect 38485 6137 38519 6171
rect 39589 6069 39623 6103
rect 32045 5865 32079 5899
rect 39037 5865 39071 5899
rect 45201 5865 45235 5899
rect 40325 5797 40359 5831
rect 32597 5729 32631 5763
rect 38393 5729 38427 5763
rect 29837 5661 29871 5695
rect 32413 5661 32447 5695
rect 38209 5661 38243 5695
rect 42257 5661 42291 5695
rect 45385 5661 45419 5695
rect 46857 5661 46891 5695
rect 47961 5661 47995 5695
rect 32505 5593 32539 5627
rect 38945 5593 38979 5627
rect 40141 5593 40175 5627
rect 40877 5593 40911 5627
rect 41061 5593 41095 5627
rect 47041 5593 47075 5627
rect 49157 5593 49191 5627
rect 29929 5525 29963 5559
rect 42073 5525 42107 5559
rect 39957 5253 39991 5287
rect 40877 5253 40911 5287
rect 46213 5185 46247 5219
rect 47961 5185 47995 5219
rect 40141 5117 40175 5151
rect 49157 5117 49191 5151
rect 41061 5049 41095 5083
rect 46029 4981 46063 5015
rect 11437 4641 11471 4675
rect 48421 4641 48455 4675
rect 46121 4573 46155 4607
rect 47961 4573 47995 4607
rect 11713 4505 11747 4539
rect 13461 4505 13495 4539
rect 47317 4505 47351 4539
rect 34161 4097 34195 4131
rect 39129 4097 39163 4131
rect 44281 4097 44315 4131
rect 46489 4097 46523 4131
rect 47961 4097 47995 4131
rect 34437 4029 34471 4063
rect 39589 4029 39623 4063
rect 44741 4029 44775 4063
rect 49157 4029 49191 4063
rect 46305 3893 46339 3927
rect 48513 3689 48547 3723
rect 20269 3553 20303 3587
rect 25053 3553 25087 3587
rect 30205 3553 30239 3587
rect 32045 3553 32079 3587
rect 35357 3553 35391 3587
rect 37197 3553 37231 3587
rect 40509 3553 40543 3587
rect 42349 3553 42383 3587
rect 45661 3553 45695 3587
rect 17233 3485 17267 3519
rect 19993 3485 20027 3519
rect 24685 3485 24719 3519
rect 29929 3485 29963 3519
rect 31677 3485 31711 3519
rect 34897 3485 34931 3519
rect 36921 3485 36955 3519
rect 40049 3485 40083 3519
rect 41889 3485 41923 3519
rect 45201 3485 45235 3519
rect 47225 3417 47259 3451
rect 17049 3349 17083 3383
rect 3985 3145 4019 3179
rect 6745 3145 6779 3179
rect 11713 3145 11747 3179
rect 49157 3077 49191 3111
rect 2605 3009 2639 3043
rect 3893 3009 3927 3043
rect 6929 3009 6963 3043
rect 9045 3009 9079 3043
rect 11897 3009 11931 3043
rect 12909 3009 12943 3043
rect 14381 3009 14415 3043
rect 18061 3009 18095 3043
rect 22477 3009 22511 3043
rect 25329 3009 25363 3043
rect 27537 3009 27571 3043
rect 29377 3009 29411 3043
rect 32505 3009 32539 3043
rect 34345 3009 34379 3043
rect 37657 3009 37691 3043
rect 39497 3009 39531 3043
rect 42625 3009 42659 3043
rect 44465 3009 44499 3043
rect 47961 3009 47995 3043
rect 2329 2941 2363 2975
rect 12633 2941 12667 2975
rect 14105 2941 14139 2975
rect 17785 2941 17819 2975
rect 19257 2941 19291 2975
rect 19533 2941 19567 2975
rect 20637 2941 20671 2975
rect 20913 2941 20947 2975
rect 22201 2941 22235 2975
rect 25605 2941 25639 2975
rect 27813 2941 27847 2975
rect 29653 2941 29687 2975
rect 32781 2941 32815 2975
rect 34621 2941 34655 2975
rect 37933 2941 37967 2975
rect 39773 2941 39807 2975
rect 43085 2941 43119 2975
rect 44925 2941 44959 2975
rect 9229 2873 9263 2907
rect 1593 2601 1627 2635
rect 15071 2601 15105 2635
rect 22569 2533 22603 2567
rect 2881 2465 2915 2499
rect 10609 2465 10643 2499
rect 12909 2465 12943 2499
rect 18061 2465 18095 2499
rect 25789 2465 25823 2499
rect 27629 2465 27663 2499
rect 30389 2465 30423 2499
rect 32781 2465 32815 2499
rect 37933 2465 37967 2499
rect 43085 2465 43119 2499
rect 45661 2465 45695 2499
rect 48329 2465 48363 2499
rect 1777 2397 1811 2431
rect 2605 2397 2639 2431
rect 7665 2397 7699 2431
rect 8493 2397 8527 2431
rect 10333 2397 10367 2431
rect 12081 2397 12115 2431
rect 13185 2397 13219 2431
rect 14841 2397 14875 2431
rect 16313 2397 16347 2431
rect 17049 2397 17083 2431
rect 22753 2397 22787 2431
rect 23213 2397 23247 2431
rect 25237 2397 25271 2431
rect 27353 2397 27387 2431
rect 29745 2397 29779 2431
rect 32505 2397 32539 2431
rect 35081 2397 35115 2431
rect 37473 2397 37507 2431
rect 40141 2397 40175 2431
rect 42625 2397 42659 2431
rect 45201 2397 45235 2431
rect 47777 2397 47811 2431
rect 4629 2329 4663 2363
rect 5365 2329 5399 2363
rect 5549 2329 5583 2363
rect 6653 2329 6687 2363
rect 8309 2329 8343 2363
rect 9689 2329 9723 2363
rect 9873 2329 9907 2363
rect 21281 2329 21315 2363
rect 21465 2329 21499 2363
rect 35817 2329 35851 2363
rect 40969 2329 41003 2363
rect 4721 2261 4755 2295
rect 6745 2261 6779 2295
rect 7481 2261 7515 2295
rect 11897 2261 11931 2295
rect 16129 2261 16163 2295
rect 16865 2261 16899 2295
rect 18291 2261 18325 2295
rect 23443 2261 23477 2295
<< metal1 >>
rect 1104 54426 49864 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 27950 54426
rect 28002 54374 28014 54426
rect 28066 54374 28078 54426
rect 28130 54374 28142 54426
rect 28194 54374 28206 54426
rect 28258 54374 37950 54426
rect 38002 54374 38014 54426
rect 38066 54374 38078 54426
rect 38130 54374 38142 54426
rect 38194 54374 38206 54426
rect 38258 54374 47950 54426
rect 48002 54374 48014 54426
rect 48066 54374 48078 54426
rect 48130 54374 48142 54426
rect 48194 54374 48206 54426
rect 48258 54374 49864 54426
rect 1104 54352 49864 54374
rect 29546 54272 29552 54324
rect 29604 54312 29610 54324
rect 33505 54315 33563 54321
rect 33505 54312 33517 54315
rect 29604 54284 33517 54312
rect 29604 54272 29610 54284
rect 33505 54281 33517 54284
rect 33551 54281 33563 54315
rect 33505 54275 33563 54281
rect 8386 54244 8392 54256
rect 4356 54216 8392 54244
rect 4356 54185 4384 54216
rect 8386 54204 8392 54216
rect 8444 54204 8450 54256
rect 36078 54204 36084 54256
rect 36136 54244 36142 54256
rect 36265 54247 36323 54253
rect 36265 54244 36277 54247
rect 36136 54216 36277 54244
rect 36136 54204 36142 54216
rect 36265 54213 36277 54216
rect 36311 54213 36323 54247
rect 36265 54207 36323 54213
rect 46750 54204 46756 54256
rect 46808 54244 46814 54256
rect 46845 54247 46903 54253
rect 46845 54244 46857 54247
rect 46808 54216 46857 54244
rect 46808 54204 46814 54216
rect 46845 54213 46857 54216
rect 46891 54213 46903 54247
rect 46845 54207 46903 54213
rect 1765 54179 1823 54185
rect 1765 54145 1777 54179
rect 1811 54176 1823 54179
rect 4341 54179 4399 54185
rect 1811 54148 4016 54176
rect 1811 54145 1823 54148
rect 1765 54139 1823 54145
rect 1394 54068 1400 54120
rect 1452 54108 1458 54120
rect 2041 54111 2099 54117
rect 2041 54108 2053 54111
rect 1452 54080 2053 54108
rect 1452 54068 1458 54080
rect 2041 54077 2053 54080
rect 2087 54077 2099 54111
rect 2041 54071 2099 54077
rect 3988 54040 4016 54148
rect 4341 54145 4353 54179
rect 4387 54145 4399 54179
rect 4341 54139 4399 54145
rect 6917 54179 6975 54185
rect 6917 54145 6929 54179
rect 6963 54176 6975 54179
rect 7098 54176 7104 54188
rect 6963 54148 7104 54176
rect 6963 54145 6975 54148
rect 6917 54139 6975 54145
rect 7098 54136 7104 54148
rect 7156 54136 7162 54188
rect 9582 54136 9588 54188
rect 9640 54136 9646 54188
rect 12250 54136 12256 54188
rect 12308 54136 12314 54188
rect 15010 54136 15016 54188
rect 15068 54136 15074 54188
rect 17678 54136 17684 54188
rect 17736 54136 17742 54188
rect 20254 54136 20260 54188
rect 20312 54136 20318 54188
rect 22830 54136 22836 54188
rect 22888 54136 22894 54188
rect 25406 54136 25412 54188
rect 25464 54176 25470 54188
rect 25685 54179 25743 54185
rect 25685 54176 25697 54179
rect 25464 54148 25697 54176
rect 25464 54136 25470 54148
rect 25685 54145 25697 54148
rect 25731 54145 25743 54179
rect 25685 54139 25743 54145
rect 28350 54136 28356 54188
rect 28408 54136 28414 54188
rect 30742 54136 30748 54188
rect 30800 54176 30806 54188
rect 31021 54179 31079 54185
rect 31021 54176 31033 54179
rect 30800 54148 31033 54176
rect 30800 54136 30806 54148
rect 31021 54145 31033 54148
rect 31067 54145 31079 54179
rect 31021 54139 31079 54145
rect 33410 54136 33416 54188
rect 33468 54176 33474 54188
rect 33689 54179 33747 54185
rect 33689 54176 33701 54179
rect 33468 54148 33701 54176
rect 33468 54136 33474 54148
rect 33689 54145 33701 54148
rect 33735 54145 33747 54179
rect 33689 54139 33747 54145
rect 38746 54136 38752 54188
rect 38804 54176 38810 54188
rect 38841 54179 38899 54185
rect 38841 54176 38853 54179
rect 38804 54148 38853 54176
rect 38804 54136 38810 54148
rect 38841 54145 38853 54148
rect 38887 54145 38899 54179
rect 38841 54139 38899 54145
rect 41414 54136 41420 54188
rect 41472 54176 41478 54188
rect 41509 54179 41567 54185
rect 41509 54176 41521 54179
rect 41472 54148 41521 54176
rect 41472 54136 41478 54148
rect 41509 54145 41521 54148
rect 41555 54145 41567 54179
rect 41509 54139 41567 54145
rect 44082 54136 44088 54188
rect 44140 54176 44146 54188
rect 44177 54179 44235 54185
rect 44177 54176 44189 54179
rect 44140 54148 44189 54176
rect 44140 54136 44146 54148
rect 44177 54145 44189 54148
rect 44223 54145 44235 54179
rect 44177 54139 44235 54145
rect 48314 54136 48320 54188
rect 48372 54136 48378 54188
rect 49050 54136 49056 54188
rect 49108 54136 49114 54188
rect 4062 54068 4068 54120
rect 4120 54108 4126 54120
rect 4617 54111 4675 54117
rect 4617 54108 4629 54111
rect 4120 54080 4629 54108
rect 4120 54068 4126 54080
rect 4617 54077 4629 54080
rect 4663 54077 4675 54111
rect 4617 54071 4675 54077
rect 7006 54068 7012 54120
rect 7064 54108 7070 54120
rect 7285 54111 7343 54117
rect 7285 54108 7297 54111
rect 7064 54080 7297 54108
rect 7064 54068 7070 54080
rect 7285 54077 7297 54080
rect 7331 54077 7343 54111
rect 7285 54071 7343 54077
rect 9398 54068 9404 54120
rect 9456 54108 9462 54120
rect 9953 54111 10011 54117
rect 9953 54108 9965 54111
rect 9456 54080 9965 54108
rect 9456 54068 9462 54080
rect 9953 54077 9965 54080
rect 9999 54077 10011 54111
rect 9953 54071 10011 54077
rect 12342 54068 12348 54120
rect 12400 54108 12406 54120
rect 12621 54111 12679 54117
rect 12621 54108 12633 54111
rect 12400 54080 12633 54108
rect 12400 54068 12406 54080
rect 12621 54077 12633 54080
rect 12667 54077 12679 54111
rect 12621 54071 12679 54077
rect 14734 54068 14740 54120
rect 14792 54108 14798 54120
rect 15289 54111 15347 54117
rect 15289 54108 15301 54111
rect 14792 54080 15301 54108
rect 14792 54068 14798 54080
rect 15289 54077 15301 54080
rect 15335 54077 15347 54111
rect 15289 54071 15347 54077
rect 17862 54068 17868 54120
rect 17920 54108 17926 54120
rect 17957 54111 18015 54117
rect 17957 54108 17969 54111
rect 17920 54080 17969 54108
rect 17920 54068 17926 54080
rect 17957 54077 17969 54080
rect 18003 54077 18015 54111
rect 17957 54071 18015 54077
rect 20162 54068 20168 54120
rect 20220 54108 20226 54120
rect 20533 54111 20591 54117
rect 20533 54108 20545 54111
rect 20220 54080 20545 54108
rect 20220 54068 20226 54080
rect 20533 54077 20545 54080
rect 20579 54077 20591 54111
rect 20533 54071 20591 54077
rect 22738 54068 22744 54120
rect 22796 54108 22802 54120
rect 23109 54111 23167 54117
rect 23109 54108 23121 54111
rect 22796 54080 23121 54108
rect 22796 54068 22802 54080
rect 23109 54077 23121 54080
rect 23155 54077 23167 54111
rect 23109 54071 23167 54077
rect 15194 54040 15200 54052
rect 3988 54012 15200 54040
rect 15194 54000 15200 54012
rect 15252 54000 15258 54052
rect 36449 54043 36507 54049
rect 36449 54040 36461 54043
rect 20548 54012 36461 54040
rect 20548 53984 20576 54012
rect 36449 54009 36461 54012
rect 36495 54009 36507 54043
rect 36449 54003 36507 54009
rect 20530 53932 20536 53984
rect 20588 53932 20594 53984
rect 24394 53932 24400 53984
rect 24452 53972 24458 53984
rect 25501 53975 25559 53981
rect 25501 53972 25513 53975
rect 24452 53944 25513 53972
rect 24452 53932 24458 53944
rect 25501 53941 25513 53944
rect 25547 53941 25559 53975
rect 25501 53935 25559 53941
rect 25682 53932 25688 53984
rect 25740 53972 25746 53984
rect 28169 53975 28227 53981
rect 28169 53972 28181 53975
rect 25740 53944 28181 53972
rect 25740 53932 25746 53944
rect 28169 53941 28181 53944
rect 28215 53941 28227 53975
rect 28169 53935 28227 53941
rect 30834 53932 30840 53984
rect 30892 53932 30898 53984
rect 39022 53932 39028 53984
rect 39080 53932 39086 53984
rect 41690 53932 41696 53984
rect 41748 53932 41754 53984
rect 44358 53932 44364 53984
rect 44416 53932 44422 53984
rect 46934 53932 46940 53984
rect 46992 53932 46998 53984
rect 48498 53932 48504 53984
rect 48556 53932 48562 53984
rect 48866 53932 48872 53984
rect 48924 53972 48930 53984
rect 49237 53975 49295 53981
rect 49237 53972 49249 53975
rect 48924 53944 49249 53972
rect 48924 53932 48930 53944
rect 49237 53941 49249 53944
rect 49283 53941 49295 53975
rect 49237 53935 49295 53941
rect 1104 53882 49864 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 32950 53882
rect 33002 53830 33014 53882
rect 33066 53830 33078 53882
rect 33130 53830 33142 53882
rect 33194 53830 33206 53882
rect 33258 53830 42950 53882
rect 43002 53830 43014 53882
rect 43066 53830 43078 53882
rect 43130 53830 43142 53882
rect 43194 53830 43206 53882
rect 43258 53830 49864 53882
rect 1104 53808 49864 53830
rect 49418 53632 49424 53644
rect 47872 53604 49424 53632
rect 47872 53573 47900 53604
rect 49418 53592 49424 53604
rect 49476 53592 49482 53644
rect 47857 53567 47915 53573
rect 47857 53533 47869 53567
rect 47903 53533 47915 53567
rect 47857 53527 47915 53533
rect 48317 53567 48375 53573
rect 48317 53533 48329 53567
rect 48363 53564 48375 53567
rect 48406 53564 48412 53576
rect 48363 53536 48412 53564
rect 48363 53533 48375 53536
rect 48317 53527 48375 53533
rect 48406 53524 48412 53536
rect 48464 53524 48470 53576
rect 49053 53567 49111 53573
rect 49053 53533 49065 53567
rect 49099 53564 49111 53567
rect 49142 53564 49148 53576
rect 49099 53536 49148 53564
rect 49099 53533 49111 53536
rect 49053 53527 49111 53533
rect 49142 53524 49148 53536
rect 49200 53524 49206 53576
rect 43438 53388 43444 53440
rect 43496 53428 43502 53440
rect 47673 53431 47731 53437
rect 47673 53428 47685 53431
rect 43496 53400 47685 53428
rect 43496 53388 43502 53400
rect 47673 53397 47685 53400
rect 47719 53397 47731 53431
rect 47673 53391 47731 53397
rect 48406 53388 48412 53440
rect 48464 53428 48470 53440
rect 48501 53431 48559 53437
rect 48501 53428 48513 53431
rect 48464 53400 48513 53428
rect 48464 53388 48470 53400
rect 48501 53397 48513 53400
rect 48547 53397 48559 53431
rect 48501 53391 48559 53397
rect 49237 53431 49295 53437
rect 49237 53397 49249 53431
rect 49283 53428 49295 53431
rect 50154 53428 50160 53440
rect 49283 53400 50160 53428
rect 49283 53397 49295 53400
rect 49237 53391 49295 53397
rect 50154 53388 50160 53400
rect 50212 53388 50218 53440
rect 1104 53338 49864 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 27950 53338
rect 28002 53286 28014 53338
rect 28066 53286 28078 53338
rect 28130 53286 28142 53338
rect 28194 53286 28206 53338
rect 28258 53286 37950 53338
rect 38002 53286 38014 53338
rect 38066 53286 38078 53338
rect 38130 53286 38142 53338
rect 38194 53286 38206 53338
rect 38258 53286 47950 53338
rect 48002 53286 48014 53338
rect 48066 53286 48078 53338
rect 48130 53286 48142 53338
rect 48194 53286 48206 53338
rect 48258 53286 49864 53338
rect 1104 53264 49864 53286
rect 8386 53184 8392 53236
rect 8444 53224 8450 53236
rect 9861 53227 9919 53233
rect 9861 53224 9873 53227
rect 8444 53196 9873 53224
rect 8444 53184 8450 53196
rect 9861 53193 9873 53196
rect 9907 53193 9919 53227
rect 9861 53187 9919 53193
rect 9769 53091 9827 53097
rect 9769 53057 9781 53091
rect 9815 53088 9827 53091
rect 13722 53088 13728 53100
rect 9815 53060 13728 53088
rect 9815 53057 9827 53060
rect 9769 53051 9827 53057
rect 13722 53048 13728 53060
rect 13780 53048 13786 53100
rect 49050 53048 49056 53100
rect 49108 53048 49114 53100
rect 34698 52844 34704 52896
rect 34756 52884 34762 52896
rect 49237 52887 49295 52893
rect 49237 52884 49249 52887
rect 34756 52856 49249 52884
rect 34756 52844 34762 52856
rect 49237 52853 49249 52856
rect 49283 52853 49295 52887
rect 49237 52847 49295 52853
rect 1104 52794 49864 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 32950 52794
rect 33002 52742 33014 52794
rect 33066 52742 33078 52794
rect 33130 52742 33142 52794
rect 33194 52742 33206 52794
rect 33258 52742 42950 52794
rect 43002 52742 43014 52794
rect 43066 52742 43078 52794
rect 43130 52742 43142 52794
rect 43194 52742 43206 52794
rect 43258 52742 49864 52794
rect 1104 52720 49864 52742
rect 49329 52479 49387 52485
rect 49329 52445 49341 52479
rect 49375 52476 49387 52479
rect 49970 52476 49976 52488
rect 49375 52448 49976 52476
rect 49375 52445 49387 52448
rect 49329 52439 49387 52445
rect 49970 52436 49976 52448
rect 50028 52436 50034 52488
rect 48958 52368 48964 52420
rect 49016 52368 49022 52420
rect 1104 52250 49864 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 27950 52250
rect 28002 52198 28014 52250
rect 28066 52198 28078 52250
rect 28130 52198 28142 52250
rect 28194 52198 28206 52250
rect 28258 52198 37950 52250
rect 38002 52198 38014 52250
rect 38066 52198 38078 52250
rect 38130 52198 38142 52250
rect 38194 52198 38206 52250
rect 38258 52198 47950 52250
rect 48002 52198 48014 52250
rect 48066 52198 48078 52250
rect 48130 52198 48142 52250
rect 48194 52198 48206 52250
rect 48258 52198 49864 52250
rect 1104 52176 49864 52198
rect 7098 52096 7104 52148
rect 7156 52136 7162 52148
rect 12805 52139 12863 52145
rect 12805 52136 12817 52139
rect 7156 52108 12817 52136
rect 7156 52096 7162 52108
rect 12805 52105 12817 52108
rect 12851 52105 12863 52139
rect 12805 52099 12863 52105
rect 12713 52003 12771 52009
rect 12713 51969 12725 52003
rect 12759 52000 12771 52003
rect 19794 52000 19800 52012
rect 12759 51972 19800 52000
rect 12759 51969 12771 51972
rect 12713 51963 12771 51969
rect 19794 51960 19800 51972
rect 19852 51960 19858 52012
rect 1104 51706 49864 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 32950 51706
rect 33002 51654 33014 51706
rect 33066 51654 33078 51706
rect 33130 51654 33142 51706
rect 33194 51654 33206 51706
rect 33258 51654 42950 51706
rect 43002 51654 43014 51706
rect 43066 51654 43078 51706
rect 43130 51654 43142 51706
rect 43194 51654 43206 51706
rect 43258 51654 49864 51706
rect 1104 51632 49864 51654
rect 15010 51552 15016 51604
rect 15068 51592 15074 51604
rect 16301 51595 16359 51601
rect 16301 51592 16313 51595
rect 15068 51564 16313 51592
rect 15068 51552 15074 51564
rect 16301 51561 16313 51564
rect 16347 51561 16359 51595
rect 16301 51555 16359 51561
rect 12250 51484 12256 51536
rect 12308 51524 12314 51536
rect 17313 51527 17371 51533
rect 17313 51524 17325 51527
rect 12308 51496 17325 51524
rect 12308 51484 12314 51496
rect 17313 51493 17325 51496
rect 17359 51493 17371 51527
rect 17313 51487 17371 51493
rect 21634 51456 21640 51468
rect 14936 51428 21640 51456
rect 14936 51397 14964 51428
rect 21634 51416 21640 51428
rect 21692 51416 21698 51468
rect 14921 51391 14979 51397
rect 14921 51357 14933 51391
rect 14967 51357 14979 51391
rect 14921 51351 14979 51357
rect 16485 51391 16543 51397
rect 16485 51357 16497 51391
rect 16531 51388 16543 51391
rect 17494 51388 17500 51400
rect 16531 51360 17500 51388
rect 16531 51357 16543 51360
rect 16485 51351 16543 51357
rect 17494 51348 17500 51360
rect 17552 51348 17558 51400
rect 17129 51323 17187 51329
rect 17129 51289 17141 51323
rect 17175 51320 17187 51323
rect 22738 51320 22744 51332
rect 17175 51292 22744 51320
rect 17175 51289 17187 51292
rect 17129 51283 17187 51289
rect 22738 51280 22744 51292
rect 22796 51280 22802 51332
rect 48958 51280 48964 51332
rect 49016 51280 49022 51332
rect 49329 51323 49387 51329
rect 49329 51289 49341 51323
rect 49375 51320 49387 51323
rect 49602 51320 49608 51332
rect 49375 51292 49608 51320
rect 49375 51289 49387 51292
rect 49329 51283 49387 51289
rect 49602 51280 49608 51292
rect 49660 51280 49666 51332
rect 9582 51212 9588 51264
rect 9640 51252 9646 51264
rect 15013 51255 15071 51261
rect 15013 51252 15025 51255
rect 9640 51224 15025 51252
rect 9640 51212 9646 51224
rect 15013 51221 15025 51224
rect 15059 51221 15071 51255
rect 15013 51215 15071 51221
rect 1104 51162 49864 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 27950 51162
rect 28002 51110 28014 51162
rect 28066 51110 28078 51162
rect 28130 51110 28142 51162
rect 28194 51110 28206 51162
rect 28258 51110 37950 51162
rect 38002 51110 38014 51162
rect 38066 51110 38078 51162
rect 38130 51110 38142 51162
rect 38194 51110 38206 51162
rect 38258 51110 47950 51162
rect 48002 51110 48014 51162
rect 48066 51110 48078 51162
rect 48130 51110 48142 51162
rect 48194 51110 48206 51162
rect 48258 51110 49864 51162
rect 1104 51088 49864 51110
rect 48958 50872 48964 50924
rect 49016 50872 49022 50924
rect 35710 50668 35716 50720
rect 35768 50708 35774 50720
rect 49053 50711 49111 50717
rect 49053 50708 49065 50711
rect 35768 50680 49065 50708
rect 35768 50668 35774 50680
rect 49053 50677 49065 50680
rect 49099 50677 49111 50711
rect 49053 50671 49111 50677
rect 1104 50618 49864 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 32950 50618
rect 33002 50566 33014 50618
rect 33066 50566 33078 50618
rect 33130 50566 33142 50618
rect 33194 50566 33206 50618
rect 33258 50566 42950 50618
rect 43002 50566 43014 50618
rect 43066 50566 43078 50618
rect 43130 50566 43142 50618
rect 43194 50566 43206 50618
rect 43258 50566 49864 50618
rect 1104 50544 49864 50566
rect 15194 50464 15200 50516
rect 15252 50504 15258 50516
rect 15289 50507 15347 50513
rect 15289 50504 15301 50507
rect 15252 50476 15301 50504
rect 15252 50464 15258 50476
rect 15289 50473 15301 50476
rect 15335 50504 15347 50507
rect 16114 50504 16120 50516
rect 15335 50476 16120 50504
rect 15335 50473 15347 50476
rect 15289 50467 15347 50473
rect 16114 50464 16120 50476
rect 16172 50464 16178 50516
rect 17678 50464 17684 50516
rect 17736 50504 17742 50516
rect 19613 50507 19671 50513
rect 19613 50504 19625 50507
rect 17736 50476 19625 50504
rect 17736 50464 17742 50476
rect 19613 50473 19625 50476
rect 19659 50473 19671 50507
rect 19613 50467 19671 50473
rect 13722 50396 13728 50448
rect 13780 50436 13786 50448
rect 15657 50439 15715 50445
rect 15657 50436 15669 50439
rect 13780 50408 15669 50436
rect 13780 50396 13786 50408
rect 15657 50405 15669 50408
rect 15703 50436 15715 50439
rect 17310 50436 17316 50448
rect 15703 50408 17316 50436
rect 15703 50405 15715 50408
rect 15657 50399 15715 50405
rect 17310 50396 17316 50408
rect 17368 50396 17374 50448
rect 15197 50303 15255 50309
rect 15197 50269 15209 50303
rect 15243 50300 15255 50303
rect 20530 50300 20536 50312
rect 15243 50272 20536 50300
rect 15243 50269 15255 50272
rect 15197 50263 15255 50269
rect 20530 50260 20536 50272
rect 20588 50260 20594 50312
rect 19521 50235 19579 50241
rect 19521 50201 19533 50235
rect 19567 50232 19579 50235
rect 20622 50232 20628 50244
rect 19567 50204 20628 50232
rect 19567 50201 19579 50204
rect 19521 50195 19579 50201
rect 20622 50192 20628 50204
rect 20680 50192 20686 50244
rect 1104 50074 49864 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 27950 50074
rect 28002 50022 28014 50074
rect 28066 50022 28078 50074
rect 28130 50022 28142 50074
rect 28194 50022 28206 50074
rect 28258 50022 37950 50074
rect 38002 50022 38014 50074
rect 38066 50022 38078 50074
rect 38130 50022 38142 50074
rect 38194 50022 38206 50074
rect 38258 50022 47950 50074
rect 48002 50022 48014 50074
rect 48066 50022 48078 50074
rect 48130 50022 48142 50074
rect 48194 50022 48206 50074
rect 48258 50022 49864 50074
rect 1104 50000 49864 50022
rect 49142 49784 49148 49836
rect 49200 49784 49206 49836
rect 49329 49759 49387 49765
rect 49329 49725 49341 49759
rect 49375 49756 49387 49759
rect 49510 49756 49516 49768
rect 49375 49728 49516 49756
rect 49375 49725 49387 49728
rect 49329 49719 49387 49725
rect 49510 49716 49516 49728
rect 49568 49716 49574 49768
rect 1104 49530 49864 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 32950 49530
rect 33002 49478 33014 49530
rect 33066 49478 33078 49530
rect 33130 49478 33142 49530
rect 33194 49478 33206 49530
rect 33258 49478 42950 49530
rect 43002 49478 43014 49530
rect 43066 49478 43078 49530
rect 43130 49478 43142 49530
rect 43194 49478 43206 49530
rect 43258 49478 49864 49530
rect 1104 49456 49864 49478
rect 20254 49376 20260 49428
rect 20312 49416 20318 49428
rect 20993 49419 21051 49425
rect 20993 49416 21005 49419
rect 20312 49388 21005 49416
rect 20312 49376 20318 49388
rect 20993 49385 21005 49388
rect 21039 49385 21051 49419
rect 20993 49379 21051 49385
rect 22830 49376 22836 49428
rect 22888 49416 22894 49428
rect 23017 49419 23075 49425
rect 23017 49416 23029 49419
rect 22888 49388 23029 49416
rect 22888 49376 22894 49388
rect 23017 49385 23029 49388
rect 23063 49385 23075 49419
rect 23017 49379 23075 49385
rect 20901 49147 20959 49153
rect 20901 49113 20913 49147
rect 20947 49144 20959 49147
rect 21450 49144 21456 49156
rect 20947 49116 21456 49144
rect 20947 49113 20959 49116
rect 20901 49107 20959 49113
rect 21450 49104 21456 49116
rect 21508 49104 21514 49156
rect 22925 49147 22983 49153
rect 22925 49113 22937 49147
rect 22971 49144 22983 49147
rect 23290 49144 23296 49156
rect 22971 49116 23296 49144
rect 22971 49113 22983 49116
rect 22925 49107 22983 49113
rect 23290 49104 23296 49116
rect 23348 49104 23354 49156
rect 49142 49104 49148 49156
rect 49200 49104 49206 49156
rect 49329 49147 49387 49153
rect 49329 49113 49341 49147
rect 49375 49144 49387 49147
rect 50430 49144 50436 49156
rect 49375 49116 50436 49144
rect 49375 49113 49387 49116
rect 49329 49107 49387 49113
rect 50430 49104 50436 49116
rect 50488 49104 50494 49156
rect 1104 48986 49864 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 27950 48986
rect 28002 48934 28014 48986
rect 28066 48934 28078 48986
rect 28130 48934 28142 48986
rect 28194 48934 28206 48986
rect 28258 48934 37950 48986
rect 38002 48934 38014 48986
rect 38066 48934 38078 48986
rect 38130 48934 38142 48986
rect 38194 48934 38206 48986
rect 38258 48934 47950 48986
rect 48002 48934 48014 48986
rect 48066 48934 48078 48986
rect 48130 48934 48142 48986
rect 48194 48934 48206 48986
rect 48258 48934 49864 48986
rect 1104 48912 49864 48934
rect 1104 48442 49864 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 32950 48442
rect 33002 48390 33014 48442
rect 33066 48390 33078 48442
rect 33130 48390 33142 48442
rect 33194 48390 33206 48442
rect 33258 48390 42950 48442
rect 43002 48390 43014 48442
rect 43066 48390 43078 48442
rect 43130 48390 43142 48442
rect 43194 48390 43206 48442
rect 43258 48390 49864 48442
rect 1104 48368 49864 48390
rect 16114 48220 16120 48272
rect 16172 48220 16178 48272
rect 14369 48195 14427 48201
rect 14369 48161 14381 48195
rect 14415 48192 14427 48195
rect 19426 48192 19432 48204
rect 14415 48164 19432 48192
rect 14415 48161 14427 48164
rect 14369 48155 14427 48161
rect 19426 48152 19432 48164
rect 19484 48152 19490 48204
rect 14645 48059 14703 48065
rect 14645 48025 14657 48059
rect 14691 48025 14703 48059
rect 18322 48056 18328 48068
rect 15870 48028 18328 48056
rect 14645 48019 14703 48025
rect 14660 47988 14688 48019
rect 18322 48016 18328 48028
rect 18380 48016 18386 48068
rect 49142 48016 49148 48068
rect 49200 48016 49206 48068
rect 19518 47988 19524 48000
rect 14660 47960 19524 47988
rect 19518 47948 19524 47960
rect 19576 47948 19582 48000
rect 33686 47948 33692 48000
rect 33744 47988 33750 48000
rect 49237 47991 49295 47997
rect 49237 47988 49249 47991
rect 33744 47960 49249 47988
rect 33744 47948 33750 47960
rect 49237 47957 49249 47960
rect 49283 47957 49295 47991
rect 49237 47951 49295 47957
rect 1104 47898 49864 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 27950 47898
rect 28002 47846 28014 47898
rect 28066 47846 28078 47898
rect 28130 47846 28142 47898
rect 28194 47846 28206 47898
rect 28258 47846 37950 47898
rect 38002 47846 38014 47898
rect 38066 47846 38078 47898
rect 38130 47846 38142 47898
rect 38194 47846 38206 47898
rect 38258 47846 47950 47898
rect 48002 47846 48014 47898
rect 48066 47846 48078 47898
rect 48130 47846 48142 47898
rect 48194 47846 48206 47898
rect 48258 47846 49864 47898
rect 1104 47824 49864 47846
rect 19794 47744 19800 47796
rect 19852 47744 19858 47796
rect 20530 47716 20536 47728
rect 19352 47688 20536 47716
rect 19352 47657 19380 47688
rect 20530 47676 20536 47688
rect 20588 47676 20594 47728
rect 19337 47651 19395 47657
rect 19337 47617 19349 47651
rect 19383 47617 19395 47651
rect 20292 47651 20350 47657
rect 20292 47648 20304 47651
rect 19337 47611 19395 47617
rect 19444 47620 20304 47648
rect 17310 47540 17316 47592
rect 17368 47580 17374 47592
rect 19444 47580 19472 47620
rect 20292 47617 20304 47620
rect 20338 47617 20350 47651
rect 20292 47611 20350 47617
rect 49326 47608 49332 47660
rect 49384 47608 49390 47660
rect 17368 47552 19472 47580
rect 17368 47540 17374 47552
rect 19518 47540 19524 47592
rect 19576 47580 19582 47592
rect 21174 47580 21180 47592
rect 19576 47552 21180 47580
rect 19576 47540 19582 47552
rect 21174 47540 21180 47552
rect 21232 47540 21238 47592
rect 19536 47453 19564 47540
rect 19521 47447 19579 47453
rect 19521 47413 19533 47447
rect 19567 47413 19579 47447
rect 19521 47407 19579 47413
rect 20395 47447 20453 47453
rect 20395 47413 20407 47447
rect 20441 47444 20453 47447
rect 22002 47444 22008 47456
rect 20441 47416 22008 47444
rect 20441 47413 20453 47416
rect 20395 47407 20453 47413
rect 22002 47404 22008 47416
rect 22060 47404 22066 47456
rect 46198 47404 46204 47456
rect 46256 47444 46262 47456
rect 49145 47447 49203 47453
rect 49145 47444 49157 47447
rect 46256 47416 49157 47444
rect 46256 47404 46262 47416
rect 49145 47413 49157 47416
rect 49191 47413 49203 47447
rect 49145 47407 49203 47413
rect 1104 47354 49864 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 32950 47354
rect 33002 47302 33014 47354
rect 33066 47302 33078 47354
rect 33130 47302 33142 47354
rect 33194 47302 33206 47354
rect 33258 47302 42950 47354
rect 43002 47302 43014 47354
rect 43066 47302 43078 47354
rect 43130 47302 43142 47354
rect 43194 47302 43206 47354
rect 43258 47302 49864 47354
rect 1104 47280 49864 47302
rect 25682 47064 25688 47116
rect 25740 47064 25746 47116
rect 19794 46996 19800 47048
rect 19852 47036 19858 47048
rect 22316 47039 22374 47045
rect 22316 47036 22328 47039
rect 19852 47008 22328 47036
rect 19852 46996 19858 47008
rect 22316 47005 22328 47008
rect 22362 47005 22374 47039
rect 22316 46999 22374 47005
rect 22419 46971 22477 46977
rect 22419 46937 22431 46971
rect 22465 46968 22477 46971
rect 25869 46971 25927 46977
rect 25869 46968 25881 46971
rect 22465 46940 25881 46968
rect 22465 46937 22477 46940
rect 22419 46931 22477 46937
rect 25869 46937 25881 46940
rect 25915 46937 25927 46971
rect 25869 46931 25927 46937
rect 27522 46928 27528 46980
rect 27580 46928 27586 46980
rect 1104 46810 49864 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 27950 46810
rect 28002 46758 28014 46810
rect 28066 46758 28078 46810
rect 28130 46758 28142 46810
rect 28194 46758 28206 46810
rect 28258 46758 37950 46810
rect 38002 46758 38014 46810
rect 38066 46758 38078 46810
rect 38130 46758 38142 46810
rect 38194 46758 38206 46810
rect 38258 46758 47950 46810
rect 48002 46758 48014 46810
rect 48066 46758 48078 46810
rect 48130 46758 48142 46810
rect 48194 46758 48206 46810
rect 48258 46758 49864 46810
rect 1104 46736 49864 46758
rect 20530 46656 20536 46708
rect 20588 46696 20594 46708
rect 22462 46696 22468 46708
rect 20588 46668 22468 46696
rect 20588 46656 20594 46668
rect 22462 46656 22468 46668
rect 22520 46656 22526 46708
rect 24394 46628 24400 46640
rect 23216 46600 24400 46628
rect 23216 46569 23244 46600
rect 24394 46588 24400 46600
rect 24452 46588 24458 46640
rect 23201 46563 23259 46569
rect 23201 46529 23213 46563
rect 23247 46529 23259 46563
rect 23201 46523 23259 46529
rect 49326 46520 49332 46572
rect 49384 46520 49390 46572
rect 22002 46452 22008 46504
rect 22060 46492 22066 46504
rect 23385 46495 23443 46501
rect 23385 46492 23397 46495
rect 22060 46464 23397 46492
rect 22060 46452 22066 46464
rect 23385 46461 23397 46464
rect 23431 46461 23443 46495
rect 23385 46455 23443 46461
rect 24762 46452 24768 46504
rect 24820 46452 24826 46504
rect 41230 46316 41236 46368
rect 41288 46356 41294 46368
rect 49145 46359 49203 46365
rect 49145 46356 49157 46359
rect 41288 46328 49157 46356
rect 41288 46316 41294 46328
rect 49145 46325 49157 46328
rect 49191 46325 49203 46359
rect 49145 46319 49203 46325
rect 1104 46266 49864 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 32950 46266
rect 33002 46214 33014 46266
rect 33066 46214 33078 46266
rect 33130 46214 33142 46266
rect 33194 46214 33206 46266
rect 33258 46214 42950 46266
rect 43002 46214 43014 46266
rect 43066 46214 43078 46266
rect 43130 46214 43142 46266
rect 43194 46214 43206 46266
rect 43258 46214 49864 46266
rect 1104 46192 49864 46214
rect 17494 46112 17500 46164
rect 17552 46112 17558 46164
rect 21453 46155 21511 46161
rect 21453 46121 21465 46155
rect 21499 46152 21511 46155
rect 21542 46152 21548 46164
rect 21499 46124 21548 46152
rect 21499 46121 21511 46124
rect 21453 46115 21511 46121
rect 21542 46112 21548 46124
rect 21600 46112 21606 46164
rect 21634 46112 21640 46164
rect 21692 46112 21698 46164
rect 20990 46044 20996 46096
rect 21048 46084 21054 46096
rect 21652 46084 21680 46112
rect 30834 46084 30840 46096
rect 21048 46056 21680 46084
rect 21048 46044 21054 46056
rect 17310 45976 17316 46028
rect 17368 45976 17374 46028
rect 17126 45908 17132 45960
rect 17184 45908 17190 45960
rect 20530 45908 20536 45960
rect 20588 45948 20594 45960
rect 21177 45951 21235 45957
rect 21177 45948 21189 45951
rect 20588 45920 21189 45948
rect 20588 45908 20594 45920
rect 21177 45917 21189 45920
rect 21223 45917 21235 45951
rect 21652 45948 21680 46056
rect 27356 46056 30840 46084
rect 27356 46025 27384 46056
rect 30834 46044 30840 46056
rect 30892 46044 30898 46096
rect 27341 46019 27399 46025
rect 27341 45985 27353 46019
rect 27387 45985 27399 46019
rect 27341 45979 27399 45985
rect 28902 45976 28908 46028
rect 28960 45976 28966 46028
rect 24616 45951 24674 45957
rect 24616 45948 24628 45951
rect 21652 45920 24628 45948
rect 21177 45911 21235 45917
rect 24616 45917 24628 45920
rect 24662 45917 24674 45951
rect 24616 45911 24674 45917
rect 49326 45908 49332 45960
rect 49384 45908 49390 45960
rect 24719 45883 24777 45889
rect 24719 45849 24731 45883
rect 24765 45880 24777 45883
rect 27525 45883 27583 45889
rect 27525 45880 27537 45883
rect 24765 45852 27537 45880
rect 24765 45849 24777 45852
rect 24719 45843 24777 45849
rect 27525 45849 27537 45852
rect 27571 45849 27583 45883
rect 27525 45843 27583 45849
rect 49145 45815 49203 45821
rect 49145 45781 49157 45815
rect 49191 45812 49203 45815
rect 49878 45812 49884 45824
rect 49191 45784 49884 45812
rect 49191 45781 49203 45784
rect 49145 45775 49203 45781
rect 49878 45772 49884 45784
rect 49936 45772 49942 45824
rect 1104 45722 49864 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 27950 45722
rect 28002 45670 28014 45722
rect 28066 45670 28078 45722
rect 28130 45670 28142 45722
rect 28194 45670 28206 45722
rect 28258 45670 37950 45722
rect 38002 45670 38014 45722
rect 38066 45670 38078 45722
rect 38130 45670 38142 45722
rect 38194 45670 38206 45722
rect 38258 45670 47950 45722
rect 48002 45670 48014 45722
rect 48066 45670 48078 45722
rect 48130 45670 48142 45722
rect 48194 45670 48206 45722
rect 48258 45670 49864 45722
rect 1104 45648 49864 45670
rect 22830 45432 22836 45484
rect 22888 45472 22894 45484
rect 25904 45475 25962 45481
rect 25904 45472 25916 45475
rect 22888 45444 25916 45472
rect 22888 45432 22894 45444
rect 25904 45441 25916 45444
rect 25950 45441 25962 45475
rect 25904 45435 25962 45441
rect 29546 45432 29552 45484
rect 29604 45432 29610 45484
rect 29733 45407 29791 45413
rect 29733 45404 29745 45407
rect 26206 45376 29745 45404
rect 26007 45271 26065 45277
rect 26007 45237 26019 45271
rect 26053 45268 26065 45271
rect 26206 45268 26234 45376
rect 29733 45373 29745 45376
rect 29779 45373 29791 45407
rect 29733 45367 29791 45373
rect 31386 45364 31392 45416
rect 31444 45364 31450 45416
rect 26053 45240 26234 45268
rect 26053 45237 26065 45240
rect 26007 45231 26065 45237
rect 1104 45178 49864 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 32950 45178
rect 33002 45126 33014 45178
rect 33066 45126 33078 45178
rect 33130 45126 33142 45178
rect 33194 45126 33206 45178
rect 33258 45126 42950 45178
rect 43002 45126 43014 45178
rect 43066 45126 43078 45178
rect 43130 45126 43142 45178
rect 43194 45126 43206 45178
rect 43258 45126 49864 45178
rect 1104 45104 49864 45126
rect 21174 45024 21180 45076
rect 21232 45024 21238 45076
rect 19705 44931 19763 44937
rect 19705 44897 19717 44931
rect 19751 44928 19763 44931
rect 21542 44928 21548 44940
rect 19751 44900 21548 44928
rect 19751 44897 19763 44900
rect 19705 44891 19763 44897
rect 21542 44888 21548 44900
rect 21600 44888 21606 44940
rect 19426 44820 19432 44872
rect 19484 44820 19490 44872
rect 49326 44820 49332 44872
rect 49384 44820 49390 44872
rect 23382 44792 23388 44804
rect 20930 44764 23388 44792
rect 18322 44684 18328 44736
rect 18380 44724 18386 44736
rect 21008 44724 21036 44764
rect 23382 44752 23388 44764
rect 23440 44752 23446 44804
rect 18380 44696 21036 44724
rect 18380 44684 18386 44696
rect 48682 44684 48688 44736
rect 48740 44724 48746 44736
rect 49145 44727 49203 44733
rect 49145 44724 49157 44727
rect 48740 44696 49157 44724
rect 48740 44684 48746 44696
rect 49145 44693 49157 44696
rect 49191 44693 49203 44727
rect 49145 44687 49203 44693
rect 1104 44634 49864 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 27950 44634
rect 28002 44582 28014 44634
rect 28066 44582 28078 44634
rect 28130 44582 28142 44634
rect 28194 44582 28206 44634
rect 28258 44582 37950 44634
rect 38002 44582 38014 44634
rect 38066 44582 38078 44634
rect 38130 44582 38142 44634
rect 38194 44582 38206 44634
rect 38258 44582 47950 44634
rect 48002 44582 48014 44634
rect 48066 44582 48078 44634
rect 48130 44582 48142 44634
rect 48194 44582 48206 44634
rect 48258 44582 49864 44634
rect 1104 44560 49864 44582
rect 20622 44480 20628 44532
rect 20680 44480 20686 44532
rect 22830 44480 22836 44532
rect 22888 44520 22894 44532
rect 22925 44523 22983 44529
rect 22925 44520 22937 44523
rect 22888 44492 22937 44520
rect 22888 44480 22894 44492
rect 22925 44489 22937 44492
rect 22971 44489 22983 44523
rect 22925 44483 22983 44489
rect 19794 44344 19800 44396
rect 19852 44384 19858 44396
rect 20165 44387 20223 44393
rect 20165 44384 20177 44387
rect 19852 44356 20177 44384
rect 19852 44344 19858 44356
rect 20165 44353 20177 44356
rect 20211 44353 20223 44387
rect 20165 44347 20223 44353
rect 22462 44344 22468 44396
rect 22520 44344 22526 44396
rect 49142 44344 49148 44396
rect 49200 44344 49206 44396
rect 19978 44276 19984 44328
rect 20036 44276 20042 44328
rect 49329 44251 49387 44257
rect 49329 44217 49341 44251
rect 49375 44248 49387 44251
rect 49694 44248 49700 44260
rect 49375 44220 49700 44248
rect 49375 44217 49387 44220
rect 49329 44211 49387 44217
rect 49694 44208 49700 44220
rect 49752 44208 49758 44260
rect 22554 44140 22560 44192
rect 22612 44140 22618 44192
rect 1104 44090 49864 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 32950 44090
rect 33002 44038 33014 44090
rect 33066 44038 33078 44090
rect 33130 44038 33142 44090
rect 33194 44038 33206 44090
rect 33258 44038 42950 44090
rect 43002 44038 43014 44090
rect 43066 44038 43078 44090
rect 43130 44038 43142 44090
rect 43194 44038 43206 44090
rect 43258 44038 49864 44090
rect 1104 44016 49864 44038
rect 41785 43843 41843 43849
rect 41785 43809 41797 43843
rect 41831 43840 41843 43843
rect 43438 43840 43444 43852
rect 41831 43812 43444 43840
rect 41831 43809 41843 43812
rect 41785 43803 41843 43809
rect 43438 43800 43444 43812
rect 43496 43800 43502 43852
rect 41414 43732 41420 43784
rect 41472 43772 41478 43784
rect 41509 43775 41567 43781
rect 41509 43772 41521 43775
rect 41472 43744 41521 43772
rect 41472 43732 41478 43744
rect 41509 43741 41521 43744
rect 41555 43741 41567 43775
rect 41509 43735 41567 43741
rect 42794 43664 42800 43716
rect 42852 43664 42858 43716
rect 34974 43596 34980 43648
rect 35032 43636 35038 43648
rect 43257 43639 43315 43645
rect 43257 43636 43269 43639
rect 35032 43608 43269 43636
rect 35032 43596 35038 43608
rect 43257 43605 43269 43608
rect 43303 43605 43315 43639
rect 43257 43599 43315 43605
rect 1104 43546 49864 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 27950 43546
rect 28002 43494 28014 43546
rect 28066 43494 28078 43546
rect 28130 43494 28142 43546
rect 28194 43494 28206 43546
rect 28258 43494 37950 43546
rect 38002 43494 38014 43546
rect 38066 43494 38078 43546
rect 38130 43494 38142 43546
rect 38194 43494 38206 43546
rect 38258 43494 47950 43546
rect 48002 43494 48014 43546
rect 48066 43494 48078 43546
rect 48130 43494 48142 43546
rect 48194 43494 48206 43546
rect 48258 43494 49864 43546
rect 1104 43472 49864 43494
rect 49142 43256 49148 43308
rect 49200 43256 49206 43308
rect 49329 43163 49387 43169
rect 49329 43129 49341 43163
rect 49375 43160 49387 43163
rect 49786 43160 49792 43172
rect 49375 43132 49792 43160
rect 49375 43129 49387 43132
rect 49329 43123 49387 43129
rect 49786 43120 49792 43132
rect 49844 43120 49850 43172
rect 1104 43002 49864 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 32950 43002
rect 33002 42950 33014 43002
rect 33066 42950 33078 43002
rect 33130 42950 33142 43002
rect 33194 42950 33206 43002
rect 33258 42950 42950 43002
rect 43002 42950 43014 43002
rect 43066 42950 43078 43002
rect 43130 42950 43142 43002
rect 43194 42950 43206 43002
rect 43258 42950 49864 43002
rect 1104 42928 49864 42950
rect 49142 42576 49148 42628
rect 49200 42576 49206 42628
rect 49234 42508 49240 42560
rect 49292 42508 49298 42560
rect 1104 42458 49864 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 27950 42458
rect 28002 42406 28014 42458
rect 28066 42406 28078 42458
rect 28130 42406 28142 42458
rect 28194 42406 28206 42458
rect 28258 42406 37950 42458
rect 38002 42406 38014 42458
rect 38066 42406 38078 42458
rect 38130 42406 38142 42458
rect 38194 42406 38206 42458
rect 38258 42406 47950 42458
rect 48002 42406 48014 42458
rect 48066 42406 48078 42458
rect 48130 42406 48142 42458
rect 48194 42406 48206 42458
rect 48258 42406 49864 42458
rect 1104 42384 49864 42406
rect 21450 42304 21456 42356
rect 21508 42304 21514 42356
rect 23017 42347 23075 42353
rect 23017 42313 23029 42347
rect 23063 42344 23075 42347
rect 23290 42344 23296 42356
rect 23063 42316 23296 42344
rect 23063 42313 23075 42316
rect 23017 42307 23075 42313
rect 23290 42304 23296 42316
rect 23348 42304 23354 42356
rect 20990 42168 20996 42220
rect 21048 42168 21054 42220
rect 22373 42211 22431 42217
rect 22373 42177 22385 42211
rect 22419 42208 22431 42211
rect 22646 42208 22652 42220
rect 22419 42180 22652 42208
rect 22419 42177 22431 42180
rect 22373 42171 22431 42177
rect 22646 42168 22652 42180
rect 22704 42168 22710 42220
rect 20806 42100 20812 42152
rect 20864 42100 20870 42152
rect 22557 42143 22615 42149
rect 22557 42109 22569 42143
rect 22603 42140 22615 42143
rect 22830 42140 22836 42152
rect 22603 42112 22836 42140
rect 22603 42109 22615 42112
rect 22557 42103 22615 42109
rect 22830 42100 22836 42112
rect 22888 42100 22894 42152
rect 1104 41914 49864 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 32950 41914
rect 33002 41862 33014 41914
rect 33066 41862 33078 41914
rect 33130 41862 33142 41914
rect 33194 41862 33206 41914
rect 33258 41862 42950 41914
rect 43002 41862 43014 41914
rect 43066 41862 43078 41914
rect 43130 41862 43142 41914
rect 43194 41862 43206 41914
rect 43258 41862 49864 41914
rect 1104 41840 49864 41862
rect 21542 41760 21548 41812
rect 21600 41800 21606 41812
rect 23293 41803 23351 41809
rect 23293 41800 23305 41803
rect 21600 41772 23305 41800
rect 21600 41760 21606 41772
rect 23293 41769 23305 41772
rect 23339 41769 23351 41803
rect 23293 41763 23351 41769
rect 19426 41624 19432 41676
rect 19484 41664 19490 41676
rect 21545 41667 21603 41673
rect 21545 41664 21557 41667
rect 19484 41636 21557 41664
rect 19484 41624 19490 41636
rect 21545 41633 21557 41636
rect 21591 41664 21603 41667
rect 22830 41664 22836 41676
rect 21591 41636 22836 41664
rect 21591 41633 21603 41636
rect 21545 41627 21603 41633
rect 22830 41624 22836 41636
rect 22888 41624 22894 41676
rect 23382 41624 23388 41676
rect 23440 41624 23446 41676
rect 23400 41596 23428 41624
rect 24302 41596 24308 41608
rect 22954 41568 24308 41596
rect 24302 41556 24308 41568
rect 24360 41556 24366 41608
rect 21821 41531 21879 41537
rect 21821 41497 21833 41531
rect 21867 41497 21879 41531
rect 23382 41528 23388 41540
rect 21821 41491 21879 41497
rect 23124 41500 23388 41528
rect 21836 41460 21864 41491
rect 22554 41460 22560 41472
rect 21836 41432 22560 41460
rect 22554 41420 22560 41432
rect 22612 41460 22618 41472
rect 23124 41460 23152 41500
rect 23382 41488 23388 41500
rect 23440 41488 23446 41540
rect 49142 41488 49148 41540
rect 49200 41488 49206 41540
rect 22612 41432 23152 41460
rect 22612 41420 22618 41432
rect 36814 41420 36820 41472
rect 36872 41460 36878 41472
rect 49237 41463 49295 41469
rect 49237 41460 49249 41463
rect 36872 41432 49249 41460
rect 36872 41420 36878 41432
rect 49237 41429 49249 41432
rect 49283 41429 49295 41463
rect 49237 41423 49295 41429
rect 1104 41370 49864 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 27950 41370
rect 28002 41318 28014 41370
rect 28066 41318 28078 41370
rect 28130 41318 28142 41370
rect 28194 41318 28206 41370
rect 28258 41318 37950 41370
rect 38002 41318 38014 41370
rect 38066 41318 38078 41370
rect 38130 41318 38142 41370
rect 38194 41318 38206 41370
rect 38258 41318 47950 41370
rect 48002 41318 48014 41370
rect 48066 41318 48078 41370
rect 48130 41318 48142 41370
rect 48194 41318 48206 41370
rect 48258 41318 49864 41370
rect 1104 41296 49864 41318
rect 49326 41080 49332 41132
rect 49384 41080 49390 41132
rect 48314 40876 48320 40928
rect 48372 40916 48378 40928
rect 49145 40919 49203 40925
rect 49145 40916 49157 40919
rect 48372 40888 49157 40916
rect 48372 40876 48378 40888
rect 49145 40885 49157 40888
rect 49191 40885 49203 40919
rect 49145 40879 49203 40885
rect 1104 40826 49864 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 32950 40826
rect 33002 40774 33014 40826
rect 33066 40774 33078 40826
rect 33130 40774 33142 40826
rect 33194 40774 33206 40826
rect 33258 40774 42950 40826
rect 43002 40774 43014 40826
rect 43066 40774 43078 40826
rect 43130 40774 43142 40826
rect 43194 40774 43206 40826
rect 43258 40774 49864 40826
rect 1104 40752 49864 40774
rect 1104 40282 49864 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 27950 40282
rect 28002 40230 28014 40282
rect 28066 40230 28078 40282
rect 28130 40230 28142 40282
rect 28194 40230 28206 40282
rect 28258 40230 37950 40282
rect 38002 40230 38014 40282
rect 38066 40230 38078 40282
rect 38130 40230 38142 40282
rect 38194 40230 38206 40282
rect 38258 40230 47950 40282
rect 48002 40230 48014 40282
rect 48066 40230 48078 40282
rect 48130 40230 48142 40282
rect 48194 40230 48206 40282
rect 48258 40230 49864 40282
rect 1104 40208 49864 40230
rect 49050 40128 49056 40180
rect 49108 40168 49114 40180
rect 49145 40171 49203 40177
rect 49145 40168 49157 40171
rect 49108 40140 49157 40168
rect 49108 40128 49114 40140
rect 49145 40137 49157 40140
rect 49191 40137 49203 40171
rect 49145 40131 49203 40137
rect 49326 39992 49332 40044
rect 49384 39992 49390 40044
rect 1104 39738 49864 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 32950 39738
rect 33002 39686 33014 39738
rect 33066 39686 33078 39738
rect 33130 39686 33142 39738
rect 33194 39686 33206 39738
rect 33258 39686 42950 39738
rect 43002 39686 43014 39738
rect 43066 39686 43078 39738
rect 43130 39686 43142 39738
rect 43194 39686 43206 39738
rect 43258 39686 49864 39738
rect 1104 39664 49864 39686
rect 49326 39380 49332 39432
rect 49384 39380 49390 39432
rect 48590 39244 48596 39296
rect 48648 39284 48654 39296
rect 49145 39287 49203 39293
rect 49145 39284 49157 39287
rect 48648 39256 49157 39284
rect 48648 39244 48654 39256
rect 49145 39253 49157 39256
rect 49191 39253 49203 39287
rect 49145 39247 49203 39253
rect 1104 39194 49864 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 27950 39194
rect 28002 39142 28014 39194
rect 28066 39142 28078 39194
rect 28130 39142 28142 39194
rect 28194 39142 28206 39194
rect 28258 39142 37950 39194
rect 38002 39142 38014 39194
rect 38066 39142 38078 39194
rect 38130 39142 38142 39194
rect 38194 39142 38206 39194
rect 38258 39142 47950 39194
rect 48002 39142 48014 39194
rect 48066 39142 48078 39194
rect 48130 39142 48142 39194
rect 48194 39142 48206 39194
rect 48258 39142 49864 39194
rect 1104 39120 49864 39142
rect 1104 38650 49864 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 32950 38650
rect 33002 38598 33014 38650
rect 33066 38598 33078 38650
rect 33130 38598 33142 38650
rect 33194 38598 33206 38650
rect 33258 38598 42950 38650
rect 43002 38598 43014 38650
rect 43066 38598 43078 38650
rect 43130 38598 43142 38650
rect 43194 38598 43206 38650
rect 43258 38598 49864 38650
rect 1104 38576 49864 38598
rect 49326 38292 49332 38344
rect 49384 38292 49390 38344
rect 48958 38156 48964 38208
rect 49016 38196 49022 38208
rect 49145 38199 49203 38205
rect 49145 38196 49157 38199
rect 49016 38168 49157 38196
rect 49016 38156 49022 38168
rect 49145 38165 49157 38168
rect 49191 38165 49203 38199
rect 49145 38159 49203 38165
rect 1104 38106 49864 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 27950 38106
rect 28002 38054 28014 38106
rect 28066 38054 28078 38106
rect 28130 38054 28142 38106
rect 28194 38054 28206 38106
rect 28258 38054 37950 38106
rect 38002 38054 38014 38106
rect 38066 38054 38078 38106
rect 38130 38054 38142 38106
rect 38194 38054 38206 38106
rect 38258 38054 47950 38106
rect 48002 38054 48014 38106
rect 48066 38054 48078 38106
rect 48130 38054 48142 38106
rect 48194 38054 48206 38106
rect 48258 38054 49864 38106
rect 1104 38032 49864 38054
rect 49142 37816 49148 37868
rect 49200 37816 49206 37868
rect 49329 37723 49387 37729
rect 49329 37689 49341 37723
rect 49375 37720 49387 37723
rect 50522 37720 50528 37732
rect 49375 37692 50528 37720
rect 49375 37689 49387 37692
rect 49329 37683 49387 37689
rect 50522 37680 50528 37692
rect 50580 37680 50586 37732
rect 1104 37562 49864 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 32950 37562
rect 33002 37510 33014 37562
rect 33066 37510 33078 37562
rect 33130 37510 33142 37562
rect 33194 37510 33206 37562
rect 33258 37510 42950 37562
rect 43002 37510 43014 37562
rect 43066 37510 43078 37562
rect 43130 37510 43142 37562
rect 43194 37510 43206 37562
rect 43258 37510 49864 37562
rect 1104 37488 49864 37510
rect 20441 37247 20499 37253
rect 20441 37213 20453 37247
rect 20487 37244 20499 37247
rect 22554 37244 22560 37256
rect 20487 37216 22560 37244
rect 20487 37213 20499 37216
rect 20441 37207 20499 37213
rect 22554 37204 22560 37216
rect 22612 37204 22618 37256
rect 17126 37068 17132 37120
rect 17184 37108 17190 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 17184 37080 20269 37108
rect 17184 37068 17190 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 1104 37018 49864 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 27950 37018
rect 28002 36966 28014 37018
rect 28066 36966 28078 37018
rect 28130 36966 28142 37018
rect 28194 36966 28206 37018
rect 28258 36966 37950 37018
rect 38002 36966 38014 37018
rect 38066 36966 38078 37018
rect 38130 36966 38142 37018
rect 38194 36966 38206 37018
rect 38258 36966 47950 37018
rect 48002 36966 48014 37018
rect 48066 36966 48078 37018
rect 48130 36966 48142 37018
rect 48194 36966 48206 37018
rect 48258 36966 49864 37018
rect 1104 36944 49864 36966
rect 49142 36728 49148 36780
rect 49200 36728 49206 36780
rect 48774 36524 48780 36576
rect 48832 36564 48838 36576
rect 49237 36567 49295 36573
rect 49237 36564 49249 36567
rect 48832 36536 49249 36564
rect 48832 36524 48838 36536
rect 49237 36533 49249 36536
rect 49283 36533 49295 36567
rect 49237 36527 49295 36533
rect 49418 36524 49424 36576
rect 49476 36564 49482 36576
rect 49694 36564 49700 36576
rect 49476 36536 49700 36564
rect 49476 36524 49482 36536
rect 49694 36524 49700 36536
rect 49752 36524 49758 36576
rect 1104 36474 49864 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 32950 36474
rect 33002 36422 33014 36474
rect 33066 36422 33078 36474
rect 33130 36422 33142 36474
rect 33194 36422 33206 36474
rect 33258 36422 42950 36474
rect 43002 36422 43014 36474
rect 43066 36422 43078 36474
rect 43130 36422 43142 36474
rect 43194 36422 43206 36474
rect 43258 36422 49864 36474
rect 1104 36400 49864 36422
rect 49326 36116 49332 36168
rect 49384 36116 49390 36168
rect 49145 36023 49203 36029
rect 49145 35989 49157 36023
rect 49191 36020 49203 36023
rect 49694 36020 49700 36032
rect 49191 35992 49700 36020
rect 49191 35989 49203 35992
rect 49145 35983 49203 35989
rect 49694 35980 49700 35992
rect 49752 35980 49758 36032
rect 1104 35930 49864 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 27950 35930
rect 28002 35878 28014 35930
rect 28066 35878 28078 35930
rect 28130 35878 28142 35930
rect 28194 35878 28206 35930
rect 28258 35878 37950 35930
rect 38002 35878 38014 35930
rect 38066 35878 38078 35930
rect 38130 35878 38142 35930
rect 38194 35878 38206 35930
rect 38258 35878 47950 35930
rect 48002 35878 48014 35930
rect 48066 35878 48078 35930
rect 48130 35878 48142 35930
rect 48194 35878 48206 35930
rect 48258 35878 49864 35930
rect 1104 35856 49864 35878
rect 1104 35386 49864 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 32950 35386
rect 33002 35334 33014 35386
rect 33066 35334 33078 35386
rect 33130 35334 33142 35386
rect 33194 35334 33206 35386
rect 33258 35334 42950 35386
rect 43002 35334 43014 35386
rect 43066 35334 43078 35386
rect 43130 35334 43142 35386
rect 43194 35334 43206 35386
rect 43258 35334 49864 35386
rect 1104 35312 49864 35334
rect 49326 35028 49332 35080
rect 49384 35028 49390 35080
rect 49145 34935 49203 34941
rect 49145 34901 49157 34935
rect 49191 34932 49203 34935
rect 50062 34932 50068 34944
rect 49191 34904 50068 34932
rect 49191 34901 49203 34904
rect 49145 34895 49203 34901
rect 50062 34892 50068 34904
rect 50120 34892 50126 34944
rect 1104 34842 49864 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 27950 34842
rect 28002 34790 28014 34842
rect 28066 34790 28078 34842
rect 28130 34790 28142 34842
rect 28194 34790 28206 34842
rect 28258 34790 37950 34842
rect 38002 34790 38014 34842
rect 38066 34790 38078 34842
rect 38130 34790 38142 34842
rect 38194 34790 38206 34842
rect 38258 34790 47950 34842
rect 48002 34790 48014 34842
rect 48066 34790 48078 34842
rect 48130 34790 48142 34842
rect 48194 34790 48206 34842
rect 48258 34790 49864 34842
rect 1104 34768 49864 34790
rect 23382 34688 23388 34740
rect 23440 34728 23446 34740
rect 24673 34731 24731 34737
rect 24673 34728 24685 34731
rect 23440 34700 24685 34728
rect 23440 34688 23446 34700
rect 24673 34697 24685 34700
rect 24719 34697 24731 34731
rect 24673 34691 24731 34697
rect 44174 34688 44180 34740
rect 44232 34728 44238 34740
rect 49145 34731 49203 34737
rect 49145 34728 49157 34731
rect 44232 34700 49157 34728
rect 44232 34688 44238 34700
rect 49145 34697 49157 34700
rect 49191 34697 49203 34731
rect 49145 34691 49203 34697
rect 24302 34552 24308 34604
rect 24360 34552 24366 34604
rect 49326 34552 49332 34604
rect 49384 34552 49390 34604
rect 22830 34484 22836 34536
rect 22888 34524 22894 34536
rect 22925 34527 22983 34533
rect 22925 34524 22937 34527
rect 22888 34496 22937 34524
rect 22888 34484 22894 34496
rect 22925 34493 22937 34496
rect 22971 34493 22983 34527
rect 22925 34487 22983 34493
rect 23188 34391 23246 34397
rect 23188 34357 23200 34391
rect 23234 34388 23246 34391
rect 24210 34388 24216 34400
rect 23234 34360 24216 34388
rect 23234 34357 23246 34360
rect 23188 34351 23246 34357
rect 24210 34348 24216 34360
rect 24268 34348 24274 34400
rect 1104 34298 49864 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 32950 34298
rect 33002 34246 33014 34298
rect 33066 34246 33078 34298
rect 33130 34246 33142 34298
rect 33194 34246 33206 34298
rect 33258 34246 42950 34298
rect 43002 34246 43014 34298
rect 43066 34246 43078 34298
rect 43130 34246 43142 34298
rect 43194 34246 43206 34298
rect 43258 34246 49864 34298
rect 1104 34224 49864 34246
rect 19978 34144 19984 34196
rect 20036 34184 20042 34196
rect 22833 34187 22891 34193
rect 22833 34184 22845 34187
rect 20036 34156 22845 34184
rect 20036 34144 20042 34156
rect 22833 34153 22845 34156
rect 22879 34153 22891 34187
rect 22833 34147 22891 34153
rect 38378 34076 38384 34128
rect 38436 34116 38442 34128
rect 42153 34119 42211 34125
rect 42153 34116 42165 34119
rect 38436 34088 42165 34116
rect 38436 34076 38442 34088
rect 42153 34085 42165 34088
rect 42199 34085 42211 34119
rect 43714 34116 43720 34128
rect 42153 34079 42211 34085
rect 42444 34088 43720 34116
rect 41230 34008 41236 34060
rect 41288 34048 41294 34060
rect 41417 34051 41475 34057
rect 41417 34048 41429 34051
rect 41288 34020 41429 34048
rect 41288 34008 41294 34020
rect 41417 34017 41429 34020
rect 41463 34017 41475 34051
rect 41417 34011 41475 34017
rect 41509 34051 41567 34057
rect 41509 34017 41521 34051
rect 41555 34017 41567 34051
rect 41509 34011 41567 34017
rect 22738 33940 22744 33992
rect 22796 33980 22802 33992
rect 23017 33983 23075 33989
rect 23017 33980 23029 33983
rect 22796 33952 23029 33980
rect 22796 33940 22802 33952
rect 23017 33949 23029 33952
rect 23063 33949 23075 33983
rect 23017 33943 23075 33949
rect 39666 33940 39672 33992
rect 39724 33980 39730 33992
rect 41524 33980 41552 34011
rect 39724 33952 41552 33980
rect 39724 33940 39730 33952
rect 41325 33915 41383 33921
rect 41325 33912 41337 33915
rect 40420 33884 41337 33912
rect 27522 33804 27528 33856
rect 27580 33844 27586 33856
rect 40420 33853 40448 33884
rect 41325 33881 41337 33884
rect 41371 33912 41383 33915
rect 42444 33912 42472 34088
rect 43714 34076 43720 34088
rect 43772 34076 43778 34128
rect 42702 34008 42708 34060
rect 42760 34008 42766 34060
rect 42886 34008 42892 34060
rect 42944 34048 42950 34060
rect 49878 34048 49884 34060
rect 42944 34020 49884 34048
rect 42944 34008 42950 34020
rect 49878 34008 49884 34020
rect 49936 34008 49942 34060
rect 42521 33983 42579 33989
rect 42521 33949 42533 33983
rect 42567 33980 42579 33983
rect 42567 33952 43852 33980
rect 42567 33949 42579 33952
rect 42521 33943 42579 33949
rect 41371 33884 42472 33912
rect 41371 33881 41383 33884
rect 41325 33875 41383 33881
rect 40405 33847 40463 33853
rect 40405 33844 40417 33847
rect 27580 33816 40417 33844
rect 27580 33804 27586 33816
rect 40405 33813 40417 33816
rect 40451 33813 40463 33847
rect 40405 33807 40463 33813
rect 40954 33804 40960 33856
rect 41012 33804 41018 33856
rect 41230 33804 41236 33856
rect 41288 33844 41294 33856
rect 42536 33844 42564 33943
rect 43824 33856 43852 33952
rect 41288 33816 42564 33844
rect 42613 33847 42671 33853
rect 41288 33804 41294 33816
rect 42613 33813 42625 33847
rect 42659 33844 42671 33847
rect 42886 33844 42892 33856
rect 42659 33816 42892 33844
rect 42659 33813 42671 33816
rect 42613 33807 42671 33813
rect 42886 33804 42892 33816
rect 42944 33804 42950 33856
rect 43441 33847 43499 33853
rect 43441 33813 43453 33847
rect 43487 33844 43499 33847
rect 43806 33844 43812 33856
rect 43487 33816 43812 33844
rect 43487 33813 43499 33816
rect 43441 33807 43499 33813
rect 43806 33804 43812 33816
rect 43864 33804 43870 33856
rect 1104 33754 49864 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 27950 33754
rect 28002 33702 28014 33754
rect 28066 33702 28078 33754
rect 28130 33702 28142 33754
rect 28194 33702 28206 33754
rect 28258 33702 37950 33754
rect 38002 33702 38014 33754
rect 38066 33702 38078 33754
rect 38130 33702 38142 33754
rect 38194 33702 38206 33754
rect 38258 33702 47950 33754
rect 48002 33702 48014 33754
rect 48066 33702 48078 33754
rect 48130 33702 48142 33754
rect 48194 33702 48206 33754
rect 48258 33702 49864 33754
rect 1104 33680 49864 33702
rect 43073 33643 43131 33649
rect 43073 33609 43085 33643
rect 43119 33640 43131 33643
rect 48682 33640 48688 33652
rect 43119 33612 48688 33640
rect 43119 33609 43131 33612
rect 43073 33603 43131 33609
rect 48682 33600 48688 33612
rect 48740 33600 48746 33652
rect 42981 33507 43039 33513
rect 42981 33504 42993 33507
rect 41386 33476 42993 33504
rect 31386 33328 31392 33380
rect 31444 33368 31450 33380
rect 41386 33368 41414 33476
rect 42981 33473 42993 33476
rect 43027 33504 43039 33507
rect 43622 33504 43628 33516
rect 43027 33476 43628 33504
rect 43027 33473 43039 33476
rect 42981 33467 43039 33473
rect 43622 33464 43628 33476
rect 43680 33464 43686 33516
rect 49326 33464 49332 33516
rect 49384 33464 49390 33516
rect 43257 33439 43315 33445
rect 43257 33405 43269 33439
rect 43303 33436 43315 33439
rect 43530 33436 43536 33448
rect 43303 33408 43536 33436
rect 43303 33405 43315 33408
rect 43257 33399 43315 33405
rect 43530 33396 43536 33408
rect 43588 33396 43594 33448
rect 31444 33340 41414 33368
rect 31444 33328 31450 33340
rect 40218 33260 40224 33312
rect 40276 33300 40282 33312
rect 42613 33303 42671 33309
rect 42613 33300 42625 33303
rect 40276 33272 42625 33300
rect 40276 33260 40282 33272
rect 42613 33269 42625 33272
rect 42659 33269 42671 33303
rect 42613 33263 42671 33269
rect 43622 33260 43628 33312
rect 43680 33300 43686 33312
rect 43809 33303 43867 33309
rect 43809 33300 43821 33303
rect 43680 33272 43821 33300
rect 43680 33260 43686 33272
rect 43809 33269 43821 33272
rect 43855 33269 43867 33303
rect 43809 33263 43867 33269
rect 46842 33260 46848 33312
rect 46900 33300 46906 33312
rect 49145 33303 49203 33309
rect 49145 33300 49157 33303
rect 46900 33272 49157 33300
rect 46900 33260 46906 33272
rect 49145 33269 49157 33272
rect 49191 33269 49203 33303
rect 49145 33263 49203 33269
rect 1104 33210 49864 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 32950 33210
rect 33002 33158 33014 33210
rect 33066 33158 33078 33210
rect 33130 33158 33142 33210
rect 33194 33158 33206 33210
rect 33258 33158 42950 33210
rect 43002 33158 43014 33210
rect 43066 33158 43078 33210
rect 43130 33158 43142 33210
rect 43194 33158 43206 33210
rect 43258 33158 49864 33210
rect 1104 33136 49864 33158
rect 49326 32852 49332 32904
rect 49384 32852 49390 32904
rect 47394 32716 47400 32768
rect 47452 32756 47458 32768
rect 49145 32759 49203 32765
rect 49145 32756 49157 32759
rect 47452 32728 49157 32756
rect 47452 32716 47458 32728
rect 49145 32725 49157 32728
rect 49191 32725 49203 32759
rect 49145 32719 49203 32725
rect 1104 32666 49864 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 27950 32666
rect 28002 32614 28014 32666
rect 28066 32614 28078 32666
rect 28130 32614 28142 32666
rect 28194 32614 28206 32666
rect 28258 32614 37950 32666
rect 38002 32614 38014 32666
rect 38066 32614 38078 32666
rect 38130 32614 38142 32666
rect 38194 32614 38206 32666
rect 38258 32614 47950 32666
rect 48002 32614 48014 32666
rect 48066 32614 48078 32666
rect 48130 32614 48142 32666
rect 48194 32614 48206 32666
rect 48258 32614 49864 32666
rect 1104 32592 49864 32614
rect 40126 32484 40132 32496
rect 39974 32456 40132 32484
rect 40126 32444 40132 32456
rect 40184 32484 40190 32496
rect 41506 32484 41512 32496
rect 40184 32456 41512 32484
rect 40184 32444 40190 32456
rect 41506 32444 41512 32456
rect 41564 32444 41570 32496
rect 38470 32308 38476 32360
rect 38528 32308 38534 32360
rect 38749 32351 38807 32357
rect 38749 32317 38761 32351
rect 38795 32348 38807 32351
rect 41782 32348 41788 32360
rect 38795 32320 41788 32348
rect 38795 32317 38807 32320
rect 38749 32311 38807 32317
rect 41782 32308 41788 32320
rect 41840 32308 41846 32360
rect 38286 32172 38292 32224
rect 38344 32212 38350 32224
rect 40221 32215 40279 32221
rect 40221 32212 40233 32215
rect 38344 32184 40233 32212
rect 38344 32172 38350 32184
rect 40221 32181 40233 32184
rect 40267 32181 40279 32215
rect 40221 32175 40279 32181
rect 1104 32122 49864 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 32950 32122
rect 33002 32070 33014 32122
rect 33066 32070 33078 32122
rect 33130 32070 33142 32122
rect 33194 32070 33206 32122
rect 33258 32070 42950 32122
rect 43002 32070 43014 32122
rect 43066 32070 43078 32122
rect 43130 32070 43142 32122
rect 43194 32070 43206 32122
rect 43258 32070 49864 32122
rect 1104 32048 49864 32070
rect 42797 32011 42855 32017
rect 42797 32008 42809 32011
rect 26206 31980 42809 32008
rect 24394 31832 24400 31884
rect 24452 31872 24458 31884
rect 24762 31872 24768 31884
rect 24452 31844 24768 31872
rect 24452 31832 24458 31844
rect 24762 31832 24768 31844
rect 24820 31872 24826 31884
rect 26206 31872 26234 31980
rect 42797 31977 42809 31980
rect 42843 32008 42855 32011
rect 42886 32008 42892 32020
rect 42843 31980 42892 32008
rect 42843 31977 42855 31980
rect 42797 31971 42855 31977
rect 42886 31968 42892 31980
rect 42944 31968 42950 32020
rect 41782 31900 41788 31952
rect 41840 31900 41846 31952
rect 41874 31900 41880 31952
rect 41932 31940 41938 31952
rect 43257 31943 43315 31949
rect 43257 31940 43269 31943
rect 41932 31912 43269 31940
rect 41932 31900 41938 31912
rect 43257 31909 43269 31912
rect 43303 31909 43315 31943
rect 43257 31903 43315 31909
rect 45646 31900 45652 31952
rect 45704 31940 45710 31952
rect 49145 31943 49203 31949
rect 49145 31940 49157 31943
rect 45704 31912 49157 31940
rect 45704 31900 45710 31912
rect 49145 31909 49157 31912
rect 49191 31909 49203 31943
rect 49145 31903 49203 31909
rect 24820 31844 26234 31872
rect 24820 31832 24826 31844
rect 40310 31832 40316 31884
rect 40368 31832 40374 31884
rect 41506 31872 41512 31884
rect 41432 31844 41512 31872
rect 40034 31764 40040 31816
rect 40092 31764 40098 31816
rect 41432 31790 41460 31844
rect 41506 31832 41512 31844
rect 41564 31832 41570 31884
rect 41800 31872 41828 31900
rect 42702 31872 42708 31884
rect 41800 31844 42708 31872
rect 42702 31832 42708 31844
rect 42760 31832 42766 31884
rect 43346 31832 43352 31884
rect 43404 31872 43410 31884
rect 43809 31875 43867 31881
rect 43809 31872 43821 31875
rect 43404 31844 43821 31872
rect 43404 31832 43410 31844
rect 43809 31841 43821 31844
rect 43855 31841 43867 31875
rect 43809 31835 43867 31841
rect 42886 31764 42892 31816
rect 42944 31804 42950 31816
rect 43625 31807 43683 31813
rect 43625 31804 43637 31807
rect 42944 31776 43637 31804
rect 42944 31764 42950 31776
rect 43625 31773 43637 31776
rect 43671 31773 43683 31807
rect 43625 31767 43683 31773
rect 43717 31807 43775 31813
rect 43717 31773 43729 31807
rect 43763 31804 43775 31807
rect 48314 31804 48320 31816
rect 43763 31776 48320 31804
rect 43763 31773 43775 31776
rect 43717 31767 43775 31773
rect 48314 31764 48320 31776
rect 48372 31764 48378 31816
rect 49326 31764 49332 31816
rect 49384 31764 49390 31816
rect 34330 31628 34336 31680
rect 34388 31668 34394 31680
rect 46934 31668 46940 31680
rect 34388 31640 46940 31668
rect 34388 31628 34394 31640
rect 46934 31628 46940 31640
rect 46992 31628 46998 31680
rect 1104 31578 49864 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 27950 31578
rect 28002 31526 28014 31578
rect 28066 31526 28078 31578
rect 28130 31526 28142 31578
rect 28194 31526 28206 31578
rect 28258 31526 37950 31578
rect 38002 31526 38014 31578
rect 38066 31526 38078 31578
rect 38130 31526 38142 31578
rect 38194 31526 38206 31578
rect 38258 31526 47950 31578
rect 48002 31526 48014 31578
rect 48066 31526 48078 31578
rect 48130 31526 48142 31578
rect 48194 31526 48206 31578
rect 48258 31526 49864 31578
rect 1104 31504 49864 31526
rect 41414 31464 41420 31476
rect 40328 31436 41420 31464
rect 38470 31396 38476 31408
rect 37936 31368 38476 31396
rect 33965 31331 34023 31337
rect 33965 31297 33977 31331
rect 34011 31328 34023 31331
rect 34330 31328 34336 31340
rect 34011 31300 34336 31328
rect 34011 31297 34023 31300
rect 33965 31291 34023 31297
rect 34330 31288 34336 31300
rect 34388 31328 34394 31340
rect 34793 31331 34851 31337
rect 34793 31328 34805 31331
rect 34388 31300 34805 31328
rect 34388 31288 34394 31300
rect 34793 31297 34805 31300
rect 34839 31297 34851 31331
rect 34793 31291 34851 31297
rect 34885 31331 34943 31337
rect 34885 31297 34897 31331
rect 34931 31328 34943 31331
rect 35158 31328 35164 31340
rect 34931 31300 35164 31328
rect 34931 31297 34943 31300
rect 34885 31291 34943 31297
rect 35158 31288 35164 31300
rect 35216 31288 35222 31340
rect 37936 31337 37964 31368
rect 38470 31356 38476 31368
rect 38528 31356 38534 31408
rect 40126 31396 40132 31408
rect 39422 31368 40132 31396
rect 40126 31356 40132 31368
rect 40184 31356 40190 31408
rect 37921 31331 37979 31337
rect 37921 31297 37933 31331
rect 37967 31297 37979 31331
rect 37921 31291 37979 31297
rect 40034 31288 40040 31340
rect 40092 31328 40098 31340
rect 40328 31337 40356 31436
rect 41414 31424 41420 31436
rect 41472 31424 41478 31476
rect 41506 31424 41512 31476
rect 41564 31464 41570 31476
rect 41564 31436 41920 31464
rect 41564 31424 41570 31436
rect 41892 31396 41920 31436
rect 43714 31424 43720 31476
rect 43772 31424 43778 31476
rect 43809 31467 43867 31473
rect 43809 31433 43821 31467
rect 43855 31464 43867 31467
rect 49050 31464 49056 31476
rect 43855 31436 49056 31464
rect 43855 31433 43867 31436
rect 43809 31427 43867 31433
rect 49050 31424 49056 31436
rect 49108 31424 49114 31476
rect 42794 31396 42800 31408
rect 41814 31368 42800 31396
rect 42794 31356 42800 31368
rect 42852 31356 42858 31408
rect 42886 31356 42892 31408
rect 42944 31396 42950 31408
rect 43898 31396 43904 31408
rect 42944 31368 43904 31396
rect 42944 31356 42950 31368
rect 43898 31356 43904 31368
rect 43956 31356 43962 31408
rect 40313 31331 40371 31337
rect 40313 31328 40325 31331
rect 40092 31300 40325 31328
rect 40092 31288 40098 31300
rect 40313 31297 40325 31300
rect 40359 31297 40371 31331
rect 40313 31291 40371 31297
rect 49326 31288 49332 31340
rect 49384 31288 49390 31340
rect 34974 31220 34980 31272
rect 35032 31260 35038 31272
rect 35069 31263 35127 31269
rect 35069 31260 35081 31263
rect 35032 31232 35081 31260
rect 35032 31220 35038 31232
rect 35069 31229 35081 31232
rect 35115 31260 35127 31263
rect 35618 31260 35624 31272
rect 35115 31232 35624 31260
rect 35115 31229 35127 31232
rect 35069 31223 35127 31229
rect 35618 31220 35624 31232
rect 35676 31220 35682 31272
rect 38197 31263 38255 31269
rect 38197 31229 38209 31263
rect 38243 31260 38255 31263
rect 38286 31260 38292 31272
rect 38243 31232 38292 31260
rect 38243 31229 38255 31232
rect 38197 31223 38255 31229
rect 38286 31220 38292 31232
rect 38344 31260 38350 31272
rect 38562 31260 38568 31272
rect 38344 31232 38568 31260
rect 38344 31220 38350 31232
rect 38562 31220 38568 31232
rect 38620 31220 38626 31272
rect 40589 31263 40647 31269
rect 40589 31229 40601 31263
rect 40635 31260 40647 31263
rect 43530 31260 43536 31272
rect 40635 31232 43536 31260
rect 40635 31229 40647 31232
rect 40589 31223 40647 31229
rect 43530 31220 43536 31232
rect 43588 31220 43594 31272
rect 43901 31263 43959 31269
rect 43901 31229 43913 31263
rect 43947 31229 43959 31263
rect 43901 31223 43959 31229
rect 31478 31152 31484 31204
rect 31536 31192 31542 31204
rect 34425 31195 34483 31201
rect 34425 31192 34437 31195
rect 31536 31164 34437 31192
rect 31536 31152 31542 31164
rect 34425 31161 34437 31164
rect 34471 31161 34483 31195
rect 34425 31155 34483 31161
rect 42518 31152 42524 31204
rect 42576 31192 42582 31204
rect 43916 31192 43944 31223
rect 42576 31164 43944 31192
rect 42576 31152 42582 31164
rect 39666 31084 39672 31136
rect 39724 31084 39730 31136
rect 40310 31084 40316 31136
rect 40368 31124 40374 31136
rect 42061 31127 42119 31133
rect 42061 31124 42073 31127
rect 40368 31096 42073 31124
rect 40368 31084 40374 31096
rect 42061 31093 42073 31096
rect 42107 31093 42119 31127
rect 42061 31087 42119 31093
rect 43349 31127 43407 31133
rect 43349 31093 43361 31127
rect 43395 31124 43407 31127
rect 43438 31124 43444 31136
rect 43395 31096 43444 31124
rect 43395 31093 43407 31096
rect 43349 31087 43407 31093
rect 43438 31084 43444 31096
rect 43496 31084 43502 31136
rect 48314 31084 48320 31136
rect 48372 31124 48378 31136
rect 49145 31127 49203 31133
rect 49145 31124 49157 31127
rect 48372 31096 49157 31124
rect 48372 31084 48378 31096
rect 49145 31093 49157 31096
rect 49191 31093 49203 31127
rect 49145 31087 49203 31093
rect 1104 31034 49864 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 32950 31034
rect 33002 30982 33014 31034
rect 33066 30982 33078 31034
rect 33130 30982 33142 31034
rect 33194 30982 33206 31034
rect 33258 30982 42950 31034
rect 43002 30982 43014 31034
rect 43066 30982 43078 31034
rect 43130 30982 43142 31034
rect 43194 30982 43206 31034
rect 43258 30982 49864 31034
rect 1104 30960 49864 30982
rect 20806 30880 20812 30932
rect 20864 30920 20870 30932
rect 22281 30923 22339 30929
rect 22281 30920 22293 30923
rect 20864 30892 22293 30920
rect 20864 30880 20870 30892
rect 22281 30889 22293 30892
rect 22327 30889 22339 30923
rect 22281 30883 22339 30889
rect 22646 30880 22652 30932
rect 22704 30920 22710 30932
rect 22925 30923 22983 30929
rect 22925 30920 22937 30923
rect 22704 30892 22937 30920
rect 22704 30880 22710 30892
rect 22925 30889 22937 30892
rect 22971 30889 22983 30923
rect 22925 30883 22983 30889
rect 43165 30923 43223 30929
rect 43165 30889 43177 30923
rect 43211 30920 43223 30923
rect 43530 30920 43536 30932
rect 43211 30892 43536 30920
rect 43211 30889 43223 30892
rect 43165 30883 43223 30889
rect 43530 30880 43536 30892
rect 43588 30880 43594 30932
rect 39942 30744 39948 30796
rect 40000 30784 40006 30796
rect 40773 30787 40831 30793
rect 40773 30784 40785 30787
rect 40000 30756 40785 30784
rect 40000 30744 40006 30756
rect 40773 30753 40785 30756
rect 40819 30753 40831 30787
rect 40773 30747 40831 30753
rect 41414 30744 41420 30796
rect 41472 30744 41478 30796
rect 22462 30676 22468 30728
rect 22520 30676 22526 30728
rect 23109 30719 23167 30725
rect 23109 30685 23121 30719
rect 23155 30716 23167 30719
rect 23382 30716 23388 30728
rect 23155 30688 23388 30716
rect 23155 30685 23167 30688
rect 23109 30679 23167 30685
rect 23382 30676 23388 30688
rect 23440 30676 23446 30728
rect 40586 30676 40592 30728
rect 40644 30676 40650 30728
rect 42794 30676 42800 30728
rect 42852 30716 42858 30728
rect 43622 30716 43628 30728
rect 42852 30688 43628 30716
rect 42852 30676 42858 30688
rect 43622 30676 43628 30688
rect 43680 30676 43686 30728
rect 32769 30651 32827 30657
rect 32769 30617 32781 30651
rect 32815 30648 32827 30651
rect 32858 30648 32864 30660
rect 32815 30620 32864 30648
rect 32815 30617 32827 30620
rect 32769 30611 32827 30617
rect 32858 30608 32864 30620
rect 32916 30608 32922 30660
rect 33502 30608 33508 30660
rect 33560 30608 33566 30660
rect 35434 30608 35440 30660
rect 35492 30608 35498 30660
rect 36265 30651 36323 30657
rect 36265 30617 36277 30651
rect 36311 30648 36323 30651
rect 37458 30648 37464 30660
rect 36311 30620 37464 30648
rect 36311 30617 36323 30620
rect 36265 30611 36323 30617
rect 37458 30608 37464 30620
rect 37516 30608 37522 30660
rect 41690 30608 41696 30660
rect 41748 30608 41754 30660
rect 38286 30540 38292 30592
rect 38344 30580 38350 30592
rect 40221 30583 40279 30589
rect 40221 30580 40233 30583
rect 38344 30552 40233 30580
rect 38344 30540 38350 30552
rect 40221 30549 40233 30552
rect 40267 30549 40279 30583
rect 40221 30543 40279 30549
rect 40681 30583 40739 30589
rect 40681 30549 40693 30583
rect 40727 30580 40739 30583
rect 48590 30580 48596 30592
rect 40727 30552 48596 30580
rect 40727 30549 40739 30552
rect 40681 30543 40739 30549
rect 48590 30540 48596 30552
rect 48648 30540 48654 30592
rect 1104 30490 49864 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 27950 30490
rect 28002 30438 28014 30490
rect 28066 30438 28078 30490
rect 28130 30438 28142 30490
rect 28194 30438 28206 30490
rect 28258 30438 37950 30490
rect 38002 30438 38014 30490
rect 38066 30438 38078 30490
rect 38130 30438 38142 30490
rect 38194 30438 38206 30490
rect 38258 30438 47950 30490
rect 48002 30438 48014 30490
rect 48066 30438 48078 30490
rect 48130 30438 48142 30490
rect 48194 30438 48206 30490
rect 48258 30438 49864 30490
rect 1104 30416 49864 30438
rect 39114 30336 39120 30388
rect 39172 30376 39178 30388
rect 39172 30348 39712 30376
rect 39172 30336 39178 30348
rect 34609 30311 34667 30317
rect 34609 30277 34621 30311
rect 34655 30308 34667 30311
rect 35437 30311 35495 30317
rect 35437 30308 35449 30311
rect 34655 30280 35449 30308
rect 34655 30277 34667 30280
rect 34609 30271 34667 30277
rect 35437 30277 35449 30280
rect 35483 30308 35495 30311
rect 35894 30308 35900 30320
rect 35483 30280 35900 30308
rect 35483 30277 35495 30280
rect 35437 30271 35495 30277
rect 35894 30268 35900 30280
rect 35952 30268 35958 30320
rect 38470 30308 38476 30320
rect 38120 30280 38476 30308
rect 35529 30243 35587 30249
rect 35529 30209 35541 30243
rect 35575 30240 35587 30243
rect 35986 30240 35992 30252
rect 35575 30212 35992 30240
rect 35575 30209 35587 30212
rect 35529 30203 35587 30209
rect 35986 30200 35992 30212
rect 36044 30200 36050 30252
rect 37458 30200 37464 30252
rect 37516 30240 37522 30252
rect 38120 30249 38148 30280
rect 38470 30268 38476 30280
rect 38528 30268 38534 30320
rect 39684 30308 39712 30348
rect 43254 30336 43260 30388
rect 43312 30376 43318 30388
rect 43530 30376 43536 30388
rect 43312 30348 43536 30376
rect 43312 30336 43318 30348
rect 43530 30336 43536 30348
rect 43588 30336 43594 30388
rect 40126 30308 40132 30320
rect 39606 30280 40132 30308
rect 40126 30268 40132 30280
rect 40184 30268 40190 30320
rect 41141 30311 41199 30317
rect 41141 30277 41153 30311
rect 41187 30308 41199 30311
rect 43272 30308 43300 30336
rect 41187 30280 43300 30308
rect 41187 30277 41199 30280
rect 41141 30271 41199 30277
rect 43622 30268 43628 30320
rect 43680 30268 43686 30320
rect 38105 30243 38163 30249
rect 38105 30240 38117 30243
rect 37516 30212 38117 30240
rect 37516 30200 37522 30212
rect 38105 30209 38117 30212
rect 38151 30209 38163 30243
rect 38105 30203 38163 30209
rect 39776 30212 41368 30240
rect 35618 30132 35624 30184
rect 35676 30132 35682 30184
rect 38381 30175 38439 30181
rect 38381 30141 38393 30175
rect 38427 30172 38439 30175
rect 39666 30172 39672 30184
rect 38427 30144 39672 30172
rect 38427 30141 38439 30144
rect 38381 30135 38439 30141
rect 39666 30132 39672 30144
rect 39724 30132 39730 30184
rect 39482 30064 39488 30116
rect 39540 30104 39546 30116
rect 39776 30104 39804 30212
rect 41340 30181 41368 30212
rect 41414 30200 41420 30252
rect 41472 30240 41478 30252
rect 42610 30240 42616 30252
rect 41472 30212 42616 30240
rect 41472 30200 41478 30212
rect 42610 30200 42616 30212
rect 42668 30200 42674 30252
rect 49326 30200 49332 30252
rect 49384 30200 49390 30252
rect 41233 30175 41291 30181
rect 41233 30141 41245 30175
rect 41279 30141 41291 30175
rect 41233 30135 41291 30141
rect 41325 30175 41383 30181
rect 41325 30141 41337 30175
rect 41371 30141 41383 30175
rect 41325 30135 41383 30141
rect 42889 30175 42947 30181
rect 42889 30141 42901 30175
rect 42935 30172 42947 30175
rect 42978 30172 42984 30184
rect 42935 30144 42984 30172
rect 42935 30141 42947 30144
rect 42889 30135 42947 30141
rect 39540 30076 39804 30104
rect 39540 30064 39546 30076
rect 34698 29996 34704 30048
rect 34756 30036 34762 30048
rect 35069 30039 35127 30045
rect 35069 30036 35081 30039
rect 34756 30008 35081 30036
rect 34756 29996 34762 30008
rect 35069 30005 35081 30008
rect 35115 30005 35127 30039
rect 35069 29999 35127 30005
rect 35158 29996 35164 30048
rect 35216 30036 35222 30048
rect 35802 30036 35808 30048
rect 35216 30008 35808 30036
rect 35216 29996 35222 30008
rect 35802 29996 35808 30008
rect 35860 30036 35866 30048
rect 39022 30036 39028 30048
rect 35860 30008 39028 30036
rect 35860 29996 35866 30008
rect 39022 29996 39028 30008
rect 39080 29996 39086 30048
rect 39758 29996 39764 30048
rect 39816 30036 39822 30048
rect 39853 30039 39911 30045
rect 39853 30036 39865 30039
rect 39816 30008 39865 30036
rect 39816 29996 39822 30008
rect 39853 30005 39865 30008
rect 39899 30005 39911 30039
rect 39853 29999 39911 30005
rect 40586 29996 40592 30048
rect 40644 30036 40650 30048
rect 40773 30039 40831 30045
rect 40773 30036 40785 30039
rect 40644 30008 40785 30036
rect 40644 29996 40650 30008
rect 40773 30005 40785 30008
rect 40819 30005 40831 30039
rect 41248 30036 41276 30135
rect 42978 30132 42984 30144
rect 43036 30172 43042 30184
rect 43530 30172 43536 30184
rect 43036 30144 43536 30172
rect 43036 30132 43042 30144
rect 43530 30132 43536 30144
rect 43588 30132 43594 30184
rect 41506 30036 41512 30048
rect 41248 30008 41512 30036
rect 40773 29999 40831 30005
rect 41506 29996 41512 30008
rect 41564 29996 41570 30048
rect 41690 29996 41696 30048
rect 41748 30036 41754 30048
rect 44361 30039 44419 30045
rect 44361 30036 44373 30039
rect 41748 30008 44373 30036
rect 41748 29996 41754 30008
rect 44361 30005 44373 30008
rect 44407 30005 44419 30039
rect 44361 29999 44419 30005
rect 48682 29996 48688 30048
rect 48740 30036 48746 30048
rect 49145 30039 49203 30045
rect 49145 30036 49157 30039
rect 48740 30008 49157 30036
rect 48740 29996 48746 30008
rect 49145 30005 49157 30008
rect 49191 30005 49203 30039
rect 49145 29999 49203 30005
rect 1104 29946 49864 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 32950 29946
rect 33002 29894 33014 29946
rect 33066 29894 33078 29946
rect 33130 29894 33142 29946
rect 33194 29894 33206 29946
rect 33258 29894 42950 29946
rect 43002 29894 43014 29946
rect 43066 29894 43078 29946
rect 43130 29894 43142 29946
rect 43194 29894 43206 29946
rect 43258 29894 49864 29946
rect 1104 29872 49864 29894
rect 31560 29835 31618 29841
rect 31560 29801 31572 29835
rect 31606 29832 31618 29835
rect 35618 29832 35624 29844
rect 31606 29804 35624 29832
rect 31606 29801 31618 29804
rect 31560 29795 31618 29801
rect 35618 29792 35624 29804
rect 35676 29792 35682 29844
rect 41506 29792 41512 29844
rect 41564 29832 41570 29844
rect 48958 29832 48964 29844
rect 41564 29804 48964 29832
rect 41564 29792 41570 29804
rect 48958 29792 48964 29804
rect 49016 29792 49022 29844
rect 34514 29724 34520 29776
rect 34572 29764 34578 29776
rect 35066 29764 35072 29776
rect 34572 29736 35072 29764
rect 34572 29724 34578 29736
rect 35066 29724 35072 29736
rect 35124 29764 35130 29776
rect 41598 29764 41604 29776
rect 35124 29736 41604 29764
rect 35124 29724 35130 29736
rect 41598 29724 41604 29736
rect 41656 29724 41662 29776
rect 48866 29764 48872 29776
rect 41800 29736 48872 29764
rect 33502 29696 33508 29708
rect 31312 29668 33508 29696
rect 22830 29588 22836 29640
rect 22888 29628 22894 29640
rect 31312 29637 31340 29668
rect 33502 29656 33508 29668
rect 33560 29656 33566 29708
rect 35526 29656 35532 29708
rect 35584 29656 35590 29708
rect 35894 29656 35900 29708
rect 35952 29696 35958 29708
rect 41506 29696 41512 29708
rect 35952 29668 41512 29696
rect 35952 29656 35958 29668
rect 41506 29656 41512 29668
rect 41564 29656 41570 29708
rect 31297 29631 31355 29637
rect 31297 29628 31309 29631
rect 22888 29600 31309 29628
rect 22888 29588 22894 29600
rect 31297 29597 31309 29600
rect 31343 29597 31355 29631
rect 31297 29591 31355 29597
rect 32674 29588 32680 29640
rect 32732 29588 32738 29640
rect 34606 29588 34612 29640
rect 34664 29628 34670 29640
rect 35345 29631 35403 29637
rect 35345 29628 35357 29631
rect 34664 29600 35357 29628
rect 34664 29588 34670 29600
rect 35345 29597 35357 29600
rect 35391 29628 35403 29631
rect 36173 29631 36231 29637
rect 36173 29628 36185 29631
rect 35391 29600 36185 29628
rect 35391 29597 35403 29600
rect 35345 29591 35403 29597
rect 36173 29597 36185 29600
rect 36219 29628 36231 29631
rect 41800 29628 41828 29736
rect 48866 29724 48872 29736
rect 48924 29724 48930 29776
rect 42610 29656 42616 29708
rect 42668 29696 42674 29708
rect 43533 29699 43591 29705
rect 43533 29696 43545 29699
rect 42668 29668 43545 29696
rect 42668 29656 42674 29668
rect 43533 29665 43545 29668
rect 43579 29665 43591 29699
rect 43533 29659 43591 29665
rect 48406 29628 48412 29640
rect 36219 29600 41828 29628
rect 41892 29600 48412 29628
rect 36219 29597 36231 29600
rect 36173 29591 36231 29597
rect 33318 29520 33324 29572
rect 33376 29560 33382 29572
rect 34057 29563 34115 29569
rect 34057 29560 34069 29563
rect 33376 29532 34069 29560
rect 33376 29520 33382 29532
rect 34057 29529 34069 29532
rect 34103 29560 34115 29563
rect 35253 29563 35311 29569
rect 35253 29560 35265 29563
rect 34103 29532 35265 29560
rect 34103 29529 34115 29532
rect 34057 29523 34115 29529
rect 35253 29529 35265 29532
rect 35299 29560 35311 29563
rect 41892 29560 41920 29600
rect 48406 29588 48412 29600
rect 48464 29588 48470 29640
rect 49326 29588 49332 29640
rect 49384 29588 49390 29640
rect 35299 29532 41920 29560
rect 35299 29529 35311 29532
rect 35253 29523 35311 29529
rect 41966 29520 41972 29572
rect 42024 29560 42030 29572
rect 42797 29563 42855 29569
rect 42797 29560 42809 29563
rect 42024 29532 42809 29560
rect 42024 29520 42030 29532
rect 42797 29529 42809 29532
rect 42843 29529 42855 29563
rect 50154 29560 50160 29572
rect 42797 29523 42855 29529
rect 42904 29532 50160 29560
rect 31662 29452 31668 29504
rect 31720 29492 31726 29504
rect 33045 29495 33103 29501
rect 33045 29492 33057 29495
rect 31720 29464 33057 29492
rect 31720 29452 31726 29464
rect 33045 29461 33057 29464
rect 33091 29461 33103 29495
rect 33045 29455 33103 29461
rect 33594 29452 33600 29504
rect 33652 29492 33658 29504
rect 34885 29495 34943 29501
rect 34885 29492 34897 29495
rect 33652 29464 34897 29492
rect 33652 29452 33658 29464
rect 34885 29461 34897 29464
rect 34931 29461 34943 29495
rect 34885 29455 34943 29461
rect 41506 29452 41512 29504
rect 41564 29492 41570 29504
rect 42904 29492 42932 29532
rect 50154 29520 50160 29532
rect 50212 29520 50218 29572
rect 41564 29464 42932 29492
rect 41564 29452 41570 29464
rect 48406 29452 48412 29504
rect 48464 29492 48470 29504
rect 49145 29495 49203 29501
rect 49145 29492 49157 29495
rect 48464 29464 49157 29492
rect 48464 29452 48470 29464
rect 49145 29461 49157 29464
rect 49191 29461 49203 29495
rect 49145 29455 49203 29461
rect 1104 29402 49864 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 27950 29402
rect 28002 29350 28014 29402
rect 28066 29350 28078 29402
rect 28130 29350 28142 29402
rect 28194 29350 28206 29402
rect 28258 29350 37950 29402
rect 38002 29350 38014 29402
rect 38066 29350 38078 29402
rect 38130 29350 38142 29402
rect 38194 29350 38206 29402
rect 38258 29350 47950 29402
rect 48002 29350 48014 29402
rect 48066 29350 48078 29402
rect 48130 29350 48142 29402
rect 48194 29350 48206 29402
rect 48258 29350 49864 29402
rect 1104 29328 49864 29350
rect 31386 29248 31392 29300
rect 31444 29288 31450 29300
rect 34241 29291 34299 29297
rect 34241 29288 34253 29291
rect 31444 29260 34253 29288
rect 31444 29248 31450 29260
rect 34241 29257 34253 29260
rect 34287 29257 34299 29291
rect 34241 29251 34299 29257
rect 34514 29248 34520 29300
rect 34572 29248 34578 29300
rect 34609 29291 34667 29297
rect 34609 29257 34621 29291
rect 34655 29288 34667 29291
rect 35250 29288 35256 29300
rect 34655 29260 35256 29288
rect 34655 29257 34667 29260
rect 34609 29251 34667 29257
rect 35250 29248 35256 29260
rect 35308 29288 35314 29300
rect 35529 29291 35587 29297
rect 35529 29288 35541 29291
rect 35308 29260 35541 29288
rect 35308 29248 35314 29260
rect 35529 29257 35541 29260
rect 35575 29288 35587 29291
rect 35575 29260 42564 29288
rect 35575 29257 35587 29260
rect 35529 29251 35587 29257
rect 32953 29223 33011 29229
rect 32953 29189 32965 29223
rect 32999 29220 33011 29223
rect 34532 29220 34560 29248
rect 32999 29192 34560 29220
rect 32999 29189 33011 29192
rect 32953 29183 33011 29189
rect 34790 29180 34796 29232
rect 34848 29180 34854 29232
rect 34882 29180 34888 29232
rect 34940 29220 34946 29232
rect 35802 29220 35808 29232
rect 34940 29192 35808 29220
rect 34940 29180 34946 29192
rect 35802 29180 35808 29192
rect 35860 29220 35866 29232
rect 36081 29223 36139 29229
rect 36081 29220 36093 29223
rect 35860 29192 36093 29220
rect 35860 29180 35866 29192
rect 36081 29189 36093 29192
rect 36127 29189 36139 29223
rect 39114 29220 39120 29232
rect 38962 29192 39120 29220
rect 36081 29183 36139 29189
rect 39114 29180 39120 29192
rect 39172 29180 39178 29232
rect 40034 29220 40040 29232
rect 39684 29192 40040 29220
rect 32861 29155 32919 29161
rect 32861 29121 32873 29155
rect 32907 29152 32919 29155
rect 34514 29152 34520 29164
rect 32907 29124 34520 29152
rect 32907 29121 32919 29124
rect 32861 29115 32919 29121
rect 34514 29112 34520 29124
rect 34572 29112 34578 29164
rect 34701 29155 34759 29161
rect 34701 29121 34713 29155
rect 34747 29152 34759 29155
rect 34808 29152 34836 29180
rect 35158 29152 35164 29164
rect 34747 29124 35164 29152
rect 34747 29121 34759 29124
rect 34701 29115 34759 29121
rect 30282 29044 30288 29096
rect 30340 29084 30346 29096
rect 33137 29087 33195 29093
rect 30340 29056 32904 29084
rect 30340 29044 30346 29056
rect 31570 28976 31576 29028
rect 31628 29016 31634 29028
rect 32493 29019 32551 29025
rect 32493 29016 32505 29019
rect 31628 28988 32505 29016
rect 31628 28976 31634 28988
rect 32493 28985 32505 28988
rect 32539 28985 32551 29019
rect 32876 29016 32904 29056
rect 33137 29053 33149 29087
rect 33183 29053 33195 29087
rect 33137 29047 33195 29053
rect 33781 29087 33839 29093
rect 33781 29053 33793 29087
rect 33827 29084 33839 29087
rect 34716 29084 34744 29115
rect 35158 29112 35164 29124
rect 35216 29112 35222 29164
rect 35989 29155 36047 29161
rect 35989 29121 36001 29155
rect 36035 29121 36047 29155
rect 35989 29115 36047 29121
rect 33827 29056 34744 29084
rect 34793 29087 34851 29093
rect 33827 29053 33839 29056
rect 33781 29047 33839 29053
rect 34793 29053 34805 29087
rect 34839 29053 34851 29087
rect 36004 29084 36032 29115
rect 37458 29112 37464 29164
rect 37516 29112 37522 29164
rect 39684 29161 39712 29192
rect 40034 29180 40040 29192
rect 40092 29180 40098 29232
rect 41414 29220 41420 29232
rect 41170 29192 41420 29220
rect 41414 29180 41420 29192
rect 41472 29180 41478 29232
rect 39669 29155 39727 29161
rect 39669 29121 39681 29155
rect 39715 29121 39727 29155
rect 39669 29115 39727 29121
rect 34793 29047 34851 29053
rect 35452 29056 36032 29084
rect 36173 29087 36231 29093
rect 33152 29016 33180 29047
rect 34808 29016 34836 29047
rect 32876 28988 34836 29016
rect 32493 28979 32551 28985
rect 34330 28908 34336 28960
rect 34388 28948 34394 28960
rect 35452 28948 35480 29056
rect 36173 29053 36185 29087
rect 36219 29053 36231 29087
rect 36173 29047 36231 29053
rect 39209 29087 39267 29093
rect 39209 29053 39221 29087
rect 39255 29084 39267 29087
rect 39942 29084 39948 29096
rect 39255 29056 39948 29084
rect 39255 29053 39267 29056
rect 39209 29047 39267 29053
rect 35621 29019 35679 29025
rect 35621 28985 35633 29019
rect 35667 29016 35679 29019
rect 35802 29016 35808 29028
rect 35667 28988 35808 29016
rect 35667 28985 35679 28988
rect 35621 28979 35679 28985
rect 35802 28976 35808 28988
rect 35860 28976 35866 29028
rect 34388 28920 35480 28948
rect 34388 28908 34394 28920
rect 35710 28908 35716 28960
rect 35768 28948 35774 28960
rect 36188 28948 36216 29047
rect 39942 29044 39948 29056
rect 40000 29044 40006 29096
rect 42536 29084 42564 29260
rect 43530 29248 43536 29300
rect 43588 29288 43594 29300
rect 44361 29291 44419 29297
rect 44361 29288 44373 29291
rect 43588 29260 44373 29288
rect 43588 29248 43594 29260
rect 44361 29257 44373 29260
rect 44407 29257 44419 29291
rect 44361 29251 44419 29257
rect 43622 29180 43628 29232
rect 43680 29180 43686 29232
rect 42610 29112 42616 29164
rect 42668 29112 42674 29164
rect 48498 29084 48504 29096
rect 42536 29056 48504 29084
rect 48498 29044 48504 29056
rect 48556 29044 48562 29096
rect 35768 28920 36216 28948
rect 37724 28951 37782 28957
rect 35768 28908 35774 28920
rect 37724 28917 37736 28951
rect 37770 28948 37782 28951
rect 38470 28948 38476 28960
rect 37770 28920 38476 28948
rect 37770 28917 37782 28920
rect 37724 28911 37782 28917
rect 38470 28908 38476 28920
rect 38528 28908 38534 28960
rect 39942 28908 39948 28960
rect 40000 28948 40006 28960
rect 41417 28951 41475 28957
rect 41417 28948 41429 28951
rect 40000 28920 41429 28948
rect 40000 28908 40006 28920
rect 41417 28917 41429 28920
rect 41463 28917 41475 28951
rect 41417 28911 41475 28917
rect 42426 28908 42432 28960
rect 42484 28948 42490 28960
rect 42870 28951 42928 28957
rect 42870 28948 42882 28951
rect 42484 28920 42882 28948
rect 42484 28908 42490 28920
rect 42870 28917 42882 28920
rect 42916 28917 42928 28951
rect 42870 28911 42928 28917
rect 1104 28858 49864 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 32950 28858
rect 33002 28806 33014 28858
rect 33066 28806 33078 28858
rect 33130 28806 33142 28858
rect 33194 28806 33206 28858
rect 33258 28806 42950 28858
rect 43002 28806 43014 28858
rect 43066 28806 43078 28858
rect 43130 28806 43142 28858
rect 43194 28806 43206 28858
rect 43258 28806 49864 28858
rect 1104 28784 49864 28806
rect 36173 28747 36231 28753
rect 36173 28713 36185 28747
rect 36219 28744 36231 28747
rect 42058 28744 42064 28756
rect 36219 28716 42064 28744
rect 36219 28713 36231 28716
rect 36173 28707 36231 28713
rect 30285 28611 30343 28617
rect 30285 28577 30297 28611
rect 30331 28608 30343 28611
rect 30650 28608 30656 28620
rect 30331 28580 30656 28608
rect 30331 28577 30343 28580
rect 30285 28571 30343 28577
rect 30650 28568 30656 28580
rect 30708 28608 30714 28620
rect 33229 28611 33287 28617
rect 33229 28608 33241 28611
rect 30708 28580 33241 28608
rect 30708 28568 30714 28580
rect 33229 28577 33241 28580
rect 33275 28577 33287 28611
rect 33229 28571 33287 28577
rect 35437 28611 35495 28617
rect 35437 28577 35449 28611
rect 35483 28608 35495 28611
rect 35526 28608 35532 28620
rect 35483 28580 35532 28608
rect 35483 28577 35495 28580
rect 35437 28571 35495 28577
rect 35452 28540 35480 28571
rect 35526 28568 35532 28580
rect 35584 28568 35590 28620
rect 36188 28608 36216 28707
rect 42058 28704 42064 28716
rect 42116 28704 42122 28756
rect 43622 28744 43628 28756
rect 42168 28716 43628 28744
rect 36004 28580 36216 28608
rect 32048 28512 35480 28540
rect 30466 28432 30472 28484
rect 30524 28472 30530 28484
rect 30561 28475 30619 28481
rect 30561 28472 30573 28475
rect 30524 28444 30573 28472
rect 30524 28432 30530 28444
rect 30561 28441 30573 28444
rect 30607 28441 30619 28475
rect 31938 28472 31944 28484
rect 31786 28444 31944 28472
rect 30561 28435 30619 28441
rect 31938 28432 31944 28444
rect 31996 28432 32002 28484
rect 32048 28416 32076 28512
rect 32493 28475 32551 28481
rect 32493 28441 32505 28475
rect 32539 28472 32551 28475
rect 32858 28472 32864 28484
rect 32539 28444 32864 28472
rect 32539 28441 32551 28444
rect 32493 28435 32551 28441
rect 32858 28432 32864 28444
rect 32916 28432 32922 28484
rect 33410 28432 33416 28484
rect 33468 28472 33474 28484
rect 35253 28475 35311 28481
rect 35253 28472 35265 28475
rect 33468 28444 35265 28472
rect 33468 28432 33474 28444
rect 35253 28441 35265 28444
rect 35299 28472 35311 28475
rect 36004 28472 36032 28580
rect 38470 28568 38476 28620
rect 38528 28608 38534 28620
rect 38749 28611 38807 28617
rect 38749 28608 38761 28611
rect 38528 28580 38761 28608
rect 38528 28568 38534 28580
rect 38749 28577 38761 28580
rect 38795 28577 38807 28611
rect 38749 28571 38807 28577
rect 36170 28500 36176 28552
rect 36228 28540 36234 28552
rect 37001 28543 37059 28549
rect 37001 28540 37013 28543
rect 36228 28512 37013 28540
rect 36228 28500 36234 28512
rect 37001 28509 37013 28512
rect 37047 28509 37059 28543
rect 39022 28540 39028 28552
rect 38410 28512 39028 28540
rect 37001 28503 37059 28509
rect 39022 28500 39028 28512
rect 39080 28500 39086 28552
rect 39390 28500 39396 28552
rect 39448 28500 39454 28552
rect 40034 28500 40040 28552
rect 40092 28500 40098 28552
rect 41414 28500 41420 28552
rect 41472 28540 41478 28552
rect 42168 28540 42196 28716
rect 43622 28704 43628 28716
rect 43680 28704 43686 28756
rect 42245 28611 42303 28617
rect 42245 28577 42257 28611
rect 42291 28608 42303 28611
rect 42610 28608 42616 28620
rect 42291 28580 42616 28608
rect 42291 28577 42303 28580
rect 42245 28571 42303 28577
rect 42610 28568 42616 28580
rect 42668 28568 42674 28620
rect 41472 28512 42196 28540
rect 41472 28500 41478 28512
rect 43622 28500 43628 28552
rect 43680 28500 43686 28552
rect 49326 28500 49332 28552
rect 49384 28500 49390 28552
rect 35299 28444 36032 28472
rect 37277 28475 37335 28481
rect 35299 28441 35311 28444
rect 35253 28435 35311 28441
rect 37277 28441 37289 28475
rect 37323 28441 37335 28475
rect 37277 28435 37335 28441
rect 32030 28364 32036 28416
rect 32088 28364 32094 28416
rect 34882 28364 34888 28416
rect 34940 28364 34946 28416
rect 35342 28364 35348 28416
rect 35400 28364 35406 28416
rect 37292 28404 37320 28435
rect 38838 28432 38844 28484
rect 38896 28472 38902 28484
rect 39942 28472 39948 28484
rect 38896 28444 39948 28472
rect 38896 28432 38902 28444
rect 39942 28432 39948 28444
rect 40000 28472 40006 28484
rect 40313 28475 40371 28481
rect 40313 28472 40325 28475
rect 40000 28444 40325 28472
rect 40000 28432 40006 28444
rect 40313 28441 40325 28444
rect 40359 28441 40371 28475
rect 42518 28472 42524 28484
rect 40313 28435 40371 28441
rect 41800 28444 42524 28472
rect 39482 28404 39488 28416
rect 37292 28376 39488 28404
rect 39482 28364 39488 28376
rect 39540 28364 39546 28416
rect 41800 28413 41828 28444
rect 42518 28432 42524 28444
rect 42576 28432 42582 28484
rect 41785 28407 41843 28413
rect 41785 28373 41797 28407
rect 41831 28373 41843 28407
rect 41785 28367 41843 28373
rect 42426 28364 42432 28416
rect 42484 28404 42490 28416
rect 43993 28407 44051 28413
rect 43993 28404 44005 28407
rect 42484 28376 44005 28404
rect 42484 28364 42490 28376
rect 43993 28373 44005 28376
rect 44039 28373 44051 28407
rect 43993 28367 44051 28373
rect 46934 28364 46940 28416
rect 46992 28404 46998 28416
rect 49145 28407 49203 28413
rect 49145 28404 49157 28407
rect 46992 28376 49157 28404
rect 46992 28364 46998 28376
rect 49145 28373 49157 28376
rect 49191 28373 49203 28407
rect 49145 28367 49203 28373
rect 1104 28314 49864 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 27950 28314
rect 28002 28262 28014 28314
rect 28066 28262 28078 28314
rect 28130 28262 28142 28314
rect 28194 28262 28206 28314
rect 28258 28262 37950 28314
rect 38002 28262 38014 28314
rect 38066 28262 38078 28314
rect 38130 28262 38142 28314
rect 38194 28262 38206 28314
rect 38258 28262 47950 28314
rect 48002 28262 48014 28314
rect 48066 28262 48078 28314
rect 48130 28262 48142 28314
rect 48194 28262 48206 28314
rect 48258 28262 49864 28314
rect 1104 28240 49864 28262
rect 22554 28160 22560 28212
rect 22612 28200 22618 28212
rect 23661 28203 23719 28209
rect 23661 28200 23673 28203
rect 22612 28172 23673 28200
rect 22612 28160 22618 28172
rect 23661 28169 23673 28172
rect 23707 28169 23719 28203
rect 30650 28200 30656 28212
rect 23661 28163 23719 28169
rect 28552 28172 30656 28200
rect 24029 28135 24087 28141
rect 24029 28101 24041 28135
rect 24075 28132 24087 28135
rect 25590 28132 25596 28144
rect 24075 28104 25596 28132
rect 24075 28101 24087 28104
rect 24029 28095 24087 28101
rect 25590 28092 25596 28104
rect 25648 28092 25654 28144
rect 24121 28067 24179 28073
rect 24121 28033 24133 28067
rect 24167 28064 24179 28067
rect 25498 28064 25504 28076
rect 24167 28036 25504 28064
rect 24167 28033 24179 28036
rect 24121 28027 24179 28033
rect 25498 28024 25504 28036
rect 25556 28024 25562 28076
rect 28442 28024 28448 28076
rect 28500 28064 28506 28076
rect 28552 28073 28580 28172
rect 30650 28160 30656 28172
rect 30708 28160 30714 28212
rect 31478 28160 31484 28212
rect 31536 28160 31542 28212
rect 32858 28160 32864 28212
rect 32916 28200 32922 28212
rect 38381 28203 38439 28209
rect 32916 28172 34836 28200
rect 32916 28160 32922 28172
rect 28810 28092 28816 28144
rect 28868 28092 28874 28144
rect 30098 28132 30104 28144
rect 30038 28104 30104 28132
rect 30098 28092 30104 28104
rect 30156 28132 30162 28144
rect 31938 28132 31944 28144
rect 30156 28104 31944 28132
rect 30156 28092 30162 28104
rect 31938 28092 31944 28104
rect 31996 28092 32002 28144
rect 33502 28132 33508 28144
rect 33244 28104 33508 28132
rect 33244 28073 33272 28104
rect 33502 28092 33508 28104
rect 33560 28092 33566 28144
rect 34808 28132 34836 28172
rect 38381 28169 38393 28203
rect 38427 28200 38439 28203
rect 39390 28200 39396 28212
rect 38427 28172 39396 28200
rect 38427 28169 38439 28172
rect 38381 28163 38439 28169
rect 39390 28160 39396 28172
rect 39448 28160 39454 28212
rect 40218 28160 40224 28212
rect 40276 28160 40282 28212
rect 43898 28200 43904 28212
rect 41708 28172 43904 28200
rect 35434 28141 35440 28144
rect 35425 28135 35440 28141
rect 35425 28132 35437 28135
rect 34808 28104 35437 28132
rect 35425 28101 35437 28104
rect 35425 28095 35440 28101
rect 35434 28092 35440 28095
rect 35492 28092 35498 28144
rect 39022 28132 39028 28144
rect 35544 28104 39028 28132
rect 28537 28067 28595 28073
rect 28537 28064 28549 28067
rect 28500 28036 28549 28064
rect 28500 28024 28506 28036
rect 28537 28033 28549 28036
rect 28583 28033 28595 28067
rect 28537 28027 28595 28033
rect 31389 28067 31447 28073
rect 31389 28033 31401 28067
rect 31435 28064 31447 28067
rect 33229 28067 33287 28073
rect 31435 28036 33180 28064
rect 31435 28033 31447 28036
rect 31389 28027 31447 28033
rect 24210 27956 24216 28008
rect 24268 27956 24274 28008
rect 27522 27956 27528 28008
rect 27580 27996 27586 28008
rect 31573 27999 31631 28005
rect 31573 27996 31585 27999
rect 27580 27968 31585 27996
rect 27580 27956 27586 27968
rect 31573 27965 31585 27968
rect 31619 27996 31631 27999
rect 31662 27996 31668 28008
rect 31619 27968 31668 27996
rect 31619 27965 31631 27968
rect 31573 27959 31631 27965
rect 31662 27956 31668 27968
rect 31720 27956 31726 28008
rect 31021 27931 31079 27937
rect 31021 27928 31033 27931
rect 29840 27900 31033 27928
rect 28902 27820 28908 27872
rect 28960 27860 28966 27872
rect 29840 27860 29868 27900
rect 31021 27897 31033 27900
rect 31067 27897 31079 27931
rect 31021 27891 31079 27897
rect 28960 27832 29868 27860
rect 28960 27820 28966 27832
rect 30282 27820 30288 27872
rect 30340 27820 30346 27872
rect 33152 27860 33180 28036
rect 33229 28033 33241 28067
rect 33275 28033 33287 28067
rect 33229 28027 33287 28033
rect 34606 28024 34612 28076
rect 34664 28064 34670 28076
rect 35544 28064 35572 28104
rect 39022 28092 39028 28104
rect 39080 28092 39086 28144
rect 34664 28036 35572 28064
rect 34664 28024 34670 28036
rect 38378 28024 38384 28076
rect 38436 28064 38442 28076
rect 38473 28067 38531 28073
rect 38473 28064 38485 28067
rect 38436 28036 38485 28064
rect 38436 28024 38442 28036
rect 38473 28033 38485 28036
rect 38519 28033 38531 28067
rect 38473 28027 38531 28033
rect 40129 28067 40187 28073
rect 40129 28033 40141 28067
rect 40175 28064 40187 28067
rect 40402 28064 40408 28076
rect 40175 28036 40408 28064
rect 40175 28033 40187 28036
rect 40129 28027 40187 28033
rect 40402 28024 40408 28036
rect 40460 28024 40466 28076
rect 41506 28024 41512 28076
rect 41564 28064 41570 28076
rect 41708 28073 41736 28172
rect 43898 28160 43904 28172
rect 43956 28160 43962 28212
rect 43993 28203 44051 28209
rect 43993 28169 44005 28203
rect 44039 28200 44051 28203
rect 46198 28200 46204 28212
rect 44039 28172 46204 28200
rect 44039 28169 44051 28172
rect 43993 28163 44051 28169
rect 46198 28160 46204 28172
rect 46256 28160 46262 28212
rect 41785 28135 41843 28141
rect 41785 28101 41797 28135
rect 41831 28132 41843 28135
rect 44174 28132 44180 28144
rect 41831 28104 44180 28132
rect 41831 28101 41843 28104
rect 41785 28095 41843 28101
rect 44174 28092 44180 28104
rect 44232 28092 44238 28144
rect 41693 28067 41751 28073
rect 41693 28064 41705 28067
rect 41564 28036 41705 28064
rect 41564 28024 41570 28036
rect 41693 28033 41705 28036
rect 41739 28033 41751 28067
rect 44358 28064 44364 28076
rect 41693 28027 41751 28033
rect 41800 28036 42012 28064
rect 33502 27956 33508 28008
rect 33560 27956 33566 28008
rect 36170 27956 36176 28008
rect 36228 27956 36234 28008
rect 38562 27956 38568 28008
rect 38620 27956 38626 28008
rect 40310 27956 40316 28008
rect 40368 27956 40374 28008
rect 35342 27888 35348 27940
rect 35400 27928 35406 27940
rect 35618 27928 35624 27940
rect 35400 27900 35624 27928
rect 35400 27888 35406 27900
rect 35618 27888 35624 27900
rect 35676 27928 35682 27940
rect 41800 27928 41828 28036
rect 41877 27999 41935 28005
rect 41877 27965 41889 27999
rect 41923 27965 41935 27999
rect 41984 27996 42012 28036
rect 44008 28036 44364 28064
rect 44008 27996 44036 28036
rect 44358 28024 44364 28036
rect 44416 28024 44422 28076
rect 49326 28024 49332 28076
rect 49384 28024 49390 28076
rect 41984 27968 44036 27996
rect 41877 27959 41935 27965
rect 35676 27900 41828 27928
rect 35676 27888 35682 27900
rect 34698 27860 34704 27872
rect 33152 27832 34704 27860
rect 34698 27820 34704 27832
rect 34756 27820 34762 27872
rect 34974 27820 34980 27872
rect 35032 27820 35038 27872
rect 37642 27820 37648 27872
rect 37700 27860 37706 27872
rect 38013 27863 38071 27869
rect 38013 27860 38025 27863
rect 37700 27832 38025 27860
rect 37700 27820 37706 27832
rect 38013 27829 38025 27832
rect 38059 27829 38071 27863
rect 38013 27823 38071 27829
rect 38378 27820 38384 27872
rect 38436 27860 38442 27872
rect 39761 27863 39819 27869
rect 39761 27860 39773 27863
rect 38436 27832 39773 27860
rect 38436 27820 38442 27832
rect 39761 27829 39773 27832
rect 39807 27829 39819 27863
rect 39761 27823 39819 27829
rect 39850 27820 39856 27872
rect 39908 27860 39914 27872
rect 41325 27863 41383 27869
rect 41325 27860 41337 27863
rect 39908 27832 41337 27860
rect 39908 27820 39914 27832
rect 41325 27829 41337 27832
rect 41371 27829 41383 27863
rect 41325 27823 41383 27829
rect 41782 27820 41788 27872
rect 41840 27860 41846 27872
rect 41892 27860 41920 27959
rect 44082 27956 44088 28008
rect 44140 27956 44146 28008
rect 42058 27888 42064 27940
rect 42116 27928 42122 27940
rect 49602 27928 49608 27940
rect 42116 27900 49608 27928
rect 42116 27888 42122 27900
rect 49602 27888 49608 27900
rect 49660 27888 49666 27940
rect 41840 27832 41920 27860
rect 41840 27820 41846 27832
rect 42610 27820 42616 27872
rect 42668 27860 42674 27872
rect 43533 27863 43591 27869
rect 43533 27860 43545 27863
rect 42668 27832 43545 27860
rect 42668 27820 42674 27832
rect 43533 27829 43545 27832
rect 43579 27829 43591 27863
rect 43533 27823 43591 27829
rect 48866 27820 48872 27872
rect 48924 27860 48930 27872
rect 49145 27863 49203 27869
rect 49145 27860 49157 27863
rect 48924 27832 49157 27860
rect 48924 27820 48930 27832
rect 49145 27829 49157 27832
rect 49191 27829 49203 27863
rect 49145 27823 49203 27829
rect 1104 27770 49864 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 32950 27770
rect 33002 27718 33014 27770
rect 33066 27718 33078 27770
rect 33130 27718 33142 27770
rect 33194 27718 33206 27770
rect 33258 27718 42950 27770
rect 43002 27718 43014 27770
rect 43066 27718 43078 27770
rect 43130 27718 43142 27770
rect 43194 27718 43206 27770
rect 43258 27718 49864 27770
rect 1104 27696 49864 27718
rect 24844 27659 24902 27665
rect 24844 27625 24856 27659
rect 24890 27656 24902 27659
rect 26142 27656 26148 27668
rect 24890 27628 26148 27656
rect 24890 27625 24902 27628
rect 24844 27619 24902 27625
rect 26142 27616 26148 27628
rect 26200 27616 26206 27668
rect 31008 27659 31066 27665
rect 31008 27625 31020 27659
rect 31054 27656 31066 27659
rect 32030 27656 32036 27668
rect 31054 27628 32036 27656
rect 31054 27625 31066 27628
rect 31008 27619 31066 27625
rect 32030 27616 32036 27628
rect 32088 27616 32094 27668
rect 32674 27656 32680 27668
rect 32140 27628 32680 27656
rect 24581 27523 24639 27529
rect 24581 27489 24593 27523
rect 24627 27520 24639 27523
rect 28442 27520 28448 27532
rect 24627 27492 28448 27520
rect 24627 27489 24639 27492
rect 24581 27483 24639 27489
rect 28442 27480 28448 27492
rect 28500 27480 28506 27532
rect 30650 27480 30656 27532
rect 30708 27520 30714 27532
rect 30745 27523 30803 27529
rect 30745 27520 30757 27523
rect 30708 27492 30757 27520
rect 30708 27480 30714 27492
rect 30745 27489 30757 27492
rect 30791 27489 30803 27523
rect 30745 27483 30803 27489
rect 32140 27464 32168 27628
rect 32674 27616 32680 27628
rect 32732 27656 32738 27668
rect 34606 27656 34612 27668
rect 32732 27628 34612 27656
rect 32732 27616 32738 27628
rect 34606 27616 34612 27628
rect 34664 27616 34670 27668
rect 40402 27616 40408 27668
rect 40460 27616 40466 27668
rect 32214 27548 32220 27600
rect 32272 27588 32278 27600
rect 37277 27591 37335 27597
rect 37277 27588 37289 27591
rect 32272 27560 37289 27588
rect 32272 27548 32278 27560
rect 37277 27557 37289 27560
rect 37323 27557 37335 27591
rect 37277 27551 37335 27557
rect 32493 27523 32551 27529
rect 32493 27489 32505 27523
rect 32539 27520 32551 27523
rect 33505 27523 33563 27529
rect 33505 27520 33517 27523
rect 32539 27492 33517 27520
rect 32539 27489 32551 27492
rect 32493 27483 32551 27489
rect 33505 27489 33517 27492
rect 33551 27489 33563 27523
rect 33505 27483 33563 27489
rect 32122 27412 32128 27464
rect 32180 27412 32186 27464
rect 24302 27344 24308 27396
rect 24360 27384 24366 27396
rect 24762 27384 24768 27396
rect 24360 27356 24768 27384
rect 24360 27344 24366 27356
rect 24762 27344 24768 27356
rect 24820 27384 24826 27396
rect 24820 27356 25346 27384
rect 24820 27344 24826 27356
rect 24210 27276 24216 27328
rect 24268 27316 24274 27328
rect 26329 27319 26387 27325
rect 26329 27316 26341 27319
rect 24268 27288 26341 27316
rect 24268 27276 24274 27288
rect 26329 27285 26341 27288
rect 26375 27285 26387 27319
rect 26329 27279 26387 27285
rect 30834 27276 30840 27328
rect 30892 27316 30898 27328
rect 32508 27316 32536 27483
rect 34974 27480 34980 27532
rect 35032 27520 35038 27532
rect 35710 27520 35716 27532
rect 35032 27492 35716 27520
rect 35032 27480 35038 27492
rect 35710 27480 35716 27492
rect 35768 27520 35774 27532
rect 36081 27523 36139 27529
rect 36081 27520 36093 27523
rect 35768 27492 36093 27520
rect 35768 27480 35774 27492
rect 36081 27489 36093 27492
rect 36127 27489 36139 27523
rect 36081 27483 36139 27489
rect 37921 27523 37979 27529
rect 37921 27489 37933 27523
rect 37967 27520 37979 27523
rect 39758 27520 39764 27532
rect 37967 27492 39764 27520
rect 37967 27489 37979 27492
rect 37921 27483 37979 27489
rect 39758 27480 39764 27492
rect 39816 27480 39822 27532
rect 43898 27480 43904 27532
rect 43956 27480 43962 27532
rect 33321 27455 33379 27461
rect 33321 27421 33333 27455
rect 33367 27452 33379 27455
rect 33367 27424 33456 27452
rect 33367 27421 33379 27424
rect 33321 27415 33379 27421
rect 33428 27384 33456 27424
rect 35894 27412 35900 27464
rect 35952 27412 35958 27464
rect 37645 27455 37703 27461
rect 37645 27421 37657 27455
rect 37691 27452 37703 27455
rect 38657 27455 38715 27461
rect 38657 27452 38669 27455
rect 37691 27424 38669 27452
rect 37691 27421 37703 27424
rect 37645 27415 37703 27421
rect 38657 27421 38669 27424
rect 38703 27421 38715 27455
rect 38657 27415 38715 27421
rect 41509 27455 41567 27461
rect 41509 27421 41521 27455
rect 41555 27452 41567 27455
rect 41690 27452 41696 27464
rect 41555 27424 41696 27452
rect 41555 27421 41567 27424
rect 41509 27415 41567 27421
rect 41690 27412 41696 27424
rect 41748 27412 41754 27464
rect 41966 27412 41972 27464
rect 42024 27412 42030 27464
rect 43714 27412 43720 27464
rect 43772 27412 43778 27464
rect 43809 27455 43867 27461
rect 43809 27421 43821 27455
rect 43855 27452 43867 27455
rect 46842 27452 46848 27464
rect 43855 27424 46848 27452
rect 43855 27421 43867 27424
rect 43809 27415 43867 27421
rect 46842 27412 46848 27424
rect 46900 27412 46906 27464
rect 33594 27384 33600 27396
rect 33428 27356 33600 27384
rect 33594 27344 33600 27356
rect 33652 27344 33658 27396
rect 37737 27387 37795 27393
rect 37737 27353 37749 27387
rect 37783 27384 37795 27387
rect 40954 27384 40960 27396
rect 37783 27356 40960 27384
rect 37783 27353 37795 27356
rect 37737 27347 37795 27353
rect 40954 27344 40960 27356
rect 41012 27344 41018 27396
rect 42702 27344 42708 27396
rect 42760 27344 42766 27396
rect 30892 27288 32536 27316
rect 32953 27319 33011 27325
rect 30892 27276 30898 27288
rect 32953 27285 32965 27319
rect 32999 27316 33011 27319
rect 33226 27316 33232 27328
rect 32999 27288 33232 27316
rect 32999 27285 33011 27288
rect 32953 27279 33011 27285
rect 33226 27276 33232 27288
rect 33284 27276 33290 27328
rect 33413 27319 33471 27325
rect 33413 27285 33425 27319
rect 33459 27316 33471 27319
rect 34882 27316 34888 27328
rect 33459 27288 34888 27316
rect 33459 27285 33471 27288
rect 33413 27279 33471 27285
rect 34882 27276 34888 27288
rect 34940 27276 34946 27328
rect 35526 27276 35532 27328
rect 35584 27276 35590 27328
rect 35986 27276 35992 27328
rect 36044 27276 36050 27328
rect 40494 27276 40500 27328
rect 40552 27316 40558 27328
rect 43349 27319 43407 27325
rect 43349 27316 43361 27319
rect 40552 27288 43361 27316
rect 40552 27276 40558 27288
rect 43349 27285 43361 27288
rect 43395 27285 43407 27319
rect 43349 27279 43407 27285
rect 1104 27226 49864 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 27950 27226
rect 28002 27174 28014 27226
rect 28066 27174 28078 27226
rect 28130 27174 28142 27226
rect 28194 27174 28206 27226
rect 28258 27174 37950 27226
rect 38002 27174 38014 27226
rect 38066 27174 38078 27226
rect 38130 27174 38142 27226
rect 38194 27174 38206 27226
rect 38258 27174 47950 27226
rect 48002 27174 48014 27226
rect 48066 27174 48078 27226
rect 48130 27174 48142 27226
rect 48194 27174 48206 27226
rect 48258 27174 49864 27226
rect 1104 27152 49864 27174
rect 30282 27112 30288 27124
rect 28736 27084 30288 27112
rect 28736 27053 28764 27084
rect 30282 27072 30288 27084
rect 30340 27072 30346 27124
rect 31386 27072 31392 27124
rect 31444 27072 31450 27124
rect 31481 27115 31539 27121
rect 31481 27081 31493 27115
rect 31527 27112 31539 27115
rect 31570 27112 31576 27124
rect 31527 27084 31576 27112
rect 31527 27081 31539 27084
rect 31481 27075 31539 27081
rect 31570 27072 31576 27084
rect 31628 27072 31634 27124
rect 33137 27115 33195 27121
rect 33137 27081 33149 27115
rect 33183 27112 33195 27115
rect 33318 27112 33324 27124
rect 33183 27084 33324 27112
rect 33183 27081 33195 27084
rect 33137 27075 33195 27081
rect 33318 27072 33324 27084
rect 33376 27112 33382 27124
rect 33594 27112 33600 27124
rect 33376 27084 33600 27112
rect 33376 27072 33382 27084
rect 33594 27072 33600 27084
rect 33652 27072 33658 27124
rect 35250 27072 35256 27124
rect 35308 27072 35314 27124
rect 39482 27072 39488 27124
rect 39540 27072 39546 27124
rect 41690 27072 41696 27124
rect 41748 27072 41754 27124
rect 41785 27115 41843 27121
rect 41785 27081 41797 27115
rect 41831 27112 41843 27115
rect 41874 27112 41880 27124
rect 41831 27084 41880 27112
rect 41831 27081 41843 27084
rect 41785 27075 41843 27081
rect 41874 27072 41880 27084
rect 41932 27072 41938 27124
rect 43806 27072 43812 27124
rect 43864 27112 43870 27124
rect 44637 27115 44695 27121
rect 44637 27112 44649 27115
rect 43864 27084 44649 27112
rect 43864 27072 43870 27084
rect 44637 27081 44649 27084
rect 44683 27081 44695 27115
rect 44637 27075 44695 27081
rect 44729 27115 44787 27121
rect 44729 27081 44741 27115
rect 44775 27112 44787 27115
rect 47394 27112 47400 27124
rect 44775 27084 47400 27112
rect 44775 27081 44787 27084
rect 44729 27075 44787 27081
rect 47394 27072 47400 27084
rect 47452 27072 47458 27124
rect 28721 27047 28779 27053
rect 28721 27013 28733 27047
rect 28767 27013 28779 27047
rect 30098 27044 30104 27056
rect 29946 27016 30104 27044
rect 28721 27007 28779 27013
rect 30098 27004 30104 27016
rect 30156 27004 30162 27056
rect 39022 27004 39028 27056
rect 39080 27004 39086 27056
rect 28442 26936 28448 26988
rect 28500 26936 28506 26988
rect 33229 26979 33287 26985
rect 33229 26945 33241 26979
rect 33275 26976 33287 26979
rect 34514 26976 34520 26988
rect 33275 26948 34520 26976
rect 33275 26945 33287 26948
rect 33229 26939 33287 26945
rect 34514 26936 34520 26948
rect 34572 26976 34578 26988
rect 34698 26976 34704 26988
rect 34572 26948 34704 26976
rect 34572 26936 34578 26948
rect 34698 26936 34704 26948
rect 34756 26936 34762 26988
rect 49326 26936 49332 26988
rect 49384 26936 49390 26988
rect 31573 26911 31631 26917
rect 31573 26908 31585 26911
rect 30024 26880 31585 26908
rect 27706 26800 27712 26852
rect 27764 26840 27770 26852
rect 27764 26812 28580 26840
rect 27764 26800 27770 26812
rect 24762 26732 24768 26784
rect 24820 26772 24826 26784
rect 28166 26772 28172 26784
rect 24820 26744 28172 26772
rect 24820 26732 24826 26744
rect 28166 26732 28172 26744
rect 28224 26732 28230 26784
rect 28552 26772 28580 26812
rect 30024 26772 30052 26880
rect 31573 26877 31585 26880
rect 31619 26877 31631 26911
rect 31573 26871 31631 26877
rect 32766 26868 32772 26920
rect 32824 26908 32830 26920
rect 33321 26911 33379 26917
rect 33321 26908 33333 26911
rect 32824 26880 33333 26908
rect 32824 26868 32830 26880
rect 33321 26877 33333 26880
rect 33367 26877 33379 26911
rect 33321 26871 33379 26877
rect 35158 26868 35164 26920
rect 35216 26908 35222 26920
rect 35345 26911 35403 26917
rect 35345 26908 35357 26911
rect 35216 26880 35357 26908
rect 35216 26868 35222 26880
rect 35345 26877 35357 26880
rect 35391 26877 35403 26911
rect 35345 26871 35403 26877
rect 35434 26868 35440 26920
rect 35492 26868 35498 26920
rect 36170 26868 36176 26920
rect 36228 26908 36234 26920
rect 37737 26911 37795 26917
rect 37737 26908 37749 26911
rect 36228 26880 37749 26908
rect 36228 26868 36234 26880
rect 37737 26877 37749 26880
rect 37783 26877 37795 26911
rect 37737 26871 37795 26877
rect 38013 26911 38071 26917
rect 38013 26877 38025 26911
rect 38059 26908 38071 26911
rect 39942 26908 39948 26920
rect 38059 26880 39948 26908
rect 38059 26877 38071 26880
rect 38013 26871 38071 26877
rect 39942 26868 39948 26880
rect 40000 26868 40006 26920
rect 41598 26868 41604 26920
rect 41656 26908 41662 26920
rect 41877 26911 41935 26917
rect 41877 26908 41889 26911
rect 41656 26880 41889 26908
rect 41656 26868 41662 26880
rect 41877 26877 41889 26880
rect 41923 26877 41935 26911
rect 41877 26871 41935 26877
rect 44913 26911 44971 26917
rect 44913 26877 44925 26911
rect 44959 26908 44971 26911
rect 45094 26908 45100 26920
rect 44959 26880 45100 26908
rect 44959 26877 44971 26880
rect 44913 26871 44971 26877
rect 45094 26868 45100 26880
rect 45152 26868 45158 26920
rect 30098 26800 30104 26852
rect 30156 26840 30162 26852
rect 30156 26812 31156 26840
rect 30156 26800 30162 26812
rect 30193 26775 30251 26781
rect 30193 26772 30205 26775
rect 28552 26744 30205 26772
rect 30193 26741 30205 26744
rect 30239 26741 30251 26775
rect 30193 26735 30251 26741
rect 30650 26732 30656 26784
rect 30708 26772 30714 26784
rect 31021 26775 31079 26781
rect 31021 26772 31033 26775
rect 30708 26744 31033 26772
rect 30708 26732 30714 26744
rect 31021 26741 31033 26744
rect 31067 26741 31079 26775
rect 31128 26772 31156 26812
rect 32674 26800 32680 26852
rect 32732 26840 32738 26852
rect 34885 26843 34943 26849
rect 34885 26840 34897 26843
rect 32732 26812 34897 26840
rect 32732 26800 32738 26812
rect 34885 26809 34897 26812
rect 34931 26809 34943 26843
rect 34885 26803 34943 26809
rect 32769 26775 32827 26781
rect 32769 26772 32781 26775
rect 31128 26744 32781 26772
rect 31021 26735 31079 26741
rect 32769 26741 32781 26744
rect 32815 26741 32827 26775
rect 32769 26735 32827 26741
rect 41138 26732 41144 26784
rect 41196 26772 41202 26784
rect 41325 26775 41383 26781
rect 41325 26772 41337 26775
rect 41196 26744 41337 26772
rect 41196 26732 41202 26744
rect 41325 26741 41337 26744
rect 41371 26741 41383 26775
rect 41325 26735 41383 26741
rect 43622 26732 43628 26784
rect 43680 26772 43686 26784
rect 44269 26775 44327 26781
rect 44269 26772 44281 26775
rect 43680 26744 44281 26772
rect 43680 26732 43686 26744
rect 44269 26741 44281 26744
rect 44315 26741 44327 26775
rect 44269 26735 44327 26741
rect 47026 26732 47032 26784
rect 47084 26772 47090 26784
rect 49145 26775 49203 26781
rect 49145 26772 49157 26775
rect 47084 26744 49157 26772
rect 47084 26732 47090 26744
rect 49145 26741 49157 26744
rect 49191 26741 49203 26775
rect 49145 26735 49203 26741
rect 1104 26682 49864 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 32950 26682
rect 33002 26630 33014 26682
rect 33066 26630 33078 26682
rect 33130 26630 33142 26682
rect 33194 26630 33206 26682
rect 33258 26630 42950 26682
rect 43002 26630 43014 26682
rect 43066 26630 43078 26682
rect 43130 26630 43142 26682
rect 43194 26630 43206 26682
rect 43258 26630 49864 26682
rect 1104 26608 49864 26630
rect 27338 26528 27344 26580
rect 27396 26568 27402 26580
rect 29181 26571 29239 26577
rect 27396 26540 29132 26568
rect 27396 26528 27402 26540
rect 29104 26500 29132 26540
rect 29181 26537 29193 26571
rect 29227 26568 29239 26571
rect 30466 26568 30472 26580
rect 29227 26540 30472 26568
rect 29227 26537 29239 26540
rect 29181 26531 29239 26537
rect 30466 26528 30472 26540
rect 30524 26528 30530 26580
rect 31478 26528 31484 26580
rect 31536 26568 31542 26580
rect 34885 26571 34943 26577
rect 34885 26568 34897 26571
rect 31536 26540 34897 26568
rect 31536 26528 31542 26540
rect 34885 26537 34897 26540
rect 34931 26537 34943 26571
rect 34885 26531 34943 26537
rect 29104 26472 30696 26500
rect 27430 26392 27436 26444
rect 27488 26432 27494 26444
rect 28442 26432 28448 26444
rect 27488 26404 28448 26432
rect 27488 26392 27494 26404
rect 28442 26392 28448 26404
rect 28500 26392 28506 26444
rect 30558 26392 30564 26444
rect 30616 26392 30622 26444
rect 30668 26432 30696 26472
rect 36262 26460 36268 26512
rect 36320 26500 36326 26512
rect 38197 26503 38255 26509
rect 38197 26500 38209 26503
rect 36320 26472 38209 26500
rect 36320 26460 36326 26472
rect 38197 26469 38209 26472
rect 38243 26469 38255 26503
rect 38197 26463 38255 26469
rect 41877 26503 41935 26509
rect 41877 26469 41889 26503
rect 41923 26500 41935 26503
rect 44082 26500 44088 26512
rect 41923 26472 44088 26500
rect 41923 26469 41935 26472
rect 41877 26463 41935 26469
rect 44082 26460 44088 26472
rect 44140 26460 44146 26512
rect 30834 26432 30840 26444
rect 30668 26404 30840 26432
rect 30834 26392 30840 26404
rect 30892 26392 30898 26444
rect 32309 26435 32367 26441
rect 32309 26401 32321 26435
rect 32355 26432 32367 26435
rect 33502 26432 33508 26444
rect 32355 26404 33508 26432
rect 32355 26401 32367 26404
rect 32309 26395 32367 26401
rect 33502 26392 33508 26404
rect 33560 26432 33566 26444
rect 34146 26432 34152 26444
rect 33560 26404 34152 26432
rect 33560 26392 33566 26404
rect 34146 26392 34152 26404
rect 34204 26392 34210 26444
rect 35066 26392 35072 26444
rect 35124 26432 35130 26444
rect 35345 26435 35403 26441
rect 35345 26432 35357 26435
rect 35124 26404 35357 26432
rect 35124 26392 35130 26404
rect 35345 26401 35357 26404
rect 35391 26401 35403 26435
rect 35345 26395 35403 26401
rect 35434 26392 35440 26444
rect 35492 26392 35498 26444
rect 38286 26392 38292 26444
rect 38344 26432 38350 26444
rect 38657 26435 38715 26441
rect 38657 26432 38669 26435
rect 38344 26404 38669 26432
rect 38344 26392 38350 26404
rect 38657 26401 38669 26404
rect 38703 26401 38715 26435
rect 38657 26395 38715 26401
rect 38838 26392 38844 26444
rect 38896 26392 38902 26444
rect 42702 26432 42708 26444
rect 40144 26404 42708 26432
rect 40144 26376 40172 26404
rect 42702 26392 42708 26404
rect 42760 26392 42766 26444
rect 42886 26392 42892 26444
rect 42944 26432 42950 26444
rect 43346 26432 43352 26444
rect 42944 26404 43352 26432
rect 42944 26392 42950 26404
rect 43346 26392 43352 26404
rect 43404 26392 43410 26444
rect 35250 26324 35256 26376
rect 35308 26324 35314 26376
rect 37737 26367 37795 26373
rect 37737 26333 37749 26367
rect 37783 26364 37795 26367
rect 38565 26367 38623 26373
rect 38565 26364 38577 26367
rect 37783 26336 38577 26364
rect 37783 26333 37795 26336
rect 37737 26327 37795 26333
rect 38565 26333 38577 26336
rect 38611 26333 38623 26367
rect 38565 26327 38623 26333
rect 40126 26324 40132 26376
rect 40184 26324 40190 26376
rect 42518 26324 42524 26376
rect 42576 26324 42582 26376
rect 48041 26367 48099 26373
rect 48041 26333 48053 26367
rect 48087 26364 48099 26367
rect 48498 26364 48504 26376
rect 48087 26336 48504 26364
rect 48087 26333 48099 26336
rect 48041 26327 48099 26333
rect 48498 26324 48504 26336
rect 48556 26324 48562 26376
rect 48590 26324 48596 26376
rect 48648 26364 48654 26376
rect 48777 26367 48835 26373
rect 48777 26364 48789 26367
rect 48648 26336 48789 26364
rect 48648 26324 48654 26336
rect 48777 26333 48789 26336
rect 48823 26333 48835 26367
rect 48777 26327 48835 26333
rect 25222 26256 25228 26308
rect 25280 26296 25286 26308
rect 27706 26296 27712 26308
rect 25280 26268 27712 26296
rect 25280 26256 25286 26268
rect 27706 26256 27712 26268
rect 27764 26256 27770 26308
rect 28166 26256 28172 26308
rect 28224 26256 28230 26308
rect 32122 26296 32128 26308
rect 32062 26268 32128 26296
rect 32122 26256 32128 26268
rect 32180 26256 32186 26308
rect 39758 26256 39764 26308
rect 39816 26296 39822 26308
rect 40405 26299 40463 26305
rect 40405 26296 40417 26299
rect 39816 26268 40417 26296
rect 39816 26256 39822 26268
rect 40405 26265 40417 26268
rect 40451 26265 40463 26299
rect 40405 26259 40463 26265
rect 40788 26268 40894 26296
rect 39022 26188 39028 26240
rect 39080 26228 39086 26240
rect 40788 26228 40816 26268
rect 43346 26256 43352 26308
rect 43404 26296 43410 26308
rect 43533 26299 43591 26305
rect 43533 26296 43545 26299
rect 43404 26268 43545 26296
rect 43404 26256 43410 26268
rect 43533 26265 43545 26268
rect 43579 26265 43591 26299
rect 43533 26259 43591 26265
rect 43717 26299 43775 26305
rect 43717 26265 43729 26299
rect 43763 26296 43775 26299
rect 45462 26296 45468 26308
rect 43763 26268 45468 26296
rect 43763 26265 43775 26268
rect 43717 26259 43775 26265
rect 45462 26256 45468 26268
rect 45520 26256 45526 26308
rect 41414 26228 41420 26240
rect 39080 26200 41420 26228
rect 39080 26188 39086 26200
rect 41414 26188 41420 26200
rect 41472 26188 41478 26240
rect 1104 26138 49864 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 27950 26138
rect 28002 26086 28014 26138
rect 28066 26086 28078 26138
rect 28130 26086 28142 26138
rect 28194 26086 28206 26138
rect 28258 26086 37950 26138
rect 38002 26086 38014 26138
rect 38066 26086 38078 26138
rect 38130 26086 38142 26138
rect 38194 26086 38206 26138
rect 38258 26086 47950 26138
rect 48002 26086 48014 26138
rect 48066 26086 48078 26138
rect 48130 26086 48142 26138
rect 48194 26086 48206 26138
rect 48258 26086 49864 26138
rect 1104 26064 49864 26086
rect 32030 25984 32036 26036
rect 32088 26024 32094 26036
rect 34885 26027 34943 26033
rect 34885 26024 34897 26027
rect 32088 25996 34897 26024
rect 32088 25984 32094 25996
rect 34885 25993 34897 25996
rect 34931 25993 34943 26027
rect 34885 25987 34943 25993
rect 27430 25956 27436 25968
rect 27172 25928 27436 25956
rect 27172 25897 27200 25928
rect 27430 25916 27436 25928
rect 27488 25916 27494 25968
rect 30469 25959 30527 25965
rect 30469 25925 30481 25959
rect 30515 25956 30527 25959
rect 31389 25959 31447 25965
rect 31389 25956 31401 25959
rect 30515 25928 31401 25956
rect 30515 25925 30527 25928
rect 30469 25919 30527 25925
rect 31389 25925 31401 25928
rect 31435 25956 31447 25959
rect 31846 25956 31852 25968
rect 31435 25928 31852 25956
rect 31435 25925 31447 25928
rect 31389 25919 31447 25925
rect 31846 25916 31852 25928
rect 31904 25956 31910 25968
rect 33042 25956 33048 25968
rect 31904 25928 33048 25956
rect 31904 25916 31910 25928
rect 33042 25916 33048 25928
rect 33100 25916 33106 25968
rect 34422 25916 34428 25968
rect 34480 25916 34486 25968
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 28534 25848 28540 25900
rect 28592 25848 28598 25900
rect 31297 25891 31355 25897
rect 31297 25857 31309 25891
rect 31343 25888 31355 25891
rect 32493 25891 32551 25897
rect 32493 25888 32505 25891
rect 31343 25860 32505 25888
rect 31343 25857 31355 25860
rect 31297 25851 31355 25857
rect 32493 25857 32505 25860
rect 32539 25857 32551 25891
rect 34900 25888 34928 25987
rect 35526 25984 35532 26036
rect 35584 26024 35590 26036
rect 35713 26027 35771 26033
rect 35713 26024 35725 26027
rect 35584 25996 35725 26024
rect 35584 25984 35590 25996
rect 35713 25993 35725 25996
rect 35759 25993 35771 26027
rect 35713 25987 35771 25993
rect 35802 25984 35808 26036
rect 35860 25984 35866 26036
rect 40126 26024 40132 26036
rect 38488 25996 40132 26024
rect 38488 25897 38516 25996
rect 40126 25984 40132 25996
rect 40184 25984 40190 26036
rect 41693 26027 41751 26033
rect 41693 25993 41705 26027
rect 41739 26024 41751 26027
rect 42518 26024 42524 26036
rect 41739 25996 42524 26024
rect 41739 25993 41751 25996
rect 41693 25987 41751 25993
rect 42518 25984 42524 25996
rect 42576 25984 42582 26036
rect 42702 26024 42708 26036
rect 42628 25996 42708 26024
rect 41414 25956 41420 25968
rect 39974 25928 41420 25956
rect 41414 25916 41420 25928
rect 41472 25956 41478 25968
rect 41874 25956 41880 25968
rect 41472 25928 41880 25956
rect 41472 25916 41478 25928
rect 41874 25916 41880 25928
rect 41932 25916 41938 25968
rect 42628 25897 42656 25996
rect 42702 25984 42708 25996
rect 42760 26024 42766 26036
rect 42760 25996 44864 26024
rect 42760 25984 42766 25996
rect 38473 25891 38531 25897
rect 34900 25860 35112 25888
rect 32493 25851 32551 25857
rect 26418 25780 26424 25832
rect 26476 25820 26482 25832
rect 27433 25823 27491 25829
rect 27433 25820 27445 25823
rect 26476 25792 27445 25820
rect 26476 25780 26482 25792
rect 27433 25789 27445 25792
rect 27479 25820 27491 25823
rect 27522 25820 27528 25832
rect 27479 25792 27528 25820
rect 27479 25789 27491 25792
rect 27433 25783 27491 25789
rect 27522 25780 27528 25792
rect 27580 25780 27586 25832
rect 31481 25823 31539 25829
rect 31481 25789 31493 25823
rect 31527 25789 31539 25823
rect 31481 25783 31539 25789
rect 33137 25823 33195 25829
rect 33137 25789 33149 25823
rect 33183 25789 33195 25823
rect 33137 25783 33195 25789
rect 33413 25823 33471 25829
rect 33413 25789 33425 25823
rect 33459 25820 33471 25823
rect 34974 25820 34980 25832
rect 33459 25792 34980 25820
rect 33459 25789 33471 25792
rect 33413 25783 33471 25789
rect 28718 25712 28724 25764
rect 28776 25752 28782 25764
rect 31496 25752 31524 25783
rect 28776 25724 31524 25752
rect 28776 25712 28782 25724
rect 28810 25644 28816 25696
rect 28868 25684 28874 25696
rect 28905 25687 28963 25693
rect 28905 25684 28917 25687
rect 28868 25656 28917 25684
rect 28868 25644 28874 25656
rect 28905 25653 28917 25656
rect 28951 25653 28963 25687
rect 28905 25647 28963 25653
rect 28994 25644 29000 25696
rect 29052 25684 29058 25696
rect 30929 25687 30987 25693
rect 30929 25684 30941 25687
rect 29052 25656 30941 25684
rect 29052 25644 29058 25656
rect 30929 25653 30941 25656
rect 30975 25653 30987 25687
rect 33152 25684 33180 25783
rect 34974 25780 34980 25792
rect 35032 25780 35038 25832
rect 35084 25820 35112 25860
rect 38473 25857 38485 25891
rect 38519 25857 38531 25891
rect 38473 25851 38531 25857
rect 42613 25891 42671 25897
rect 42613 25857 42625 25891
rect 42659 25857 42671 25891
rect 44358 25888 44364 25900
rect 44022 25860 44364 25888
rect 42613 25851 42671 25857
rect 44358 25848 44364 25860
rect 44416 25888 44422 25900
rect 44836 25897 44864 25996
rect 45094 25916 45100 25968
rect 45152 25916 45158 25968
rect 46106 25916 46112 25968
rect 46164 25916 46170 25968
rect 44821 25891 44879 25897
rect 44416 25860 44772 25888
rect 44416 25848 44422 25860
rect 35897 25823 35955 25829
rect 35897 25820 35909 25823
rect 35084 25792 35909 25820
rect 35897 25789 35909 25792
rect 35943 25789 35955 25823
rect 35897 25783 35955 25789
rect 38749 25823 38807 25829
rect 38749 25789 38761 25823
rect 38795 25820 38807 25823
rect 41690 25820 41696 25832
rect 38795 25792 41696 25820
rect 38795 25789 38807 25792
rect 38749 25783 38807 25789
rect 41690 25780 41696 25792
rect 41748 25780 41754 25832
rect 41785 25823 41843 25829
rect 41785 25789 41797 25823
rect 41831 25789 41843 25823
rect 41785 25783 41843 25789
rect 41969 25823 42027 25829
rect 41969 25789 41981 25823
rect 42015 25820 42027 25823
rect 42426 25820 42432 25832
rect 42015 25792 42432 25820
rect 42015 25789 42027 25792
rect 41969 25783 42027 25789
rect 36170 25752 36176 25764
rect 34808 25724 36176 25752
rect 33594 25684 33600 25696
rect 33152 25656 33600 25684
rect 30929 25647 30987 25653
rect 33594 25644 33600 25656
rect 33652 25684 33658 25696
rect 34808 25684 34836 25724
rect 36170 25712 36176 25724
rect 36228 25712 36234 25764
rect 39942 25712 39948 25764
rect 40000 25752 40006 25764
rect 40221 25755 40279 25761
rect 40221 25752 40233 25755
rect 40000 25724 40233 25752
rect 40000 25712 40006 25724
rect 40221 25721 40233 25724
rect 40267 25721 40279 25755
rect 40221 25715 40279 25721
rect 33652 25656 34836 25684
rect 33652 25644 33658 25656
rect 35342 25644 35348 25696
rect 35400 25644 35406 25696
rect 37734 25644 37740 25696
rect 37792 25684 37798 25696
rect 37921 25687 37979 25693
rect 37921 25684 37933 25687
rect 37792 25656 37933 25684
rect 37792 25644 37798 25656
rect 37921 25653 37933 25656
rect 37967 25653 37979 25687
rect 37921 25647 37979 25653
rect 40402 25644 40408 25696
rect 40460 25684 40466 25696
rect 41325 25687 41383 25693
rect 41325 25684 41337 25687
rect 40460 25656 41337 25684
rect 40460 25644 40466 25656
rect 41325 25653 41337 25656
rect 41371 25653 41383 25687
rect 41800 25684 41828 25783
rect 42426 25780 42432 25792
rect 42484 25780 42490 25832
rect 42889 25823 42947 25829
rect 42889 25789 42901 25823
rect 42935 25820 42947 25823
rect 43530 25820 43536 25832
rect 42935 25792 43536 25820
rect 42935 25789 42947 25792
rect 42889 25783 42947 25789
rect 43530 25780 43536 25792
rect 43588 25820 43594 25832
rect 44744 25820 44772 25860
rect 44821 25857 44833 25891
rect 44867 25857 44879 25891
rect 44821 25851 44879 25857
rect 46124 25820 46152 25916
rect 43588 25792 44496 25820
rect 44744 25792 46152 25820
rect 43588 25780 43594 25792
rect 43438 25684 43444 25696
rect 41800 25656 43444 25684
rect 41325 25647 41383 25653
rect 43438 25644 43444 25656
rect 43496 25644 43502 25696
rect 43990 25644 43996 25696
rect 44048 25684 44054 25696
rect 44361 25687 44419 25693
rect 44361 25684 44373 25687
rect 44048 25656 44373 25684
rect 44048 25644 44054 25656
rect 44361 25653 44373 25656
rect 44407 25653 44419 25687
rect 44468 25684 44496 25792
rect 46569 25687 46627 25693
rect 46569 25684 46581 25687
rect 44468 25656 46581 25684
rect 44361 25647 44419 25653
rect 46569 25653 46581 25656
rect 46615 25653 46627 25687
rect 46569 25647 46627 25653
rect 1104 25594 49864 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 32950 25594
rect 33002 25542 33014 25594
rect 33066 25542 33078 25594
rect 33130 25542 33142 25594
rect 33194 25542 33206 25594
rect 33258 25542 42950 25594
rect 43002 25542 43014 25594
rect 43066 25542 43078 25594
rect 43130 25542 43142 25594
rect 43194 25542 43206 25594
rect 43258 25542 49864 25594
rect 1104 25520 49864 25542
rect 24854 25440 24860 25492
rect 24912 25480 24918 25492
rect 28718 25480 28724 25492
rect 24912 25452 28724 25480
rect 24912 25440 24918 25452
rect 28718 25440 28724 25452
rect 28776 25440 28782 25492
rect 32490 25440 32496 25492
rect 32548 25480 32554 25492
rect 34885 25483 34943 25489
rect 34885 25480 34897 25483
rect 32548 25452 34897 25480
rect 32548 25440 32554 25452
rect 34885 25449 34897 25452
rect 34931 25449 34943 25483
rect 43993 25483 44051 25489
rect 43993 25480 44005 25483
rect 34885 25443 34943 25449
rect 41386 25452 44005 25480
rect 30466 25372 30472 25424
rect 30524 25412 30530 25424
rect 33597 25415 33655 25421
rect 30524 25384 30788 25412
rect 30524 25372 30530 25384
rect 30650 25304 30656 25356
rect 30708 25304 30714 25356
rect 30760 25353 30788 25384
rect 33597 25381 33609 25415
rect 33643 25412 33655 25415
rect 38562 25412 38568 25424
rect 33643 25384 38568 25412
rect 33643 25381 33655 25384
rect 33597 25375 33655 25381
rect 38562 25372 38568 25384
rect 38620 25372 38626 25424
rect 30745 25347 30803 25353
rect 30745 25313 30757 25347
rect 30791 25313 30803 25347
rect 30745 25307 30803 25313
rect 32766 25304 32772 25356
rect 32824 25344 32830 25356
rect 32950 25344 32956 25356
rect 32824 25316 32956 25344
rect 32824 25304 32830 25316
rect 32950 25304 32956 25316
rect 33008 25304 33014 25356
rect 33318 25304 33324 25356
rect 33376 25344 33382 25356
rect 34057 25347 34115 25353
rect 34057 25344 34069 25347
rect 33376 25316 34069 25344
rect 33376 25304 33382 25316
rect 34057 25313 34069 25316
rect 34103 25313 34115 25347
rect 34057 25307 34115 25313
rect 34146 25304 34152 25356
rect 34204 25304 34210 25356
rect 34514 25304 34520 25356
rect 34572 25344 34578 25356
rect 35437 25347 35495 25353
rect 35437 25344 35449 25347
rect 34572 25316 35449 25344
rect 34572 25304 34578 25316
rect 35437 25313 35449 25316
rect 35483 25313 35495 25347
rect 35437 25307 35495 25313
rect 38013 25347 38071 25353
rect 38013 25313 38025 25347
rect 38059 25344 38071 25347
rect 38470 25344 38476 25356
rect 38059 25316 38476 25344
rect 38059 25313 38071 25316
rect 38013 25307 38071 25313
rect 38470 25304 38476 25316
rect 38528 25304 38534 25356
rect 40313 25347 40371 25353
rect 40313 25313 40325 25347
rect 40359 25344 40371 25347
rect 40678 25344 40684 25356
rect 40359 25316 40684 25344
rect 40359 25313 40371 25316
rect 40313 25307 40371 25313
rect 40678 25304 40684 25316
rect 40736 25344 40742 25356
rect 41386 25344 41414 25452
rect 43993 25449 44005 25452
rect 44039 25449 44051 25483
rect 43993 25443 44051 25449
rect 41782 25372 41788 25424
rect 41840 25372 41846 25424
rect 43898 25372 43904 25424
rect 43956 25412 43962 25424
rect 45189 25415 45247 25421
rect 45189 25412 45201 25415
rect 43956 25384 45201 25412
rect 43956 25372 43962 25384
rect 45189 25381 45201 25384
rect 45235 25381 45247 25415
rect 45189 25375 45247 25381
rect 40736 25316 41414 25344
rect 42245 25347 42303 25353
rect 40736 25304 40742 25316
rect 42245 25313 42257 25347
rect 42291 25344 42303 25347
rect 44082 25344 44088 25356
rect 42291 25316 44088 25344
rect 42291 25313 42303 25316
rect 42245 25307 42303 25313
rect 44082 25304 44088 25316
rect 44140 25304 44146 25356
rect 45646 25304 45652 25356
rect 45704 25304 45710 25356
rect 45833 25347 45891 25353
rect 45833 25313 45845 25347
rect 45879 25344 45891 25347
rect 45922 25344 45928 25356
rect 45879 25316 45928 25344
rect 45879 25313 45891 25316
rect 45833 25307 45891 25313
rect 45922 25304 45928 25316
rect 45980 25304 45986 25356
rect 36909 25279 36967 25285
rect 36909 25276 36921 25279
rect 30208 25248 36921 25276
rect 30208 25149 30236 25248
rect 36909 25245 36921 25248
rect 36955 25245 36967 25279
rect 36909 25239 36967 25245
rect 37734 25236 37740 25288
rect 37792 25236 37798 25288
rect 40034 25236 40040 25288
rect 40092 25236 40098 25288
rect 44358 25276 44364 25288
rect 43654 25248 44364 25276
rect 44358 25236 44364 25248
rect 44416 25236 44422 25288
rect 45462 25236 45468 25288
rect 45520 25276 45526 25288
rect 47949 25279 48007 25285
rect 47949 25276 47961 25279
rect 45520 25248 47961 25276
rect 45520 25236 45526 25248
rect 47949 25245 47961 25248
rect 47995 25245 48007 25279
rect 47949 25239 48007 25245
rect 49142 25236 49148 25288
rect 49200 25236 49206 25288
rect 30374 25168 30380 25220
rect 30432 25208 30438 25220
rect 30432 25180 30696 25208
rect 30432 25168 30438 25180
rect 30193 25143 30251 25149
rect 30193 25109 30205 25143
rect 30239 25109 30251 25143
rect 30193 25103 30251 25109
rect 30558 25100 30564 25152
rect 30616 25100 30622 25152
rect 30668 25140 30696 25180
rect 31294 25168 31300 25220
rect 31352 25208 31358 25220
rect 31389 25211 31447 25217
rect 31389 25208 31401 25211
rect 31352 25180 31401 25208
rect 31352 25168 31358 25180
rect 31389 25177 31401 25180
rect 31435 25177 31447 25211
rect 33965 25211 34023 25217
rect 33965 25208 33977 25211
rect 31389 25171 31447 25177
rect 31496 25180 33977 25208
rect 31496 25140 31524 25180
rect 33965 25177 33977 25180
rect 34011 25177 34023 25211
rect 33965 25171 34023 25177
rect 35253 25211 35311 25217
rect 35253 25177 35265 25211
rect 35299 25208 35311 25211
rect 35894 25208 35900 25220
rect 35299 25180 35900 25208
rect 35299 25177 35311 25180
rect 35253 25171 35311 25177
rect 35894 25168 35900 25180
rect 35952 25168 35958 25220
rect 37829 25211 37887 25217
rect 37829 25177 37841 25211
rect 37875 25208 37887 25211
rect 40586 25208 40592 25220
rect 37875 25180 40592 25208
rect 37875 25177 37887 25180
rect 37829 25171 37887 25177
rect 40586 25168 40592 25180
rect 40644 25168 40650 25220
rect 41874 25208 41880 25220
rect 41538 25180 41880 25208
rect 41874 25168 41880 25180
rect 41932 25168 41938 25220
rect 42521 25211 42579 25217
rect 42521 25177 42533 25211
rect 42567 25177 42579 25211
rect 42521 25171 42579 25177
rect 30668 25112 31524 25140
rect 32858 25100 32864 25152
rect 32916 25100 32922 25152
rect 35066 25100 35072 25152
rect 35124 25140 35130 25152
rect 35345 25143 35403 25149
rect 35345 25140 35357 25143
rect 35124 25112 35357 25140
rect 35124 25100 35130 25112
rect 35345 25109 35357 25112
rect 35391 25140 35403 25143
rect 36630 25140 36636 25152
rect 35391 25112 36636 25140
rect 35391 25109 35403 25112
rect 35345 25103 35403 25109
rect 36630 25100 36636 25112
rect 36688 25100 36694 25152
rect 36722 25100 36728 25152
rect 36780 25100 36786 25152
rect 37366 25100 37372 25152
rect 37424 25100 37430 25152
rect 42536 25140 42564 25171
rect 43990 25140 43996 25152
rect 42536 25112 43996 25140
rect 43990 25100 43996 25112
rect 44048 25100 44054 25152
rect 45554 25100 45560 25152
rect 45612 25100 45618 25152
rect 1104 25050 49864 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 27950 25050
rect 28002 24998 28014 25050
rect 28066 24998 28078 25050
rect 28130 24998 28142 25050
rect 28194 24998 28206 25050
rect 28258 24998 37950 25050
rect 38002 24998 38014 25050
rect 38066 24998 38078 25050
rect 38130 24998 38142 25050
rect 38194 24998 38206 25050
rect 38258 24998 47950 25050
rect 48002 24998 48014 25050
rect 48066 24998 48078 25050
rect 48130 24998 48142 25050
rect 48194 24998 48206 25050
rect 48258 24998 49864 25050
rect 1104 24976 49864 24998
rect 31389 24939 31447 24945
rect 31389 24905 31401 24939
rect 31435 24936 31447 24939
rect 32674 24936 32680 24948
rect 31435 24908 32680 24936
rect 31435 24905 31447 24908
rect 31389 24899 31447 24905
rect 32674 24896 32680 24908
rect 32732 24896 32738 24948
rect 33410 24936 33416 24948
rect 32784 24908 33416 24936
rect 32784 24868 32812 24908
rect 33410 24896 33416 24908
rect 33468 24936 33474 24948
rect 34606 24936 34612 24948
rect 33468 24908 34612 24936
rect 33468 24896 33474 24908
rect 34606 24896 34612 24908
rect 34664 24896 34670 24948
rect 35894 24896 35900 24948
rect 35952 24936 35958 24948
rect 36538 24936 36544 24948
rect 35952 24908 36544 24936
rect 35952 24896 35958 24908
rect 36538 24896 36544 24908
rect 36596 24896 36602 24948
rect 36722 24896 36728 24948
rect 36780 24936 36786 24948
rect 43990 24936 43996 24948
rect 36780 24908 43996 24936
rect 36780 24896 36786 24908
rect 43990 24896 43996 24908
rect 44048 24896 44054 24948
rect 32692 24840 32812 24868
rect 31478 24760 31484 24812
rect 31536 24760 31542 24812
rect 32692 24809 32720 24840
rect 34422 24828 34428 24880
rect 34480 24828 34486 24880
rect 41874 24828 41880 24880
rect 41932 24868 41938 24880
rect 44358 24868 44364 24880
rect 41932 24840 44364 24868
rect 41932 24828 41938 24840
rect 44358 24828 44364 24840
rect 44416 24828 44422 24880
rect 46014 24868 46020 24880
rect 45678 24840 46020 24868
rect 46014 24828 46020 24840
rect 46072 24828 46078 24880
rect 32677 24803 32735 24809
rect 32677 24769 32689 24803
rect 32723 24769 32735 24803
rect 32677 24763 32735 24769
rect 36630 24760 36636 24812
rect 36688 24760 36694 24812
rect 37734 24760 37740 24812
rect 37792 24760 37798 24812
rect 38562 24760 38568 24812
rect 38620 24760 38626 24812
rect 41690 24760 41696 24812
rect 41748 24800 41754 24812
rect 42978 24800 42984 24812
rect 41748 24772 42984 24800
rect 41748 24760 41754 24772
rect 42978 24760 42984 24772
rect 43036 24760 43042 24812
rect 43073 24803 43131 24809
rect 43073 24769 43085 24803
rect 43119 24800 43131 24803
rect 43119 24772 43392 24800
rect 43119 24769 43131 24772
rect 43073 24763 43131 24769
rect 29454 24692 29460 24744
rect 29512 24732 29518 24744
rect 31573 24735 31631 24741
rect 31573 24732 31585 24735
rect 29512 24704 31585 24732
rect 29512 24692 29518 24704
rect 31573 24701 31585 24704
rect 31619 24732 31631 24735
rect 31619 24704 31754 24732
rect 31619 24701 31631 24704
rect 31573 24695 31631 24701
rect 31726 24664 31754 24704
rect 32582 24692 32588 24744
rect 32640 24732 32646 24744
rect 32769 24735 32827 24741
rect 32769 24732 32781 24735
rect 32640 24704 32781 24732
rect 32640 24692 32646 24704
rect 32769 24701 32781 24704
rect 32815 24701 32827 24735
rect 32769 24695 32827 24701
rect 32950 24692 32956 24744
rect 33008 24692 33014 24744
rect 33594 24692 33600 24744
rect 33652 24692 33658 24744
rect 33870 24692 33876 24744
rect 33928 24692 33934 24744
rect 36725 24735 36783 24741
rect 36725 24701 36737 24735
rect 36771 24701 36783 24735
rect 36725 24695 36783 24701
rect 43165 24735 43223 24741
rect 43165 24701 43177 24735
rect 43211 24701 43223 24735
rect 43165 24695 43223 24701
rect 33502 24664 33508 24676
rect 31726 24636 33508 24664
rect 33502 24624 33508 24636
rect 33560 24624 33566 24676
rect 34882 24624 34888 24676
rect 34940 24664 34946 24676
rect 36740 24664 36768 24695
rect 34940 24636 36768 24664
rect 34940 24624 34946 24636
rect 42058 24624 42064 24676
rect 42116 24664 42122 24676
rect 43180 24664 43208 24695
rect 42116 24636 43208 24664
rect 42116 24624 42122 24636
rect 27062 24556 27068 24608
rect 27120 24596 27126 24608
rect 28994 24596 29000 24608
rect 27120 24568 29000 24596
rect 27120 24556 27126 24568
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 31018 24556 31024 24608
rect 31076 24556 31082 24608
rect 31110 24556 31116 24608
rect 31168 24596 31174 24608
rect 32309 24599 32367 24605
rect 32309 24596 32321 24599
rect 31168 24568 32321 24596
rect 31168 24556 31174 24568
rect 32309 24565 32321 24568
rect 32355 24565 32367 24599
rect 32309 24559 32367 24565
rect 32398 24556 32404 24608
rect 32456 24596 32462 24608
rect 35345 24599 35403 24605
rect 35345 24596 35357 24599
rect 32456 24568 35357 24596
rect 32456 24556 32462 24568
rect 35345 24565 35357 24568
rect 35391 24596 35403 24599
rect 35434 24596 35440 24608
rect 35391 24568 35440 24596
rect 35391 24565 35403 24568
rect 35345 24559 35403 24565
rect 35434 24556 35440 24568
rect 35492 24556 35498 24608
rect 36173 24599 36231 24605
rect 36173 24565 36185 24599
rect 36219 24596 36231 24599
rect 36630 24596 36636 24608
rect 36219 24568 36636 24596
rect 36219 24565 36231 24568
rect 36173 24559 36231 24565
rect 36630 24556 36636 24568
rect 36688 24556 36694 24608
rect 37826 24556 37832 24608
rect 37884 24556 37890 24608
rect 38378 24556 38384 24608
rect 38436 24556 38442 24608
rect 39206 24556 39212 24608
rect 39264 24596 39270 24608
rect 42613 24599 42671 24605
rect 42613 24596 42625 24599
rect 39264 24568 42625 24596
rect 39264 24556 39270 24568
rect 42613 24565 42625 24568
rect 42659 24565 42671 24599
rect 43364 24596 43392 24772
rect 44082 24760 44088 24812
rect 44140 24800 44146 24812
rect 44177 24803 44235 24809
rect 44177 24800 44189 24803
rect 44140 24772 44189 24800
rect 44140 24760 44146 24772
rect 44177 24769 44189 24772
rect 44223 24769 44235 24803
rect 44177 24763 44235 24769
rect 45830 24760 45836 24812
rect 45888 24800 45894 24812
rect 47949 24803 48007 24809
rect 47949 24800 47961 24803
rect 45888 24772 47961 24800
rect 45888 24760 45894 24772
rect 47949 24769 47961 24772
rect 47995 24769 48007 24803
rect 47949 24763 48007 24769
rect 43438 24692 43444 24744
rect 43496 24732 43502 24744
rect 44453 24735 44511 24741
rect 44453 24732 44465 24735
rect 43496 24704 44465 24732
rect 43496 24692 43502 24704
rect 44453 24701 44465 24704
rect 44499 24701 44511 24735
rect 44453 24695 44511 24701
rect 45094 24692 45100 24744
rect 45152 24732 45158 24744
rect 45925 24735 45983 24741
rect 45925 24732 45937 24735
rect 45152 24704 45937 24732
rect 45152 24692 45158 24704
rect 45925 24701 45937 24704
rect 45971 24701 45983 24735
rect 45925 24695 45983 24701
rect 49142 24692 49148 24744
rect 49200 24692 49206 24744
rect 48406 24596 48412 24608
rect 43364 24568 48412 24596
rect 42613 24559 42671 24565
rect 48406 24556 48412 24568
rect 48464 24556 48470 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 22830 24352 22836 24404
rect 22888 24392 22894 24404
rect 25961 24395 26019 24401
rect 25961 24392 25973 24395
rect 22888 24364 25973 24392
rect 22888 24352 22894 24364
rect 25961 24361 25973 24364
rect 26007 24361 26019 24395
rect 25961 24355 26019 24361
rect 28445 24395 28503 24401
rect 28445 24361 28457 24395
rect 28491 24392 28503 24395
rect 28491 24364 36308 24392
rect 28491 24361 28503 24364
rect 28445 24355 28503 24361
rect 27154 24284 27160 24336
rect 27212 24324 27218 24336
rect 27212 24296 27660 24324
rect 27212 24284 27218 24296
rect 26605 24259 26663 24265
rect 26605 24225 26617 24259
rect 26651 24256 26663 24259
rect 27522 24256 27528 24268
rect 26651 24228 27528 24256
rect 26651 24225 26663 24228
rect 26605 24219 26663 24225
rect 27522 24216 27528 24228
rect 27580 24216 27586 24268
rect 27632 24256 27660 24296
rect 28810 24284 28816 24336
rect 28868 24324 28874 24336
rect 28868 24296 29040 24324
rect 28868 24284 28874 24296
rect 27632 24228 28856 24256
rect 26329 24123 26387 24129
rect 26329 24089 26341 24123
rect 26375 24120 26387 24123
rect 27798 24120 27804 24132
rect 26375 24092 27804 24120
rect 26375 24089 26387 24092
rect 26329 24083 26387 24089
rect 27798 24080 27804 24092
rect 27856 24080 27862 24132
rect 28828 24129 28856 24228
rect 28902 24216 28908 24268
rect 28960 24216 28966 24268
rect 29012 24265 29040 24296
rect 33502 24284 33508 24336
rect 33560 24324 33566 24336
rect 33689 24327 33747 24333
rect 33689 24324 33701 24327
rect 33560 24296 33701 24324
rect 33560 24284 33566 24296
rect 33689 24293 33701 24296
rect 33735 24293 33747 24327
rect 35618 24324 35624 24336
rect 33689 24287 33747 24293
rect 35360 24296 35624 24324
rect 28997 24259 29055 24265
rect 28997 24225 29009 24259
rect 29043 24225 29055 24259
rect 28997 24219 29055 24225
rect 30009 24259 30067 24265
rect 30009 24225 30021 24259
rect 30055 24256 30067 24259
rect 31202 24256 31208 24268
rect 30055 24228 31208 24256
rect 30055 24225 30067 24228
rect 30009 24219 30067 24225
rect 31202 24216 31208 24228
rect 31260 24216 31266 24268
rect 31941 24259 31999 24265
rect 31941 24225 31953 24259
rect 31987 24256 31999 24259
rect 33594 24256 33600 24268
rect 31987 24228 33600 24256
rect 31987 24225 31999 24228
rect 31941 24219 31999 24225
rect 33594 24216 33600 24228
rect 33652 24216 33658 24268
rect 35360 24265 35388 24296
rect 35618 24284 35624 24296
rect 35676 24284 35682 24336
rect 35345 24259 35403 24265
rect 35345 24225 35357 24259
rect 35391 24225 35403 24259
rect 35345 24219 35403 24225
rect 35437 24259 35495 24265
rect 35437 24225 35449 24259
rect 35483 24225 35495 24259
rect 35437 24219 35495 24225
rect 29730 24148 29736 24200
rect 29788 24148 29794 24200
rect 34422 24188 34428 24200
rect 33350 24160 34428 24188
rect 34422 24148 34428 24160
rect 34480 24148 34486 24200
rect 35250 24148 35256 24200
rect 35308 24148 35314 24200
rect 28813 24123 28871 24129
rect 28813 24089 28825 24123
rect 28859 24089 28871 24123
rect 31386 24120 31392 24132
rect 31234 24092 31392 24120
rect 28813 24083 28871 24089
rect 31386 24080 31392 24092
rect 31444 24120 31450 24132
rect 32122 24120 32128 24132
rect 31444 24092 32128 24120
rect 31444 24080 31450 24092
rect 32122 24080 32128 24092
rect 32180 24080 32186 24132
rect 32217 24123 32275 24129
rect 32217 24089 32229 24123
rect 32263 24120 32275 24123
rect 32306 24120 32312 24132
rect 32263 24092 32312 24120
rect 32263 24089 32275 24092
rect 32217 24083 32275 24089
rect 32306 24080 32312 24092
rect 32364 24080 32370 24132
rect 35452 24120 35480 24219
rect 36280 24197 36308 24364
rect 43162 24352 43168 24404
rect 43220 24392 43226 24404
rect 49510 24392 49516 24404
rect 43220 24364 49516 24392
rect 43220 24352 43226 24364
rect 49510 24352 49516 24364
rect 49568 24352 49574 24404
rect 38378 24284 38384 24336
rect 38436 24324 38442 24336
rect 46566 24324 46572 24336
rect 38436 24296 41414 24324
rect 38436 24284 38442 24296
rect 41386 24256 41414 24296
rect 42720 24296 46572 24324
rect 42720 24256 42748 24296
rect 46566 24284 46572 24296
rect 46624 24284 46630 24336
rect 41386 24228 42748 24256
rect 42794 24216 42800 24268
rect 42852 24256 42858 24268
rect 44085 24259 44143 24265
rect 44085 24256 44097 24259
rect 42852 24228 44097 24256
rect 42852 24216 42858 24228
rect 44085 24225 44097 24228
rect 44131 24225 44143 24259
rect 44085 24219 44143 24225
rect 45738 24216 45744 24268
rect 45796 24216 45802 24268
rect 48682 24256 48688 24268
rect 46492 24228 48688 24256
rect 36265 24191 36323 24197
rect 36265 24157 36277 24191
rect 36311 24157 36323 24191
rect 36265 24151 36323 24157
rect 38654 24148 38660 24200
rect 38712 24188 38718 24200
rect 38933 24191 38991 24197
rect 38933 24188 38945 24191
rect 38712 24160 38945 24188
rect 38712 24148 38718 24160
rect 38933 24157 38945 24160
rect 38979 24157 38991 24191
rect 38933 24151 38991 24157
rect 40310 24148 40316 24200
rect 40368 24188 40374 24200
rect 41693 24191 41751 24197
rect 41693 24188 41705 24191
rect 40368 24160 41705 24188
rect 40368 24148 40374 24160
rect 41693 24157 41705 24160
rect 41739 24157 41751 24191
rect 41693 24151 41751 24157
rect 43254 24148 43260 24200
rect 43312 24188 43318 24200
rect 43530 24188 43536 24200
rect 43312 24160 43536 24188
rect 43312 24148 43318 24160
rect 43530 24148 43536 24160
rect 43588 24148 43594 24200
rect 43806 24148 43812 24200
rect 43864 24188 43870 24200
rect 43901 24191 43959 24197
rect 43901 24188 43913 24191
rect 43864 24160 43913 24188
rect 43864 24148 43870 24160
rect 43901 24157 43913 24160
rect 43947 24157 43959 24191
rect 43901 24151 43959 24157
rect 43993 24191 44051 24197
rect 43993 24157 44005 24191
rect 44039 24188 44051 24191
rect 46492 24188 46520 24228
rect 48682 24216 48688 24228
rect 48740 24216 48746 24268
rect 44039 24160 46520 24188
rect 44039 24157 44051 24160
rect 43993 24151 44051 24157
rect 46566 24148 46572 24200
rect 46624 24148 46630 24200
rect 33520 24092 35480 24120
rect 26421 24055 26479 24061
rect 26421 24021 26433 24055
rect 26467 24052 26479 24055
rect 28626 24052 28632 24064
rect 26467 24024 28632 24052
rect 26467 24021 26479 24024
rect 26421 24015 26479 24021
rect 28626 24012 28632 24024
rect 28684 24012 28690 24064
rect 29362 24012 29368 24064
rect 29420 24052 29426 24064
rect 31481 24055 31539 24061
rect 31481 24052 31493 24055
rect 29420 24024 31493 24052
rect 29420 24012 29426 24024
rect 31481 24021 31493 24024
rect 31527 24052 31539 24055
rect 32582 24052 32588 24064
rect 31527 24024 32588 24052
rect 31527 24021 31539 24024
rect 31481 24015 31539 24021
rect 32582 24012 32588 24024
rect 32640 24012 32646 24064
rect 32950 24012 32956 24064
rect 33008 24052 33014 24064
rect 33520 24052 33548 24092
rect 37734 24080 37740 24132
rect 37792 24120 37798 24132
rect 43162 24120 43168 24132
rect 37792 24092 43168 24120
rect 37792 24080 37798 24092
rect 43162 24080 43168 24092
rect 43220 24080 43226 24132
rect 43714 24080 43720 24132
rect 43772 24120 43778 24132
rect 45557 24123 45615 24129
rect 45557 24120 45569 24123
rect 43772 24092 45569 24120
rect 43772 24080 43778 24092
rect 45557 24089 45569 24092
rect 45603 24089 45615 24123
rect 45557 24083 45615 24089
rect 45649 24123 45707 24129
rect 45649 24089 45661 24123
rect 45695 24120 45707 24123
rect 48314 24120 48320 24132
rect 45695 24092 48320 24120
rect 45695 24089 45707 24092
rect 45649 24083 45707 24089
rect 48314 24080 48320 24092
rect 48372 24080 48378 24132
rect 33008 24024 33548 24052
rect 33008 24012 33014 24024
rect 33778 24012 33784 24064
rect 33836 24052 33842 24064
rect 34885 24055 34943 24061
rect 34885 24052 34897 24055
rect 33836 24024 34897 24052
rect 33836 24012 33842 24024
rect 34885 24021 34897 24024
rect 34931 24021 34943 24055
rect 34885 24015 34943 24021
rect 36081 24055 36139 24061
rect 36081 24021 36093 24055
rect 36127 24052 36139 24055
rect 43346 24052 43352 24064
rect 36127 24024 43352 24052
rect 36127 24021 36139 24024
rect 36081 24015 36139 24021
rect 43346 24012 43352 24024
rect 43404 24012 43410 24064
rect 43530 24012 43536 24064
rect 43588 24012 43594 24064
rect 45186 24012 45192 24064
rect 45244 24012 45250 24064
rect 46382 24012 46388 24064
rect 46440 24012 46446 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 25590 23808 25596 23860
rect 25648 23808 25654 23860
rect 25961 23851 26019 23857
rect 25961 23817 25973 23851
rect 26007 23848 26019 23851
rect 27062 23848 27068 23860
rect 26007 23820 27068 23848
rect 26007 23817 26019 23820
rect 25961 23811 26019 23817
rect 27062 23808 27068 23820
rect 27120 23808 27126 23860
rect 29730 23848 29736 23860
rect 27172 23820 29736 23848
rect 27172 23721 27200 23820
rect 27157 23715 27215 23721
rect 27157 23681 27169 23715
rect 27203 23681 27215 23715
rect 27157 23675 27215 23681
rect 28534 23672 28540 23724
rect 28592 23672 28598 23724
rect 29472 23721 29500 23820
rect 29730 23808 29736 23820
rect 29788 23848 29794 23860
rect 29788 23820 31754 23848
rect 29788 23808 29794 23820
rect 31386 23780 31392 23792
rect 30958 23766 31392 23780
rect 30944 23752 31392 23766
rect 29457 23715 29515 23721
rect 29457 23681 29469 23715
rect 29503 23681 29515 23715
rect 29457 23675 29515 23681
rect 26050 23604 26056 23656
rect 26108 23604 26114 23656
rect 26142 23604 26148 23656
rect 26200 23604 26206 23656
rect 27433 23647 27491 23653
rect 27433 23613 27445 23647
rect 27479 23644 27491 23647
rect 29362 23644 29368 23656
rect 27479 23616 29368 23644
rect 27479 23613 27491 23616
rect 27433 23607 27491 23613
rect 29362 23604 29368 23616
rect 29420 23604 29426 23656
rect 29733 23647 29791 23653
rect 29733 23644 29745 23647
rect 29472 23616 29745 23644
rect 29472 23588 29500 23616
rect 29733 23613 29745 23616
rect 29779 23613 29791 23647
rect 29733 23607 29791 23613
rect 28534 23536 28540 23588
rect 28592 23576 28598 23588
rect 28994 23576 29000 23588
rect 28592 23548 29000 23576
rect 28592 23536 28598 23548
rect 28994 23536 29000 23548
rect 29052 23576 29058 23588
rect 29052 23548 29408 23576
rect 29052 23536 29058 23548
rect 28902 23468 28908 23520
rect 28960 23468 28966 23520
rect 29380 23508 29408 23548
rect 29454 23536 29460 23588
rect 29512 23536 29518 23588
rect 30944 23520 30972 23752
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 31726 23712 31754 23820
rect 32398 23808 32404 23860
rect 32456 23848 32462 23860
rect 32858 23848 32864 23860
rect 32456 23820 32864 23848
rect 32456 23808 32462 23820
rect 32858 23808 32864 23820
rect 32916 23848 32922 23860
rect 32916 23820 41184 23848
rect 32916 23808 32922 23820
rect 32030 23740 32036 23792
rect 32088 23780 32094 23792
rect 32585 23783 32643 23789
rect 32585 23780 32597 23783
rect 32088 23752 32597 23780
rect 32088 23740 32094 23752
rect 32585 23749 32597 23752
rect 32631 23749 32643 23783
rect 34422 23780 34428 23792
rect 33810 23752 34428 23780
rect 32585 23743 32643 23749
rect 34422 23740 34428 23752
rect 34480 23740 34486 23792
rect 34698 23740 34704 23792
rect 34756 23780 34762 23792
rect 34974 23780 34980 23792
rect 34756 23752 34980 23780
rect 34756 23740 34762 23752
rect 34974 23740 34980 23752
rect 35032 23780 35038 23792
rect 35032 23752 35204 23780
rect 35032 23740 35038 23752
rect 32309 23715 32367 23721
rect 32309 23712 32321 23715
rect 31726 23684 32321 23712
rect 32309 23681 32321 23684
rect 32355 23681 32367 23715
rect 32309 23675 32367 23681
rect 34790 23672 34796 23724
rect 34848 23672 34854 23724
rect 35176 23712 35204 23752
rect 35250 23740 35256 23792
rect 35308 23780 35314 23792
rect 36541 23783 36599 23789
rect 36541 23780 36553 23783
rect 35308 23752 36553 23780
rect 35308 23740 35314 23752
rect 36541 23749 36553 23752
rect 36587 23780 36599 23783
rect 36587 23752 38608 23780
rect 36587 23749 36599 23752
rect 36541 23743 36599 23749
rect 35345 23715 35403 23721
rect 35345 23712 35357 23715
rect 35176 23684 35357 23712
rect 35345 23681 35357 23684
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 37734 23672 37740 23724
rect 37792 23712 37798 23724
rect 37829 23715 37887 23721
rect 37829 23712 37841 23715
rect 37792 23684 37841 23712
rect 37792 23672 37798 23684
rect 37829 23681 37841 23684
rect 37875 23681 37887 23715
rect 38580 23712 38608 23752
rect 38654 23740 38660 23792
rect 38712 23740 38718 23792
rect 38749 23783 38807 23789
rect 38749 23749 38761 23783
rect 38795 23780 38807 23783
rect 39850 23780 39856 23792
rect 38795 23752 39856 23780
rect 38795 23749 38807 23752
rect 38749 23743 38807 23749
rect 39850 23740 39856 23752
rect 39908 23740 39914 23792
rect 40310 23740 40316 23792
rect 40368 23740 40374 23792
rect 40405 23783 40463 23789
rect 40405 23749 40417 23783
rect 40451 23780 40463 23783
rect 40494 23780 40500 23792
rect 40451 23752 40500 23780
rect 40451 23749 40463 23752
rect 40405 23743 40463 23749
rect 40494 23740 40500 23752
rect 40552 23740 40558 23792
rect 41156 23789 41184 23820
rect 41141 23783 41199 23789
rect 41141 23749 41153 23783
rect 41187 23780 41199 23783
rect 41966 23780 41972 23792
rect 41187 23752 41972 23780
rect 41187 23749 41199 23752
rect 41141 23743 41199 23749
rect 41966 23740 41972 23752
rect 42024 23780 42030 23792
rect 43257 23783 43315 23789
rect 43257 23780 43269 23783
rect 42024 23752 43269 23780
rect 42024 23740 42030 23752
rect 43257 23749 43269 23752
rect 43303 23749 43315 23783
rect 43257 23743 43315 23749
rect 44082 23740 44088 23792
rect 44140 23740 44146 23792
rect 39022 23712 39028 23724
rect 38580 23684 39028 23712
rect 37829 23675 37887 23681
rect 39022 23672 39028 23684
rect 39080 23672 39086 23724
rect 44100 23712 44128 23740
rect 44634 23712 44640 23724
rect 44100 23684 44640 23712
rect 44634 23672 44640 23684
rect 44692 23672 44698 23724
rect 46014 23672 46020 23724
rect 46072 23672 46078 23724
rect 46382 23672 46388 23724
rect 46440 23712 46446 23724
rect 47949 23715 48007 23721
rect 47949 23712 47961 23715
rect 46440 23684 47961 23712
rect 46440 23672 46446 23684
rect 47949 23681 47961 23684
rect 47995 23681 48007 23715
rect 47949 23675 48007 23681
rect 31202 23604 31208 23656
rect 31260 23604 31266 23656
rect 33870 23604 33876 23656
rect 33928 23644 33934 23656
rect 34057 23647 34115 23653
rect 34057 23644 34069 23647
rect 33928 23616 34069 23644
rect 33928 23604 33934 23616
rect 34057 23613 34069 23616
rect 34103 23613 34115 23647
rect 34808 23644 34836 23672
rect 35434 23644 35440 23656
rect 34808 23616 35440 23644
rect 34057 23607 34115 23613
rect 35434 23604 35440 23616
rect 35492 23604 35498 23656
rect 35529 23647 35587 23653
rect 35529 23613 35541 23647
rect 35575 23613 35587 23647
rect 35529 23607 35587 23613
rect 34790 23536 34796 23588
rect 34848 23576 34854 23588
rect 35544 23576 35572 23607
rect 35618 23604 35624 23656
rect 35676 23644 35682 23656
rect 36633 23647 36691 23653
rect 36633 23644 36645 23647
rect 35676 23616 36645 23644
rect 35676 23604 35682 23616
rect 36633 23613 36645 23616
rect 36679 23613 36691 23647
rect 36633 23607 36691 23613
rect 36817 23647 36875 23653
rect 36817 23613 36829 23647
rect 36863 23644 36875 23647
rect 36998 23644 37004 23656
rect 36863 23616 37004 23644
rect 36863 23613 36875 23616
rect 36817 23607 36875 23613
rect 34848 23548 35572 23576
rect 34848 23536 34854 23548
rect 30926 23508 30932 23520
rect 29380 23480 30932 23508
rect 30926 23468 30932 23480
rect 30984 23468 30990 23520
rect 32674 23468 32680 23520
rect 32732 23508 32738 23520
rect 32950 23508 32956 23520
rect 32732 23480 32956 23508
rect 32732 23468 32738 23480
rect 32950 23468 32956 23480
rect 33008 23468 33014 23520
rect 34977 23511 35035 23517
rect 34977 23477 34989 23511
rect 35023 23508 35035 23511
rect 35250 23508 35256 23520
rect 35023 23480 35256 23508
rect 35023 23477 35035 23480
rect 34977 23471 35035 23477
rect 35250 23468 35256 23480
rect 35308 23468 35314 23520
rect 35526 23468 35532 23520
rect 35584 23508 35590 23520
rect 36173 23511 36231 23517
rect 36173 23508 36185 23511
rect 35584 23480 36185 23508
rect 35584 23468 35590 23480
rect 36173 23477 36185 23480
rect 36219 23477 36231 23511
rect 36648 23508 36676 23607
rect 36998 23604 37004 23616
rect 37056 23604 37062 23656
rect 37550 23604 37556 23656
rect 37608 23644 37614 23656
rect 38933 23647 38991 23653
rect 37608 23616 38424 23644
rect 37608 23604 37614 23616
rect 36906 23536 36912 23588
rect 36964 23576 36970 23588
rect 38289 23579 38347 23585
rect 38289 23576 38301 23579
rect 36964 23548 38301 23576
rect 36964 23536 36970 23548
rect 38289 23545 38301 23548
rect 38335 23545 38347 23579
rect 38396 23576 38424 23616
rect 38933 23613 38945 23647
rect 38979 23644 38991 23647
rect 39942 23644 39948 23656
rect 38979 23616 39948 23644
rect 38979 23613 38991 23616
rect 38933 23607 38991 23613
rect 39942 23604 39948 23616
rect 40000 23604 40006 23656
rect 40589 23647 40647 23653
rect 40589 23613 40601 23647
rect 40635 23644 40647 23647
rect 40678 23644 40684 23656
rect 40635 23616 40684 23644
rect 40635 23613 40647 23616
rect 40589 23607 40647 23613
rect 40678 23604 40684 23616
rect 40736 23604 40742 23656
rect 41877 23647 41935 23653
rect 41877 23644 41889 23647
rect 41386 23616 41889 23644
rect 41386 23588 41414 23616
rect 41877 23613 41889 23616
rect 41923 23613 41935 23647
rect 41877 23607 41935 23613
rect 44913 23647 44971 23653
rect 44913 23613 44925 23647
rect 44959 23644 44971 23647
rect 45922 23644 45928 23656
rect 44959 23616 45928 23644
rect 44959 23613 44971 23616
rect 44913 23607 44971 23613
rect 45922 23604 45928 23616
rect 45980 23644 45986 23656
rect 46658 23644 46664 23656
rect 45980 23616 46664 23644
rect 45980 23604 45986 23616
rect 46658 23604 46664 23616
rect 46716 23604 46722 23656
rect 49142 23604 49148 23656
rect 49200 23604 49206 23656
rect 38396 23548 39988 23576
rect 38289 23539 38347 23545
rect 38838 23508 38844 23520
rect 36648 23480 38844 23508
rect 36173 23471 36231 23477
rect 38838 23468 38844 23480
rect 38896 23468 38902 23520
rect 39960 23517 39988 23548
rect 40034 23536 40040 23588
rect 40092 23576 40098 23588
rect 41322 23576 41328 23588
rect 40092 23548 41328 23576
rect 40092 23536 40098 23548
rect 41322 23536 41328 23548
rect 41380 23548 41414 23588
rect 41380 23536 41386 23548
rect 39945 23511 40003 23517
rect 39945 23477 39957 23511
rect 39991 23477 40003 23511
rect 39945 23471 40003 23477
rect 43438 23468 43444 23520
rect 43496 23508 43502 23520
rect 46385 23511 46443 23517
rect 46385 23508 46397 23511
rect 43496 23480 46397 23508
rect 43496 23468 43502 23480
rect 46385 23477 46397 23480
rect 46431 23477 46443 23511
rect 46385 23471 46443 23477
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 24026 23264 24032 23316
rect 24084 23304 24090 23316
rect 24084 23276 25912 23304
rect 24084 23264 24090 23276
rect 24854 23128 24860 23180
rect 24912 23168 24918 23180
rect 25406 23168 25412 23180
rect 24912 23140 25412 23168
rect 24912 23128 24918 23140
rect 25406 23128 25412 23140
rect 25464 23128 25470 23180
rect 25884 23168 25912 23276
rect 26142 23264 26148 23316
rect 26200 23304 26206 23316
rect 26329 23307 26387 23313
rect 26329 23304 26341 23307
rect 26200 23276 26341 23304
rect 26200 23264 26206 23276
rect 26329 23273 26341 23276
rect 26375 23273 26387 23307
rect 34974 23304 34980 23316
rect 26329 23267 26387 23273
rect 31312 23276 32076 23304
rect 28902 23168 28908 23180
rect 25884 23140 28908 23168
rect 28902 23128 28908 23140
rect 28960 23168 28966 23180
rect 30285 23171 30343 23177
rect 30285 23168 30297 23171
rect 28960 23140 30297 23168
rect 28960 23128 28966 23140
rect 30285 23137 30297 23140
rect 30331 23137 30343 23171
rect 30285 23131 30343 23137
rect 24578 23060 24584 23112
rect 24636 23060 24642 23112
rect 30098 23060 30104 23112
rect 30156 23060 30162 23112
rect 30193 23103 30251 23109
rect 30193 23069 30205 23103
rect 30239 23100 30251 23103
rect 31110 23100 31116 23112
rect 30239 23072 31116 23100
rect 30239 23069 30251 23072
rect 30193 23063 30251 23069
rect 31110 23060 31116 23072
rect 31168 23060 31174 23112
rect 31312 23109 31340 23276
rect 31404 23208 31754 23236
rect 31404 23177 31432 23208
rect 31389 23171 31447 23177
rect 31389 23137 31401 23171
rect 31435 23137 31447 23171
rect 31389 23131 31447 23137
rect 31481 23171 31539 23177
rect 31481 23137 31493 23171
rect 31527 23137 31539 23171
rect 31481 23131 31539 23137
rect 31297 23103 31355 23109
rect 31297 23069 31309 23103
rect 31343 23069 31355 23103
rect 31297 23063 31355 23069
rect 26602 23032 26608 23044
rect 26082 23004 26608 23032
rect 26602 22992 26608 23004
rect 26660 22992 26666 23044
rect 26694 22992 26700 23044
rect 26752 23032 26758 23044
rect 31496 23032 31524 23131
rect 31726 23100 31754 23208
rect 32048 23168 32076 23276
rect 32508 23276 34980 23304
rect 32508 23168 32536 23276
rect 34974 23264 34980 23276
rect 35032 23264 35038 23316
rect 40862 23264 40868 23316
rect 40920 23304 40926 23316
rect 43441 23307 43499 23313
rect 43441 23304 43453 23307
rect 40920 23276 43453 23304
rect 40920 23264 40926 23276
rect 43441 23273 43453 23276
rect 43487 23273 43499 23307
rect 43441 23267 43499 23273
rect 35434 23236 35440 23248
rect 32048 23140 32536 23168
rect 32692 23208 35440 23236
rect 32692 23100 32720 23208
rect 35434 23196 35440 23208
rect 35492 23196 35498 23248
rect 38105 23239 38163 23245
rect 38105 23205 38117 23239
rect 38151 23236 38163 23239
rect 39114 23236 39120 23248
rect 38151 23208 39120 23236
rect 38151 23205 38163 23208
rect 38105 23199 38163 23205
rect 39114 23196 39120 23208
rect 39172 23196 39178 23248
rect 42245 23239 42303 23245
rect 42245 23205 42257 23239
rect 42291 23236 42303 23239
rect 42794 23236 42800 23248
rect 42291 23208 42800 23236
rect 42291 23205 42303 23208
rect 42245 23199 42303 23205
rect 42794 23196 42800 23208
rect 42852 23196 42858 23248
rect 46934 23236 46940 23248
rect 43916 23208 46940 23236
rect 33410 23128 33416 23180
rect 33468 23128 33474 23180
rect 38378 23128 38384 23180
rect 38436 23168 38442 23180
rect 38749 23171 38807 23177
rect 38436 23140 38608 23168
rect 38436 23128 38442 23140
rect 31726 23072 32720 23100
rect 33229 23103 33287 23109
rect 33229 23069 33241 23103
rect 33275 23100 33287 23103
rect 34241 23103 34299 23109
rect 34241 23100 34253 23103
rect 33275 23072 34253 23100
rect 33275 23069 33287 23072
rect 33229 23063 33287 23069
rect 34241 23069 34253 23072
rect 34287 23069 34299 23103
rect 34241 23063 34299 23069
rect 37734 23060 37740 23112
rect 37792 23100 37798 23112
rect 38580 23109 38608 23140
rect 38749 23137 38761 23171
rect 38795 23168 38807 23171
rect 39298 23168 39304 23180
rect 38795 23140 39304 23168
rect 38795 23137 38807 23140
rect 38749 23131 38807 23137
rect 39298 23128 39304 23140
rect 39356 23128 39362 23180
rect 39408 23140 39620 23168
rect 38473 23103 38531 23109
rect 38473 23100 38485 23103
rect 37792 23072 38485 23100
rect 37792 23060 37798 23072
rect 38473 23069 38485 23072
rect 38519 23069 38531 23103
rect 38473 23063 38531 23069
rect 38565 23103 38623 23109
rect 38565 23069 38577 23103
rect 38611 23100 38623 23103
rect 39408 23100 39436 23140
rect 38611 23072 39436 23100
rect 39485 23103 39543 23109
rect 38611 23069 38623 23072
rect 38565 23063 38623 23069
rect 39485 23069 39497 23103
rect 39531 23069 39543 23103
rect 39592 23100 39620 23140
rect 40034 23128 40040 23180
rect 40092 23168 40098 23180
rect 40497 23171 40555 23177
rect 40497 23168 40509 23171
rect 40092 23140 40509 23168
rect 40092 23128 40098 23140
rect 40497 23137 40509 23140
rect 40543 23137 40555 23171
rect 40497 23131 40555 23137
rect 41506 23128 41512 23180
rect 41564 23168 41570 23180
rect 43916 23177 43944 23208
rect 46934 23196 46940 23208
rect 46992 23196 46998 23248
rect 43901 23171 43959 23177
rect 41564 23140 41920 23168
rect 41564 23128 41570 23140
rect 41892 23112 41920 23140
rect 43901 23137 43913 23171
rect 43947 23137 43959 23171
rect 43901 23131 43959 23137
rect 44085 23171 44143 23177
rect 44085 23137 44097 23171
rect 44131 23168 44143 23171
rect 44358 23168 44364 23180
rect 44131 23140 44364 23168
rect 44131 23137 44143 23140
rect 44085 23131 44143 23137
rect 44358 23128 44364 23140
rect 44416 23128 44422 23180
rect 40126 23100 40132 23112
rect 39592 23072 40132 23100
rect 39485 23063 39543 23069
rect 26752 23004 31524 23032
rect 32401 23035 32459 23041
rect 26752 22992 26758 23004
rect 32401 23001 32413 23035
rect 32447 23032 32459 23035
rect 32447 23004 33364 23032
rect 32447 23001 32459 23004
rect 32401 22995 32459 23001
rect 27246 22924 27252 22976
rect 27304 22964 27310 22976
rect 29733 22967 29791 22973
rect 29733 22964 29745 22967
rect 27304 22936 29745 22964
rect 27304 22924 27310 22936
rect 29733 22933 29745 22936
rect 29779 22933 29791 22967
rect 29733 22927 29791 22933
rect 30098 22924 30104 22976
rect 30156 22964 30162 22976
rect 30929 22967 30987 22973
rect 30929 22964 30941 22967
rect 30156 22936 30941 22964
rect 30156 22924 30162 22936
rect 30929 22933 30941 22936
rect 30975 22933 30987 22967
rect 30929 22927 30987 22933
rect 32214 22924 32220 22976
rect 32272 22964 32278 22976
rect 32490 22964 32496 22976
rect 32272 22936 32496 22964
rect 32272 22924 32278 22936
rect 32490 22924 32496 22936
rect 32548 22924 32554 22976
rect 32858 22924 32864 22976
rect 32916 22924 32922 22976
rect 33336 22973 33364 23004
rect 33502 22992 33508 23044
rect 33560 23032 33566 23044
rect 39500 23032 39528 23063
rect 40126 23060 40132 23072
rect 40184 23060 40190 23112
rect 41874 23060 41880 23112
rect 41932 23060 41938 23112
rect 42889 23103 42947 23109
rect 42889 23069 42901 23103
rect 42935 23100 42947 23103
rect 42978 23100 42984 23112
rect 42935 23072 42984 23100
rect 42935 23069 42947 23072
rect 42889 23063 42947 23069
rect 42978 23060 42984 23072
rect 43036 23060 43042 23112
rect 46109 23103 46167 23109
rect 46109 23100 46121 23103
rect 43088 23072 46121 23100
rect 33560 23004 39528 23032
rect 33560 22992 33566 23004
rect 40770 22992 40776 23044
rect 40828 22992 40834 23044
rect 43088 23032 43116 23072
rect 46109 23069 46121 23072
rect 46155 23069 46167 23103
rect 46109 23063 46167 23069
rect 47949 23103 48007 23109
rect 47949 23069 47961 23103
rect 47995 23069 48007 23103
rect 47949 23063 48007 23069
rect 42168 23004 43116 23032
rect 33321 22967 33379 22973
rect 33321 22933 33333 22967
rect 33367 22964 33379 22967
rect 34054 22964 34060 22976
rect 33367 22936 34060 22964
rect 33367 22933 33379 22936
rect 33321 22927 33379 22933
rect 34054 22924 34060 22936
rect 34112 22924 34118 22976
rect 39301 22967 39359 22973
rect 39301 22933 39313 22967
rect 39347 22964 39359 22967
rect 42168 22964 42196 23004
rect 43714 22992 43720 23044
rect 43772 23032 43778 23044
rect 43809 23035 43867 23041
rect 43809 23032 43821 23035
rect 43772 23004 43821 23032
rect 43772 22992 43778 23004
rect 43809 23001 43821 23004
rect 43855 23001 43867 23035
rect 43809 22995 43867 23001
rect 44174 22992 44180 23044
rect 44232 23032 44238 23044
rect 45281 23035 45339 23041
rect 45281 23032 45293 23035
rect 44232 23004 45293 23032
rect 44232 22992 44238 23004
rect 45281 23001 45293 23004
rect 45327 23001 45339 23035
rect 45281 22995 45339 23001
rect 45465 23035 45523 23041
rect 45465 23001 45477 23035
rect 45511 23032 45523 23035
rect 46750 23032 46756 23044
rect 45511 23004 46756 23032
rect 45511 23001 45523 23004
rect 45465 22995 45523 23001
rect 46750 22992 46756 23004
rect 46808 22992 46814 23044
rect 39347 22936 42196 22964
rect 45925 22967 45983 22973
rect 39347 22933 39359 22936
rect 39301 22927 39359 22933
rect 45925 22933 45937 22967
rect 45971 22964 45983 22967
rect 47964 22964 47992 23063
rect 49142 22992 49148 23044
rect 49200 22992 49206 23044
rect 45971 22936 47992 22964
rect 45971 22933 45983 22936
rect 45925 22927 45983 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 27614 22720 27620 22772
rect 27672 22760 27678 22772
rect 33410 22760 33416 22772
rect 27672 22732 33416 22760
rect 27672 22720 27678 22732
rect 33410 22720 33416 22732
rect 33468 22720 33474 22772
rect 33873 22763 33931 22769
rect 33873 22729 33885 22763
rect 33919 22760 33931 22763
rect 35342 22760 35348 22772
rect 33919 22732 35348 22760
rect 33919 22729 33931 22732
rect 33873 22723 33931 22729
rect 35342 22720 35348 22732
rect 35400 22720 35406 22772
rect 36538 22720 36544 22772
rect 36596 22760 36602 22772
rect 37829 22763 37887 22769
rect 37829 22760 37841 22763
rect 36596 22732 37841 22760
rect 36596 22720 36602 22732
rect 37829 22729 37841 22732
rect 37875 22729 37887 22763
rect 40034 22760 40040 22772
rect 37829 22723 37887 22729
rect 39040 22732 40040 22760
rect 36722 22652 36728 22704
rect 36780 22692 36786 22704
rect 37921 22695 37979 22701
rect 37921 22692 37933 22695
rect 36780 22664 37933 22692
rect 36780 22652 36786 22664
rect 37921 22661 37933 22664
rect 37967 22661 37979 22695
rect 37921 22655 37979 22661
rect 33410 22584 33416 22636
rect 33468 22624 33474 22636
rect 39040 22633 39068 22732
rect 40034 22720 40040 22732
rect 40092 22720 40098 22772
rect 40126 22720 40132 22772
rect 40184 22760 40190 22772
rect 41414 22760 41420 22772
rect 40184 22732 41420 22760
rect 40184 22720 40190 22732
rect 41414 22720 41420 22732
rect 41472 22720 41478 22772
rect 41601 22763 41659 22769
rect 41601 22729 41613 22763
rect 41647 22760 41659 22763
rect 41690 22760 41696 22772
rect 41647 22732 41696 22760
rect 41647 22729 41659 22732
rect 41601 22723 41659 22729
rect 41690 22720 41696 22732
rect 41748 22720 41754 22772
rect 42978 22720 42984 22772
rect 43036 22720 43042 22772
rect 43073 22763 43131 22769
rect 43073 22729 43085 22763
rect 43119 22760 43131 22763
rect 43622 22760 43628 22772
rect 43119 22732 43628 22760
rect 43119 22729 43131 22732
rect 43073 22723 43131 22729
rect 43622 22720 43628 22732
rect 43680 22720 43686 22772
rect 45830 22760 45836 22772
rect 44192 22732 45836 22760
rect 40586 22652 40592 22704
rect 40644 22692 40650 22704
rect 40644 22664 41828 22692
rect 40644 22652 40650 22664
rect 33781 22627 33839 22633
rect 33781 22624 33793 22627
rect 33468 22596 33793 22624
rect 33468 22584 33474 22596
rect 33781 22593 33793 22596
rect 33827 22593 33839 22627
rect 33781 22587 33839 22593
rect 39025 22627 39083 22633
rect 39025 22593 39037 22627
rect 39071 22593 39083 22627
rect 41506 22624 41512 22636
rect 40434 22596 41512 22624
rect 39025 22587 39083 22593
rect 41506 22584 41512 22596
rect 41564 22584 41570 22636
rect 33962 22516 33968 22568
rect 34020 22516 34026 22568
rect 38013 22559 38071 22565
rect 38013 22525 38025 22559
rect 38059 22525 38071 22559
rect 38013 22519 38071 22525
rect 33413 22491 33471 22497
rect 33413 22457 33425 22491
rect 33459 22488 33471 22491
rect 33502 22488 33508 22500
rect 33459 22460 33508 22488
rect 33459 22457 33471 22460
rect 33413 22451 33471 22457
rect 33502 22448 33508 22460
rect 33560 22448 33566 22500
rect 37734 22448 37740 22500
rect 37792 22488 37798 22500
rect 38028 22488 38056 22519
rect 39298 22516 39304 22568
rect 39356 22516 39362 22568
rect 39390 22516 39396 22568
rect 39448 22556 39454 22568
rect 40770 22556 40776 22568
rect 39448 22528 40776 22556
rect 39448 22516 39454 22528
rect 40770 22516 40776 22528
rect 40828 22516 40834 22568
rect 41800 22565 41828 22664
rect 43990 22652 43996 22704
rect 44048 22652 44054 22704
rect 44192 22701 44220 22732
rect 45830 22720 45836 22732
rect 45888 22720 45894 22772
rect 46658 22720 46664 22772
rect 46716 22720 46722 22772
rect 44177 22695 44235 22701
rect 44177 22661 44189 22695
rect 44223 22661 44235 22695
rect 44177 22655 44235 22661
rect 45922 22652 45928 22704
rect 45980 22652 45986 22704
rect 44634 22584 44640 22636
rect 44692 22624 44698 22636
rect 44910 22624 44916 22636
rect 44692 22596 44916 22624
rect 44692 22584 44698 22596
rect 44910 22584 44916 22596
rect 44968 22584 44974 22636
rect 41693 22559 41751 22565
rect 41693 22525 41705 22559
rect 41739 22525 41751 22559
rect 41693 22519 41751 22525
rect 41785 22559 41843 22565
rect 41785 22525 41797 22559
rect 41831 22525 41843 22559
rect 41785 22519 41843 22525
rect 43257 22559 43315 22565
rect 43257 22525 43269 22559
rect 43303 22556 43315 22559
rect 43346 22556 43352 22568
rect 43303 22528 43352 22556
rect 43303 22525 43315 22528
rect 43257 22519 43315 22525
rect 41233 22491 41291 22497
rect 41233 22488 41245 22491
rect 37792 22460 38056 22488
rect 40328 22460 41245 22488
rect 37792 22448 37798 22460
rect 37461 22423 37519 22429
rect 37461 22389 37473 22423
rect 37507 22420 37519 22423
rect 38470 22420 38476 22432
rect 37507 22392 38476 22420
rect 37507 22389 37519 22392
rect 37461 22383 37519 22389
rect 38470 22380 38476 22392
rect 38528 22380 38534 22432
rect 39666 22380 39672 22432
rect 39724 22420 39730 22432
rect 40328 22420 40356 22460
rect 41233 22457 41245 22460
rect 41279 22457 41291 22491
rect 41708 22488 41736 22519
rect 43346 22516 43352 22528
rect 43404 22516 43410 22568
rect 44542 22516 44548 22568
rect 44600 22556 44606 22568
rect 45189 22559 45247 22565
rect 45189 22556 45201 22559
rect 44600 22528 45201 22556
rect 44600 22516 44606 22528
rect 45189 22525 45201 22528
rect 45235 22525 45247 22559
rect 45189 22519 45247 22525
rect 41708 22460 42748 22488
rect 41233 22451 41291 22457
rect 39724 22392 40356 22420
rect 39724 22380 39730 22392
rect 40402 22380 40408 22432
rect 40460 22420 40466 22432
rect 42613 22423 42671 22429
rect 42613 22420 42625 22423
rect 40460 22392 42625 22420
rect 40460 22380 40466 22392
rect 42613 22389 42625 22392
rect 42659 22389 42671 22423
rect 42720 22420 42748 22460
rect 47026 22420 47032 22432
rect 42720 22392 47032 22420
rect 42613 22383 42671 22389
rect 47026 22380 47032 22392
rect 47084 22380 47090 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 30190 22225 30196 22228
rect 26040 22219 26098 22225
rect 26040 22185 26052 22219
rect 26086 22216 26098 22219
rect 30180 22219 30196 22225
rect 26086 22188 28488 22216
rect 26086 22185 26098 22188
rect 26040 22179 26098 22185
rect 24578 22108 24584 22160
rect 24636 22148 24642 22160
rect 28460 22148 28488 22188
rect 30180 22185 30192 22219
rect 30248 22216 30254 22228
rect 34514 22216 34520 22228
rect 30248 22188 34520 22216
rect 30180 22179 30196 22185
rect 30190 22176 30196 22179
rect 30248 22176 30254 22188
rect 34514 22176 34520 22188
rect 34572 22176 34578 22228
rect 39482 22176 39488 22228
rect 39540 22216 39546 22228
rect 40402 22216 40408 22228
rect 39540 22188 40408 22216
rect 39540 22176 39546 22188
rect 40402 22176 40408 22188
rect 40460 22176 40466 22228
rect 42600 22219 42658 22225
rect 42600 22185 42612 22219
rect 42646 22216 42658 22219
rect 42794 22216 42800 22228
rect 42646 22188 42800 22216
rect 42646 22185 42658 22188
rect 42600 22179 42658 22185
rect 42794 22176 42800 22188
rect 42852 22176 42858 22228
rect 29178 22148 29184 22160
rect 24636 22120 24808 22148
rect 28460 22120 29184 22148
rect 24636 22108 24642 22120
rect 24780 22080 24808 22120
rect 24780 22052 25452 22080
rect 25424 22024 25452 22052
rect 26786 22040 26792 22092
rect 26844 22080 26850 22092
rect 28552 22089 28580 22120
rect 29178 22108 29184 22120
rect 29236 22108 29242 22160
rect 29656 22120 30052 22148
rect 28445 22083 28503 22089
rect 28445 22080 28457 22083
rect 26844 22052 28457 22080
rect 26844 22040 26850 22052
rect 28445 22049 28457 22052
rect 28491 22049 28503 22083
rect 28445 22043 28503 22049
rect 28537 22083 28595 22089
rect 28537 22049 28549 22083
rect 28583 22080 28595 22083
rect 28583 22052 28617 22080
rect 28583 22049 28595 22052
rect 28537 22043 28595 22049
rect 25406 21972 25412 22024
rect 25464 22012 25470 22024
rect 25777 22015 25835 22021
rect 25777 22012 25789 22015
rect 25464 21984 25789 22012
rect 25464 21972 25470 21984
rect 25777 21981 25789 21984
rect 25823 21981 25835 22015
rect 25777 21975 25835 21981
rect 28353 22015 28411 22021
rect 28353 21981 28365 22015
rect 28399 22012 28411 22015
rect 29656 22012 29684 22120
rect 30024 22080 30052 22120
rect 33318 22108 33324 22160
rect 33376 22148 33382 22160
rect 33502 22148 33508 22160
rect 33376 22120 33508 22148
rect 33376 22108 33382 22120
rect 33502 22108 33508 22120
rect 33560 22108 33566 22160
rect 35894 22108 35900 22160
rect 35952 22148 35958 22160
rect 37553 22151 37611 22157
rect 35952 22120 36952 22148
rect 35952 22108 35958 22120
rect 32858 22080 32864 22092
rect 30024 22052 32864 22080
rect 32858 22040 32864 22052
rect 32916 22040 32922 22092
rect 35434 22040 35440 22092
rect 35492 22080 35498 22092
rect 36924 22089 36952 22120
rect 37553 22117 37565 22151
rect 37599 22148 37611 22151
rect 37599 22120 37633 22148
rect 37599 22117 37611 22120
rect 37553 22111 37611 22117
rect 36817 22083 36875 22089
rect 36817 22080 36829 22083
rect 35492 22052 36829 22080
rect 35492 22040 35498 22052
rect 36817 22049 36829 22052
rect 36863 22049 36875 22083
rect 36817 22043 36875 22049
rect 36909 22083 36967 22089
rect 36909 22049 36921 22083
rect 36955 22080 36967 22083
rect 37568 22080 37596 22111
rect 39298 22108 39304 22160
rect 39356 22148 39362 22160
rect 42058 22148 42064 22160
rect 39356 22120 42064 22148
rect 39356 22108 39362 22120
rect 42058 22108 42064 22120
rect 42116 22108 42122 22160
rect 36955 22052 36989 22080
rect 37568 22052 37872 22080
rect 36955 22049 36967 22052
rect 36909 22043 36967 22049
rect 28399 21984 29684 22012
rect 28399 21981 28411 21984
rect 28353 21975 28411 21981
rect 29730 21972 29736 22024
rect 29788 22012 29794 22024
rect 29917 22015 29975 22021
rect 29917 22012 29929 22015
rect 29788 21984 29929 22012
rect 29788 21972 29794 21984
rect 29917 21981 29929 21984
rect 29963 21981 29975 22015
rect 37737 22015 37795 22021
rect 37737 22012 37749 22015
rect 29917 21975 29975 21981
rect 31496 21984 37749 22012
rect 27062 21904 27068 21956
rect 27120 21904 27126 21956
rect 30926 21904 30932 21956
rect 30984 21904 30990 21956
rect 26418 21836 26424 21888
rect 26476 21876 26482 21888
rect 27522 21876 27528 21888
rect 26476 21848 27528 21876
rect 26476 21836 26482 21848
rect 27522 21836 27528 21848
rect 27580 21836 27586 21888
rect 27798 21836 27804 21888
rect 27856 21876 27862 21888
rect 27985 21879 28043 21885
rect 27985 21876 27997 21879
rect 27856 21848 27997 21876
rect 27856 21836 27862 21848
rect 27985 21845 27997 21848
rect 28031 21845 28043 21879
rect 27985 21839 28043 21845
rect 30834 21836 30840 21888
rect 30892 21876 30898 21888
rect 31496 21876 31524 21984
rect 37737 21981 37749 21984
rect 37783 21981 37795 22015
rect 37737 21975 37795 21981
rect 34974 21904 34980 21956
rect 35032 21944 35038 21956
rect 36725 21947 36783 21953
rect 36725 21944 36737 21947
rect 35032 21916 36737 21944
rect 35032 21904 35038 21916
rect 36725 21913 36737 21916
rect 36771 21913 36783 21947
rect 37274 21944 37280 21956
rect 36725 21907 36783 21913
rect 37108 21916 37280 21944
rect 30892 21848 31524 21876
rect 30892 21836 30898 21848
rect 31662 21836 31668 21888
rect 31720 21836 31726 21888
rect 36357 21879 36415 21885
rect 36357 21845 36369 21879
rect 36403 21876 36415 21879
rect 37108 21876 37136 21916
rect 37274 21904 37280 21916
rect 37332 21904 37338 21956
rect 37844 21944 37872 22052
rect 39206 22040 39212 22092
rect 39264 22040 39270 22092
rect 39390 22040 39396 22092
rect 39448 22040 39454 22092
rect 44174 22080 44180 22092
rect 39500 22052 44180 22080
rect 39114 21972 39120 22024
rect 39172 21972 39178 22024
rect 39500 21944 39528 22052
rect 44174 22040 44180 22052
rect 44232 22040 44238 22092
rect 45465 22083 45523 22089
rect 45465 22049 45477 22083
rect 45511 22080 45523 22083
rect 45554 22080 45560 22092
rect 45511 22052 45560 22080
rect 45511 22049 45523 22052
rect 45465 22043 45523 22049
rect 45554 22040 45560 22052
rect 45612 22040 45618 22092
rect 41322 21972 41328 22024
rect 41380 22012 41386 22024
rect 42337 22015 42395 22021
rect 42337 22012 42349 22015
rect 41380 21984 42349 22012
rect 41380 21972 41386 21984
rect 42337 21981 42349 21984
rect 42383 21981 42395 22015
rect 42337 21975 42395 21981
rect 44910 21972 44916 22024
rect 44968 22012 44974 22024
rect 45189 22015 45247 22021
rect 45189 22012 45201 22015
rect 44968 21984 45201 22012
rect 44968 21972 44974 21984
rect 45189 21981 45201 21984
rect 45235 21981 45247 22015
rect 45189 21975 45247 21981
rect 46750 21972 46756 22024
rect 46808 22012 46814 22024
rect 47949 22015 48007 22021
rect 47949 22012 47961 22015
rect 46808 21984 47961 22012
rect 46808 21972 46814 21984
rect 47949 21981 47961 21984
rect 47995 21981 48007 22015
rect 47949 21975 48007 21981
rect 49142 21972 49148 22024
rect 49200 21972 49206 22024
rect 37844 21916 39528 21944
rect 41598 21904 41604 21956
rect 41656 21944 41662 21956
rect 41656 21916 43102 21944
rect 41656 21904 41662 21916
rect 45922 21904 45928 21956
rect 45980 21904 45986 21956
rect 36403 21848 37136 21876
rect 36403 21845 36415 21848
rect 36357 21839 36415 21845
rect 37182 21836 37188 21888
rect 37240 21876 37246 21888
rect 38749 21879 38807 21885
rect 38749 21876 38761 21879
rect 37240 21848 38761 21876
rect 37240 21836 37246 21848
rect 38749 21845 38761 21848
rect 38795 21845 38807 21879
rect 38749 21839 38807 21845
rect 43898 21836 43904 21888
rect 43956 21876 43962 21888
rect 44085 21879 44143 21885
rect 44085 21876 44097 21879
rect 43956 21848 44097 21876
rect 43956 21836 43962 21848
rect 44085 21845 44097 21848
rect 44131 21845 44143 21879
rect 44085 21839 44143 21845
rect 44542 21836 44548 21888
rect 44600 21876 44606 21888
rect 46937 21879 46995 21885
rect 46937 21876 46949 21879
rect 44600 21848 46949 21876
rect 44600 21836 44606 21848
rect 46937 21845 46949 21848
rect 46983 21845 46995 21879
rect 46937 21839 46995 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 25498 21632 25504 21684
rect 25556 21632 25562 21684
rect 26602 21632 26608 21684
rect 26660 21672 26666 21684
rect 26878 21672 26884 21684
rect 26660 21644 26884 21672
rect 26660 21632 26666 21644
rect 26878 21632 26884 21644
rect 26936 21672 26942 21684
rect 27157 21675 27215 21681
rect 26936 21644 27108 21672
rect 26936 21632 26942 21644
rect 25961 21607 26019 21613
rect 25961 21573 25973 21607
rect 26007 21604 26019 21607
rect 26970 21604 26976 21616
rect 26007 21576 26976 21604
rect 26007 21573 26019 21576
rect 25961 21567 26019 21573
rect 26970 21564 26976 21576
rect 27028 21564 27034 21616
rect 27080 21604 27108 21644
rect 27157 21641 27169 21675
rect 27203 21672 27215 21675
rect 30374 21672 30380 21684
rect 27203 21644 30380 21672
rect 27203 21641 27215 21644
rect 27157 21635 27215 21641
rect 30374 21632 30380 21644
rect 30432 21632 30438 21684
rect 30653 21675 30711 21681
rect 30653 21641 30665 21675
rect 30699 21672 30711 21675
rect 30834 21672 30840 21684
rect 30699 21644 30840 21672
rect 30699 21641 30711 21644
rect 30653 21635 30711 21641
rect 30834 21632 30840 21644
rect 30892 21632 30898 21684
rect 31018 21632 31024 21684
rect 31076 21672 31082 21684
rect 31113 21675 31171 21681
rect 31113 21672 31125 21675
rect 31076 21644 31125 21672
rect 31076 21632 31082 21644
rect 31113 21641 31125 21644
rect 31159 21641 31171 21675
rect 31113 21635 31171 21641
rect 32766 21632 32772 21684
rect 32824 21672 32830 21684
rect 33045 21675 33103 21681
rect 33045 21672 33057 21675
rect 32824 21644 33057 21672
rect 32824 21632 32830 21644
rect 33045 21641 33057 21644
rect 33091 21641 33103 21675
rect 33045 21635 33103 21641
rect 37921 21675 37979 21681
rect 37921 21641 37933 21675
rect 37967 21672 37979 21675
rect 38378 21672 38384 21684
rect 37967 21644 38384 21672
rect 37967 21641 37979 21644
rect 37921 21635 37979 21641
rect 38378 21632 38384 21644
rect 38436 21632 38442 21684
rect 39022 21632 39028 21684
rect 39080 21632 39086 21684
rect 43165 21675 43223 21681
rect 43165 21641 43177 21675
rect 43211 21672 43223 21675
rect 43714 21672 43720 21684
rect 43211 21644 43720 21672
rect 43211 21641 43223 21644
rect 43165 21635 43223 21641
rect 43714 21632 43720 21644
rect 43772 21632 43778 21684
rect 43990 21632 43996 21684
rect 44048 21672 44054 21684
rect 44910 21672 44916 21684
rect 44048 21644 44916 21672
rect 44048 21632 44054 21644
rect 44910 21632 44916 21644
rect 44968 21632 44974 21684
rect 45738 21632 45744 21684
rect 45796 21632 45802 21684
rect 28994 21604 29000 21616
rect 27080 21576 29000 21604
rect 28994 21564 29000 21576
rect 29052 21604 29058 21616
rect 29052 21576 29210 21604
rect 29052 21564 29058 21576
rect 30466 21564 30472 21616
rect 30524 21604 30530 21616
rect 32953 21607 33011 21613
rect 32953 21604 32965 21607
rect 30524 21576 32965 21604
rect 30524 21564 30530 21576
rect 32953 21573 32965 21576
rect 32999 21573 33011 21607
rect 32953 21567 33011 21573
rect 34422 21564 34428 21616
rect 34480 21604 34486 21616
rect 35342 21604 35348 21616
rect 34480 21576 35348 21604
rect 34480 21564 34486 21576
rect 35342 21564 35348 21576
rect 35400 21604 35406 21616
rect 35400 21576 35558 21604
rect 35400 21564 35406 21576
rect 38838 21564 38844 21616
rect 38896 21604 38902 21616
rect 39117 21607 39175 21613
rect 39117 21604 39129 21607
rect 38896 21576 39129 21604
rect 38896 21564 38902 21576
rect 39117 21573 39129 21576
rect 39163 21573 39175 21607
rect 39117 21567 39175 21573
rect 43806 21564 43812 21616
rect 43864 21604 43870 21616
rect 44269 21607 44327 21613
rect 44269 21604 44281 21607
rect 43864 21576 44281 21604
rect 43864 21564 43870 21576
rect 44269 21573 44281 21576
rect 44315 21573 44327 21607
rect 45922 21604 45928 21616
rect 45494 21576 45928 21604
rect 44269 21567 44327 21573
rect 45922 21564 45928 21576
rect 45980 21564 45986 21616
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 25884 21400 25912 21499
rect 27522 21496 27528 21548
rect 27580 21496 27586 21548
rect 31021 21539 31079 21545
rect 31021 21505 31033 21539
rect 31067 21505 31079 21539
rect 31021 21499 31079 21505
rect 26142 21428 26148 21480
rect 26200 21428 26206 21480
rect 26510 21428 26516 21480
rect 26568 21468 26574 21480
rect 27617 21471 27675 21477
rect 27617 21468 27629 21471
rect 26568 21440 27629 21468
rect 26568 21428 26574 21440
rect 27617 21437 27629 21440
rect 27663 21437 27675 21471
rect 27617 21431 27675 21437
rect 27709 21471 27767 21477
rect 27709 21437 27721 21471
rect 27755 21437 27767 21471
rect 27709 21431 27767 21437
rect 26694 21400 26700 21412
rect 25884 21372 26700 21400
rect 26694 21360 26700 21372
rect 26752 21360 26758 21412
rect 27338 21360 27344 21412
rect 27396 21400 27402 21412
rect 27724 21400 27752 21431
rect 27798 21428 27804 21480
rect 27856 21468 27862 21480
rect 28445 21471 28503 21477
rect 28445 21468 28457 21471
rect 27856 21440 28457 21468
rect 27856 21428 27862 21440
rect 28445 21437 28457 21440
rect 28491 21437 28503 21471
rect 28445 21431 28503 21437
rect 28718 21428 28724 21480
rect 28776 21428 28782 21480
rect 31036 21468 31064 21499
rect 37826 21496 37832 21548
rect 37884 21496 37890 21548
rect 40586 21536 40592 21548
rect 38764 21508 40592 21536
rect 38764 21480 38792 21508
rect 40586 21496 40592 21508
rect 40644 21496 40650 21548
rect 43257 21539 43315 21545
rect 43257 21505 43269 21539
rect 43303 21536 43315 21539
rect 43303 21508 43944 21536
rect 43303 21505 43315 21508
rect 43257 21499 43315 21505
rect 29748 21440 31064 21468
rect 27396 21372 27752 21400
rect 27396 21360 27402 21372
rect 24946 21292 24952 21344
rect 25004 21292 25010 21344
rect 25130 21292 25136 21344
rect 25188 21332 25194 21344
rect 29748 21332 29776 21440
rect 31202 21428 31208 21480
rect 31260 21428 31266 21480
rect 33137 21471 33195 21477
rect 33137 21437 33149 21471
rect 33183 21437 33195 21471
rect 33137 21431 33195 21437
rect 31018 21360 31024 21412
rect 31076 21400 31082 21412
rect 31662 21400 31668 21412
rect 31076 21372 31668 21400
rect 31076 21360 31082 21372
rect 31662 21360 31668 21372
rect 31720 21400 31726 21412
rect 33152 21400 33180 21431
rect 34514 21428 34520 21480
rect 34572 21468 34578 21480
rect 34793 21471 34851 21477
rect 34793 21468 34805 21471
rect 34572 21440 34805 21468
rect 34572 21428 34578 21440
rect 34793 21437 34805 21440
rect 34839 21437 34851 21471
rect 34793 21431 34851 21437
rect 35066 21428 35072 21480
rect 35124 21468 35130 21480
rect 35434 21468 35440 21480
rect 35124 21440 35440 21468
rect 35124 21428 35130 21440
rect 35434 21428 35440 21440
rect 35492 21428 35498 21480
rect 38105 21471 38163 21477
rect 38105 21437 38117 21471
rect 38151 21468 38163 21471
rect 38746 21468 38752 21480
rect 38151 21440 38752 21468
rect 38151 21437 38163 21440
rect 38105 21431 38163 21437
rect 38746 21428 38752 21440
rect 38804 21428 38810 21480
rect 39022 21428 39028 21480
rect 39080 21468 39086 21480
rect 39209 21471 39267 21477
rect 39209 21468 39221 21471
rect 39080 21440 39221 21468
rect 39080 21428 39086 21440
rect 39209 21437 39221 21440
rect 39255 21437 39267 21471
rect 39209 21431 39267 21437
rect 43349 21471 43407 21477
rect 43349 21437 43361 21471
rect 43395 21437 43407 21471
rect 43349 21431 43407 21437
rect 31720 21372 33180 21400
rect 37461 21403 37519 21409
rect 31720 21360 31726 21372
rect 37461 21369 37473 21403
rect 37507 21400 37519 21403
rect 38838 21400 38844 21412
rect 37507 21372 38844 21400
rect 37507 21369 37519 21372
rect 37461 21363 37519 21369
rect 38838 21360 38844 21372
rect 38896 21360 38902 21412
rect 41782 21360 41788 21412
rect 41840 21400 41846 21412
rect 43364 21400 43392 21431
rect 41840 21372 43392 21400
rect 43916 21400 43944 21508
rect 47026 21496 47032 21548
rect 47084 21536 47090 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47084 21508 47961 21536
rect 47084 21496 47090 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 43990 21428 43996 21480
rect 44048 21428 44054 21480
rect 48866 21468 48872 21480
rect 44100 21440 48872 21468
rect 44100 21400 44128 21440
rect 48866 21428 48872 21440
rect 48924 21428 48930 21480
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 43916 21372 44128 21400
rect 41840 21360 41846 21372
rect 25188 21304 29776 21332
rect 25188 21292 25194 21304
rect 30190 21292 30196 21344
rect 30248 21292 30254 21344
rect 32585 21335 32643 21341
rect 32585 21301 32597 21335
rect 32631 21332 32643 21335
rect 36446 21332 36452 21344
rect 32631 21304 36452 21332
rect 32631 21301 32643 21304
rect 32585 21295 32643 21301
rect 36446 21292 36452 21304
rect 36504 21292 36510 21344
rect 36538 21292 36544 21344
rect 36596 21292 36602 21344
rect 38657 21335 38715 21341
rect 38657 21301 38669 21335
rect 38703 21332 38715 21335
rect 39206 21332 39212 21344
rect 38703 21304 39212 21332
rect 38703 21301 38715 21304
rect 38657 21295 38715 21301
rect 39206 21292 39212 21304
rect 39264 21292 39270 21344
rect 42794 21292 42800 21344
rect 42852 21292 42858 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 24581 21131 24639 21137
rect 24581 21097 24593 21131
rect 24627 21128 24639 21131
rect 24627 21100 27476 21128
rect 24627 21097 24639 21100
rect 24581 21091 24639 21097
rect 27448 21060 27476 21100
rect 27522 21088 27528 21140
rect 27580 21128 27586 21140
rect 28813 21131 28871 21137
rect 28813 21128 28825 21131
rect 27580 21100 28825 21128
rect 27580 21088 27586 21100
rect 28813 21097 28825 21100
rect 28859 21097 28871 21131
rect 28813 21091 28871 21097
rect 30282 21088 30288 21140
rect 30340 21128 30346 21140
rect 32493 21131 32551 21137
rect 32493 21128 32505 21131
rect 30340 21100 32505 21128
rect 30340 21088 30346 21100
rect 32493 21097 32505 21100
rect 32539 21128 32551 21131
rect 32674 21128 32680 21140
rect 32539 21100 32680 21128
rect 32539 21097 32551 21100
rect 32493 21091 32551 21097
rect 32674 21088 32680 21100
rect 32732 21088 32738 21140
rect 36725 21131 36783 21137
rect 36725 21097 36737 21131
rect 36771 21128 36783 21131
rect 36998 21128 37004 21140
rect 36771 21100 37004 21128
rect 36771 21097 36783 21100
rect 36725 21091 36783 21097
rect 36998 21088 37004 21100
rect 37056 21088 37062 21140
rect 37826 21088 37832 21140
rect 37884 21128 37890 21140
rect 38013 21131 38071 21137
rect 38013 21128 38025 21131
rect 37884 21100 38025 21128
rect 37884 21088 37890 21100
rect 38013 21097 38025 21100
rect 38059 21097 38071 21131
rect 38013 21091 38071 21097
rect 41969 21131 42027 21137
rect 41969 21097 41981 21131
rect 42015 21128 42027 21131
rect 42058 21128 42064 21140
rect 42015 21100 42064 21128
rect 42015 21097 42027 21100
rect 41969 21091 42027 21097
rect 42058 21088 42064 21100
rect 42116 21088 42122 21140
rect 30558 21060 30564 21072
rect 27448 21032 30564 21060
rect 30558 21020 30564 21032
rect 30616 21020 30622 21072
rect 36446 21020 36452 21072
rect 36504 21060 36510 21072
rect 42889 21063 42947 21069
rect 36504 21032 38884 21060
rect 36504 21020 36510 21032
rect 25222 20952 25228 21004
rect 25280 20952 25286 21004
rect 26418 20952 26424 21004
rect 26476 20952 26482 21004
rect 31018 20952 31024 21004
rect 31076 20952 31082 21004
rect 31754 20952 31760 21004
rect 31812 20992 31818 21004
rect 33505 20995 33563 21001
rect 33505 20992 33517 20995
rect 31812 20964 33517 20992
rect 31812 20952 31818 20964
rect 33505 20961 33517 20964
rect 33551 20961 33563 20995
rect 33505 20955 33563 20961
rect 33594 20952 33600 21004
rect 33652 20992 33658 21004
rect 34977 20995 35035 21001
rect 34977 20992 34989 20995
rect 33652 20964 34989 20992
rect 33652 20952 33658 20964
rect 34977 20961 34989 20964
rect 35023 20961 35035 20995
rect 34977 20955 35035 20961
rect 35253 20995 35311 21001
rect 35253 20961 35265 20995
rect 35299 20992 35311 20995
rect 36538 20992 36544 21004
rect 35299 20964 36544 20992
rect 35299 20961 35311 20964
rect 35253 20955 35311 20961
rect 36538 20952 36544 20964
rect 36596 20952 36602 21004
rect 24946 20884 24952 20936
rect 25004 20884 25010 20936
rect 25406 20884 25412 20936
rect 25464 20924 25470 20936
rect 26145 20927 26203 20933
rect 26145 20924 26157 20927
rect 25464 20896 26157 20924
rect 25464 20884 25470 20896
rect 26145 20893 26157 20896
rect 26191 20893 26203 20927
rect 26145 20887 26203 20893
rect 29730 20884 29736 20936
rect 29788 20924 29794 20936
rect 30745 20927 30803 20933
rect 30745 20924 30757 20927
rect 29788 20896 30757 20924
rect 29788 20884 29794 20896
rect 30745 20893 30757 20896
rect 30791 20893 30803 20927
rect 30745 20887 30803 20893
rect 33413 20927 33471 20933
rect 33413 20893 33425 20927
rect 33459 20924 33471 20927
rect 33778 20924 33784 20936
rect 33459 20896 33784 20924
rect 33459 20893 33471 20896
rect 33413 20887 33471 20893
rect 33778 20884 33784 20896
rect 33836 20884 33842 20936
rect 38856 20933 38884 21032
rect 42889 21029 42901 21063
rect 42935 21060 42947 21063
rect 43622 21060 43628 21072
rect 42935 21032 43628 21060
rect 42935 21029 42947 21032
rect 42889 21023 42947 21029
rect 43622 21020 43628 21032
rect 43680 21020 43686 21072
rect 43438 20952 43444 21004
rect 43496 20952 43502 21004
rect 38841 20927 38899 20933
rect 38841 20893 38853 20927
rect 38887 20893 38899 20927
rect 38841 20887 38899 20893
rect 40034 20884 40040 20936
rect 40092 20924 40098 20936
rect 40221 20927 40279 20933
rect 40221 20924 40233 20927
rect 40092 20896 40233 20924
rect 40092 20884 40098 20896
rect 40221 20893 40233 20896
rect 40267 20893 40279 20927
rect 40221 20887 40279 20893
rect 41598 20884 41604 20936
rect 41656 20884 41662 20936
rect 43257 20927 43315 20933
rect 43257 20893 43269 20927
rect 43303 20924 43315 20927
rect 44269 20927 44327 20933
rect 44269 20924 44281 20927
rect 43303 20896 44281 20924
rect 43303 20893 43315 20896
rect 43257 20887 43315 20893
rect 44269 20893 44281 20896
rect 44315 20893 44327 20927
rect 44269 20887 44327 20893
rect 26878 20816 26884 20868
rect 26936 20816 26942 20868
rect 27706 20816 27712 20868
rect 27764 20856 27770 20868
rect 28169 20859 28227 20865
rect 28169 20856 28181 20859
rect 27764 20828 28181 20856
rect 27764 20816 27770 20828
rect 28169 20825 28181 20828
rect 28215 20825 28227 20859
rect 28169 20819 28227 20825
rect 30926 20816 30932 20868
rect 30984 20856 30990 20868
rect 33321 20859 33379 20865
rect 33321 20856 33333 20859
rect 30984 20828 31510 20856
rect 32416 20828 33333 20856
rect 30984 20816 30990 20828
rect 25038 20748 25044 20800
rect 25096 20748 25102 20800
rect 29270 20748 29276 20800
rect 29328 20788 29334 20800
rect 32416 20788 32444 20828
rect 33321 20825 33333 20828
rect 33367 20825 33379 20859
rect 33321 20819 33379 20825
rect 35342 20816 35348 20868
rect 35400 20856 35406 20868
rect 35400 20828 35742 20856
rect 35400 20816 35406 20828
rect 37090 20816 37096 20868
rect 37148 20856 37154 20868
rect 38746 20856 38752 20868
rect 37148 20828 38752 20856
rect 37148 20816 37154 20828
rect 38746 20816 38752 20828
rect 38804 20816 38810 20868
rect 40494 20816 40500 20868
rect 40552 20816 40558 20868
rect 43349 20859 43407 20865
rect 42812 20828 43024 20856
rect 29328 20760 32444 20788
rect 32953 20791 33011 20797
rect 29328 20748 29334 20760
rect 32953 20757 32965 20791
rect 32999 20788 33011 20791
rect 34422 20788 34428 20800
rect 32999 20760 34428 20788
rect 32999 20757 33011 20760
rect 32953 20751 33011 20757
rect 34422 20748 34428 20760
rect 34480 20748 34486 20800
rect 38657 20791 38715 20797
rect 38657 20757 38669 20791
rect 38703 20788 38715 20791
rect 42812 20788 42840 20828
rect 38703 20760 42840 20788
rect 42996 20788 43024 20828
rect 43349 20825 43361 20859
rect 43395 20856 43407 20859
rect 44082 20856 44088 20868
rect 43395 20828 44088 20856
rect 43395 20825 43407 20828
rect 43349 20819 43407 20825
rect 44082 20816 44088 20828
rect 44140 20816 44146 20868
rect 43898 20788 43904 20800
rect 42996 20760 43904 20788
rect 38703 20757 38715 20760
rect 38657 20751 38715 20757
rect 43898 20748 43904 20760
rect 43956 20748 43962 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 28718 20544 28724 20596
rect 28776 20584 28782 20596
rect 28905 20587 28963 20593
rect 28905 20584 28917 20587
rect 28776 20556 28917 20584
rect 28776 20544 28782 20556
rect 28905 20553 28917 20556
rect 28951 20553 28963 20587
rect 28905 20547 28963 20553
rect 31754 20544 31760 20596
rect 31812 20544 31818 20596
rect 36173 20587 36231 20593
rect 36173 20553 36185 20587
rect 36219 20553 36231 20587
rect 36173 20547 36231 20553
rect 27522 20516 27528 20528
rect 26896 20488 27528 20516
rect 26896 20460 26924 20488
rect 27522 20476 27528 20488
rect 27580 20516 27586 20528
rect 27580 20488 27922 20516
rect 27580 20476 27586 20488
rect 29638 20476 29644 20528
rect 29696 20516 29702 20528
rect 30282 20516 30288 20528
rect 29696 20488 30288 20516
rect 29696 20476 29702 20488
rect 30282 20476 30288 20488
rect 30340 20476 30346 20528
rect 30926 20476 30932 20528
rect 30984 20476 30990 20528
rect 34514 20516 34520 20528
rect 33980 20488 34520 20516
rect 25314 20448 25320 20460
rect 25162 20420 25320 20448
rect 25314 20408 25320 20420
rect 25372 20448 25378 20460
rect 26878 20448 26884 20460
rect 25372 20420 26884 20448
rect 25372 20408 25378 20420
rect 26878 20408 26884 20420
rect 26936 20408 26942 20460
rect 33980 20457 34008 20488
rect 34514 20476 34520 20488
rect 34572 20476 34578 20528
rect 36188 20516 36216 20547
rect 36630 20544 36636 20596
rect 36688 20544 36694 20596
rect 44361 20587 44419 20593
rect 44361 20553 44373 20587
rect 44407 20584 44419 20587
rect 45186 20584 45192 20596
rect 44407 20556 45192 20584
rect 44407 20553 44419 20556
rect 44361 20547 44419 20553
rect 45186 20544 45192 20556
rect 45244 20544 45250 20596
rect 38654 20516 38660 20528
rect 36188 20488 38660 20516
rect 38654 20476 38660 20488
rect 38712 20476 38718 20528
rect 41598 20516 41604 20528
rect 39882 20488 41604 20516
rect 41598 20476 41604 20488
rect 41656 20476 41662 20528
rect 43073 20519 43131 20525
rect 43073 20485 43085 20519
rect 43119 20516 43131 20519
rect 47026 20516 47032 20528
rect 43119 20488 47032 20516
rect 43119 20485 43131 20488
rect 43073 20479 43131 20485
rect 47026 20476 47032 20488
rect 47084 20476 47090 20528
rect 33965 20451 34023 20457
rect 33965 20417 33977 20451
rect 34011 20417 34023 20451
rect 33965 20411 34023 20417
rect 35342 20408 35348 20460
rect 35400 20408 35406 20460
rect 35986 20408 35992 20460
rect 36044 20448 36050 20460
rect 36541 20451 36599 20457
rect 36541 20448 36553 20451
rect 36044 20420 36553 20448
rect 36044 20408 36050 20420
rect 36541 20417 36553 20420
rect 36587 20417 36599 20451
rect 36541 20411 36599 20417
rect 39942 20408 39948 20460
rect 40000 20448 40006 20460
rect 42889 20451 42947 20457
rect 42889 20448 42901 20451
rect 40000 20420 42901 20448
rect 40000 20408 40006 20420
rect 42889 20417 42901 20420
rect 42935 20417 42947 20451
rect 42889 20411 42947 20417
rect 44269 20451 44327 20457
rect 44269 20417 44281 20451
rect 44315 20448 44327 20451
rect 45281 20451 45339 20457
rect 45281 20448 45293 20451
rect 44315 20420 45293 20448
rect 44315 20417 44327 20420
rect 44269 20411 44327 20417
rect 45281 20417 45293 20420
rect 45327 20417 45339 20451
rect 45281 20411 45339 20417
rect 46934 20408 46940 20460
rect 46992 20448 46998 20460
rect 47949 20451 48007 20457
rect 47949 20448 47961 20451
rect 46992 20420 47961 20448
rect 46992 20408 46998 20420
rect 47949 20417 47961 20420
rect 47995 20417 48007 20451
rect 47949 20411 48007 20417
rect 23750 20340 23756 20392
rect 23808 20340 23814 20392
rect 24026 20340 24032 20392
rect 24084 20340 24090 20392
rect 25406 20340 25412 20392
rect 25464 20380 25470 20392
rect 27157 20383 27215 20389
rect 27157 20380 27169 20383
rect 25464 20352 27169 20380
rect 25464 20340 25470 20352
rect 27157 20349 27169 20352
rect 27203 20349 27215 20383
rect 27433 20383 27491 20389
rect 27433 20380 27445 20383
rect 27157 20343 27215 20349
rect 27264 20352 27445 20380
rect 26602 20272 26608 20324
rect 26660 20312 26666 20324
rect 27264 20312 27292 20352
rect 27433 20349 27445 20352
rect 27479 20349 27491 20383
rect 27433 20343 27491 20349
rect 29730 20340 29736 20392
rect 29788 20380 29794 20392
rect 30009 20383 30067 20389
rect 30009 20380 30021 20383
rect 29788 20352 30021 20380
rect 29788 20340 29794 20352
rect 30009 20349 30021 20352
rect 30055 20349 30067 20383
rect 30009 20343 30067 20349
rect 34241 20383 34299 20389
rect 34241 20349 34253 20383
rect 34287 20380 34299 20383
rect 34698 20380 34704 20392
rect 34287 20352 34704 20380
rect 34287 20349 34299 20352
rect 34241 20343 34299 20349
rect 34698 20340 34704 20352
rect 34756 20340 34762 20392
rect 36630 20340 36636 20392
rect 36688 20380 36694 20392
rect 36725 20383 36783 20389
rect 36725 20380 36737 20383
rect 36688 20352 36737 20380
rect 36688 20340 36694 20352
rect 36725 20349 36737 20352
rect 36771 20349 36783 20383
rect 36725 20343 36783 20349
rect 38381 20383 38439 20389
rect 38381 20349 38393 20383
rect 38427 20349 38439 20383
rect 38381 20343 38439 20349
rect 38657 20383 38715 20389
rect 38657 20349 38669 20383
rect 38703 20380 38715 20383
rect 38746 20380 38752 20392
rect 38703 20352 38752 20380
rect 38703 20349 38715 20352
rect 38657 20343 38715 20349
rect 26660 20284 27292 20312
rect 26660 20272 26666 20284
rect 25501 20247 25559 20253
rect 25501 20213 25513 20247
rect 25547 20244 25559 20247
rect 26234 20244 26240 20256
rect 25547 20216 26240 20244
rect 25547 20213 25559 20216
rect 25501 20207 25559 20213
rect 26234 20204 26240 20216
rect 26292 20204 26298 20256
rect 35434 20204 35440 20256
rect 35492 20244 35498 20256
rect 35713 20247 35771 20253
rect 35713 20244 35725 20247
rect 35492 20216 35725 20244
rect 35492 20204 35498 20216
rect 35713 20213 35725 20216
rect 35759 20213 35771 20247
rect 38396 20244 38424 20343
rect 38746 20340 38752 20352
rect 38804 20340 38810 20392
rect 44542 20340 44548 20392
rect 44600 20340 44606 20392
rect 49142 20340 49148 20392
rect 49200 20340 49206 20392
rect 40034 20244 40040 20256
rect 38396 20216 40040 20244
rect 35713 20207 35771 20213
rect 40034 20204 40040 20216
rect 40092 20204 40098 20256
rect 40126 20204 40132 20256
rect 40184 20204 40190 20256
rect 42150 20204 42156 20256
rect 42208 20244 42214 20256
rect 43901 20247 43959 20253
rect 43901 20244 43913 20247
rect 42208 20216 43913 20244
rect 42208 20204 42214 20216
rect 43901 20213 43913 20216
rect 43947 20213 43959 20247
rect 43901 20207 43959 20213
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 29178 20000 29184 20052
rect 29236 20000 29242 20052
rect 32848 20043 32906 20049
rect 32848 20009 32860 20043
rect 32894 20040 32906 20043
rect 34790 20040 34796 20052
rect 32894 20012 34796 20040
rect 32894 20009 32906 20012
rect 32848 20003 32906 20009
rect 34790 20000 34796 20012
rect 34848 20000 34854 20052
rect 34885 20043 34943 20049
rect 34885 20009 34897 20043
rect 34931 20040 34943 20043
rect 39942 20040 39948 20052
rect 34931 20012 39948 20040
rect 34931 20009 34943 20012
rect 34885 20003 34943 20009
rect 39942 20000 39948 20012
rect 40000 20000 40006 20052
rect 40126 20000 40132 20052
rect 40184 20040 40190 20052
rect 40294 20043 40352 20049
rect 40294 20040 40306 20043
rect 40184 20012 40306 20040
rect 40184 20000 40190 20012
rect 40294 20009 40306 20012
rect 40340 20009 40352 20043
rect 40294 20003 40352 20009
rect 41782 20000 41788 20052
rect 41840 20000 41846 20052
rect 42508 20043 42566 20049
rect 42508 20009 42520 20043
rect 42554 20040 42566 20043
rect 44358 20040 44364 20052
rect 42554 20012 44364 20040
rect 42554 20009 42566 20012
rect 42508 20003 42566 20009
rect 44358 20000 44364 20012
rect 44416 20000 44422 20052
rect 40144 19972 40172 20000
rect 39132 19944 40172 19972
rect 23750 19864 23756 19916
rect 23808 19904 23814 19916
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 23808 19876 24593 19904
rect 23808 19864 23814 19876
rect 24581 19873 24593 19876
rect 24627 19904 24639 19907
rect 25406 19904 25412 19916
rect 24627 19876 25412 19904
rect 24627 19873 24639 19876
rect 24581 19867 24639 19873
rect 25406 19864 25412 19876
rect 25464 19904 25470 19916
rect 27433 19907 27491 19913
rect 27433 19904 27445 19907
rect 25464 19876 27445 19904
rect 25464 19864 25470 19876
rect 27433 19873 27445 19876
rect 27479 19904 27491 19907
rect 27798 19904 27804 19916
rect 27479 19876 27804 19904
rect 27479 19873 27491 19876
rect 27433 19867 27491 19873
rect 27798 19864 27804 19876
rect 27856 19864 27862 19916
rect 28902 19864 28908 19916
rect 28960 19904 28966 19916
rect 39132 19913 39160 19944
rect 39117 19907 39175 19913
rect 28960 19876 36676 19904
rect 28960 19864 28966 19876
rect 32582 19796 32588 19848
rect 32640 19796 32646 19848
rect 35066 19796 35072 19848
rect 35124 19796 35130 19848
rect 36648 19845 36676 19876
rect 39117 19873 39129 19907
rect 39163 19873 39175 19907
rect 39117 19867 39175 19873
rect 40034 19864 40040 19916
rect 40092 19904 40098 19916
rect 41322 19904 41328 19916
rect 40092 19876 41328 19904
rect 40092 19864 40098 19876
rect 41322 19864 41328 19876
rect 41380 19864 41386 19916
rect 42245 19907 42303 19913
rect 42245 19873 42257 19907
rect 42291 19904 42303 19907
rect 43990 19904 43996 19916
rect 42291 19876 43996 19904
rect 42291 19873 42303 19876
rect 42245 19867 42303 19873
rect 43990 19864 43996 19876
rect 44048 19864 44054 19916
rect 36633 19839 36691 19845
rect 36633 19805 36645 19839
rect 36679 19805 36691 19839
rect 36633 19799 36691 19805
rect 38838 19796 38844 19848
rect 38896 19796 38902 19848
rect 38933 19839 38991 19845
rect 38933 19805 38945 19839
rect 38979 19836 38991 19839
rect 39666 19836 39672 19848
rect 38979 19808 39672 19836
rect 38979 19805 38991 19808
rect 38933 19799 38991 19805
rect 39666 19796 39672 19808
rect 39724 19796 39730 19848
rect 41598 19836 41604 19848
rect 41446 19808 41604 19836
rect 41598 19796 41604 19808
rect 41656 19836 41662 19848
rect 41656 19808 42288 19836
rect 41656 19796 41662 19808
rect 24857 19771 24915 19777
rect 24857 19737 24869 19771
rect 24903 19737 24915 19771
rect 24857 19731 24915 19737
rect 24872 19700 24900 19731
rect 25314 19728 25320 19780
rect 25372 19728 25378 19780
rect 27614 19728 27620 19780
rect 27672 19768 27678 19780
rect 27709 19771 27767 19777
rect 27709 19768 27721 19771
rect 27672 19740 27721 19768
rect 27672 19728 27678 19740
rect 27709 19737 27721 19740
rect 27755 19737 27767 19771
rect 34146 19768 34152 19780
rect 27709 19731 27767 19737
rect 28092 19740 28198 19768
rect 34086 19740 34152 19768
rect 26234 19700 26240 19712
rect 24872 19672 26240 19700
rect 26234 19660 26240 19672
rect 26292 19660 26298 19712
rect 26329 19703 26387 19709
rect 26329 19669 26341 19703
rect 26375 19700 26387 19703
rect 26602 19700 26608 19712
rect 26375 19672 26608 19700
rect 26375 19669 26387 19672
rect 26329 19663 26387 19669
rect 26602 19660 26608 19672
rect 26660 19660 26666 19712
rect 27522 19660 27528 19712
rect 27580 19700 27586 19712
rect 28092 19700 28120 19740
rect 34146 19728 34152 19740
rect 34204 19768 34210 19780
rect 35342 19768 35348 19780
rect 34204 19740 35348 19768
rect 34204 19728 34210 19740
rect 35342 19728 35348 19740
rect 35400 19768 35406 19780
rect 36170 19768 36176 19780
rect 35400 19740 36176 19768
rect 35400 19728 35406 19740
rect 36170 19728 36176 19740
rect 36228 19728 36234 19780
rect 40586 19768 40592 19780
rect 36464 19740 40592 19768
rect 27580 19672 28120 19700
rect 34333 19703 34391 19709
rect 27580 19660 27586 19672
rect 34333 19669 34345 19703
rect 34379 19700 34391 19703
rect 34698 19700 34704 19712
rect 34379 19672 34704 19700
rect 34379 19669 34391 19672
rect 34333 19663 34391 19669
rect 34698 19660 34704 19672
rect 34756 19700 34762 19712
rect 35618 19700 35624 19712
rect 34756 19672 35624 19700
rect 34756 19660 34762 19672
rect 35618 19660 35624 19672
rect 35676 19660 35682 19712
rect 36464 19709 36492 19740
rect 40586 19728 40592 19740
rect 40644 19728 40650 19780
rect 42260 19768 42288 19808
rect 43898 19796 43904 19848
rect 43956 19836 43962 19848
rect 45373 19839 45431 19845
rect 45373 19836 45385 19839
rect 43956 19808 45385 19836
rect 43956 19796 43962 19808
rect 45373 19805 45385 19808
rect 45419 19805 45431 19839
rect 45373 19799 45431 19805
rect 47949 19839 48007 19845
rect 47949 19805 47961 19839
rect 47995 19805 48007 19839
rect 47949 19799 48007 19805
rect 42978 19768 42984 19780
rect 41708 19740 41920 19768
rect 42260 19740 42984 19768
rect 36449 19703 36507 19709
rect 36449 19669 36461 19703
rect 36495 19669 36507 19703
rect 36449 19663 36507 19669
rect 36538 19660 36544 19712
rect 36596 19700 36602 19712
rect 38473 19703 38531 19709
rect 38473 19700 38485 19703
rect 36596 19672 38485 19700
rect 36596 19660 36602 19672
rect 38473 19669 38485 19672
rect 38519 19669 38531 19703
rect 38473 19663 38531 19669
rect 40494 19660 40500 19712
rect 40552 19700 40558 19712
rect 41046 19700 41052 19712
rect 40552 19672 41052 19700
rect 40552 19660 40558 19672
rect 41046 19660 41052 19672
rect 41104 19700 41110 19712
rect 41708 19700 41736 19740
rect 41104 19672 41736 19700
rect 41892 19700 41920 19740
rect 42978 19728 42984 19740
rect 43036 19728 43042 19780
rect 43993 19703 44051 19709
rect 43993 19700 44005 19703
rect 41892 19672 44005 19700
rect 41104 19660 41110 19672
rect 43993 19669 44005 19672
rect 44039 19669 44051 19703
rect 43993 19663 44051 19669
rect 45189 19703 45247 19709
rect 45189 19669 45201 19703
rect 45235 19700 45247 19703
rect 47964 19700 47992 19799
rect 49142 19728 49148 19780
rect 49200 19728 49206 19780
rect 45235 19672 47992 19700
rect 45235 19669 45247 19672
rect 45189 19663 45247 19669
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 23382 19456 23388 19508
rect 23440 19496 23446 19508
rect 23569 19499 23627 19505
rect 23569 19496 23581 19499
rect 23440 19468 23581 19496
rect 23440 19456 23446 19468
rect 23569 19465 23581 19468
rect 23615 19465 23627 19499
rect 23569 19459 23627 19465
rect 28813 19499 28871 19505
rect 28813 19465 28825 19499
rect 28859 19496 28871 19499
rect 28902 19496 28908 19508
rect 28859 19468 28908 19496
rect 28859 19465 28871 19468
rect 28813 19459 28871 19465
rect 28902 19456 28908 19468
rect 28960 19456 28966 19508
rect 29273 19499 29331 19505
rect 29273 19465 29285 19499
rect 29319 19496 29331 19499
rect 30098 19496 30104 19508
rect 29319 19468 30104 19496
rect 29319 19465 29331 19468
rect 29273 19459 29331 19465
rect 30098 19456 30104 19468
rect 30156 19456 30162 19508
rect 33502 19456 33508 19508
rect 33560 19496 33566 19508
rect 33873 19499 33931 19505
rect 33873 19496 33885 19499
rect 33560 19468 33885 19496
rect 33560 19456 33566 19468
rect 33873 19465 33885 19468
rect 33919 19496 33931 19499
rect 35069 19499 35127 19505
rect 35069 19496 35081 19499
rect 33919 19468 35081 19496
rect 33919 19465 33931 19468
rect 33873 19459 33931 19465
rect 35069 19465 35081 19468
rect 35115 19465 35127 19499
rect 35069 19459 35127 19465
rect 35158 19456 35164 19508
rect 35216 19456 35222 19508
rect 38841 19499 38899 19505
rect 38841 19465 38853 19499
rect 38887 19496 38899 19499
rect 44913 19499 44971 19505
rect 38887 19468 43576 19496
rect 38887 19465 38899 19468
rect 38841 19459 38899 19465
rect 27798 19388 27804 19440
rect 27856 19428 27862 19440
rect 28077 19431 28135 19437
rect 28077 19428 28089 19431
rect 27856 19400 28089 19428
rect 27856 19388 27862 19400
rect 28077 19397 28089 19400
rect 28123 19397 28135 19431
rect 28077 19391 28135 19397
rect 30926 19388 30932 19440
rect 30984 19388 30990 19440
rect 32490 19388 32496 19440
rect 32548 19388 32554 19440
rect 33962 19388 33968 19440
rect 34020 19428 34026 19440
rect 34330 19428 34336 19440
rect 34020 19400 34336 19428
rect 34020 19388 34026 19400
rect 34330 19388 34336 19400
rect 34388 19388 34394 19440
rect 23290 19320 23296 19372
rect 23348 19360 23354 19372
rect 23937 19363 23995 19369
rect 23937 19360 23949 19363
rect 23348 19332 23949 19360
rect 23348 19320 23354 19332
rect 23937 19329 23949 19332
rect 23983 19329 23995 19363
rect 23937 19323 23995 19329
rect 24029 19363 24087 19369
rect 24029 19329 24041 19363
rect 24075 19360 24087 19363
rect 25314 19360 25320 19372
rect 24075 19332 25320 19360
rect 24075 19329 24087 19332
rect 24029 19323 24087 19329
rect 25314 19320 25320 19332
rect 25372 19320 25378 19372
rect 27341 19363 27399 19369
rect 27341 19329 27353 19363
rect 27387 19360 27399 19363
rect 27430 19360 27436 19372
rect 27387 19332 27436 19360
rect 27387 19329 27399 19332
rect 27341 19323 27399 19329
rect 27430 19320 27436 19332
rect 27488 19320 27494 19372
rect 28810 19320 28816 19372
rect 28868 19360 28874 19372
rect 29181 19363 29239 19369
rect 29181 19360 29193 19363
rect 28868 19332 29193 19360
rect 28868 19320 28874 19332
rect 29181 19329 29193 19332
rect 29227 19329 29239 19363
rect 29181 19323 29239 19329
rect 32766 19320 32772 19372
rect 32824 19360 32830 19372
rect 32824 19332 34376 19360
rect 32824 19320 32830 19332
rect 24118 19252 24124 19304
rect 24176 19252 24182 19304
rect 29365 19295 29423 19301
rect 29365 19261 29377 19295
rect 29411 19261 29423 19295
rect 29365 19255 29423 19261
rect 28718 19184 28724 19236
rect 28776 19224 28782 19236
rect 29380 19224 29408 19255
rect 29730 19252 29736 19304
rect 29788 19292 29794 19304
rect 30009 19295 30067 19301
rect 30009 19292 30021 19295
rect 29788 19264 30021 19292
rect 29788 19252 29794 19264
rect 30009 19261 30021 19264
rect 30055 19261 30067 19295
rect 30009 19255 30067 19261
rect 30285 19295 30343 19301
rect 30285 19261 30297 19295
rect 30331 19292 30343 19295
rect 31754 19292 31760 19304
rect 30331 19264 31760 19292
rect 30331 19261 30343 19264
rect 30285 19255 30343 19261
rect 31754 19252 31760 19264
rect 31812 19252 31818 19304
rect 34057 19295 34115 19301
rect 34057 19261 34069 19295
rect 34103 19261 34115 19295
rect 34348 19292 34376 19332
rect 34422 19320 34428 19372
rect 34480 19360 34486 19372
rect 39025 19363 39083 19369
rect 39025 19360 39037 19363
rect 34480 19332 39037 19360
rect 34480 19320 34486 19332
rect 39025 19329 39037 19332
rect 39071 19329 39083 19363
rect 39025 19323 39083 19329
rect 42981 19363 43039 19369
rect 42981 19329 42993 19363
rect 43027 19329 43039 19363
rect 42981 19323 43039 19329
rect 43073 19363 43131 19369
rect 43073 19329 43085 19363
rect 43119 19360 43131 19363
rect 43346 19360 43352 19372
rect 43119 19332 43352 19360
rect 43119 19329 43131 19332
rect 43073 19323 43131 19329
rect 34348 19264 34744 19292
rect 34057 19255 34115 19261
rect 28776 19196 29408 19224
rect 28776 19184 28782 19196
rect 32214 19184 32220 19236
rect 32272 19224 32278 19236
rect 33505 19227 33563 19233
rect 33505 19224 33517 19227
rect 32272 19196 33517 19224
rect 32272 19184 32278 19196
rect 33505 19193 33517 19196
rect 33551 19193 33563 19227
rect 33505 19187 33563 19193
rect 33870 19184 33876 19236
rect 33928 19224 33934 19236
rect 34072 19224 34100 19255
rect 34716 19233 34744 19264
rect 35342 19252 35348 19304
rect 35400 19252 35406 19304
rect 42061 19295 42119 19301
rect 42061 19261 42073 19295
rect 42107 19292 42119 19295
rect 42996 19292 43024 19323
rect 43346 19320 43352 19332
rect 43404 19320 43410 19372
rect 43548 19360 43576 19468
rect 44913 19465 44925 19499
rect 44959 19496 44971 19499
rect 47946 19496 47952 19508
rect 44959 19468 47952 19496
rect 44959 19465 44971 19468
rect 44913 19459 44971 19465
rect 47946 19456 47952 19468
rect 48004 19456 48010 19508
rect 43898 19388 43904 19440
rect 43956 19388 43962 19440
rect 45097 19363 45155 19369
rect 45097 19360 45109 19363
rect 43548 19332 45109 19360
rect 45097 19329 45109 19332
rect 45143 19329 45155 19363
rect 45097 19323 45155 19329
rect 42107 19264 43024 19292
rect 43257 19295 43315 19301
rect 42107 19261 42119 19264
rect 42061 19255 42119 19261
rect 43257 19261 43269 19295
rect 43303 19292 43315 19295
rect 43806 19292 43812 19304
rect 43303 19264 43812 19292
rect 43303 19261 43315 19264
rect 43257 19255 43315 19261
rect 43806 19252 43812 19264
rect 43864 19252 43870 19304
rect 44085 19295 44143 19301
rect 44085 19261 44097 19295
rect 44131 19292 44143 19295
rect 46934 19292 46940 19304
rect 44131 19264 46940 19292
rect 44131 19261 44143 19264
rect 44085 19255 44143 19261
rect 46934 19252 46940 19264
rect 46992 19252 46998 19304
rect 33928 19196 34100 19224
rect 34701 19227 34759 19233
rect 33928 19184 33934 19196
rect 34701 19193 34713 19227
rect 34747 19193 34759 19227
rect 34701 19187 34759 19193
rect 42978 19184 42984 19236
rect 43036 19224 43042 19236
rect 43990 19224 43996 19236
rect 43036 19196 43996 19224
rect 43036 19184 43042 19196
rect 43990 19184 43996 19196
rect 44048 19184 44054 19236
rect 30374 19116 30380 19168
rect 30432 19156 30438 19168
rect 31757 19159 31815 19165
rect 31757 19156 31769 19159
rect 30432 19128 31769 19156
rect 30432 19116 30438 19128
rect 31757 19125 31769 19128
rect 31803 19125 31815 19159
rect 31757 19119 31815 19125
rect 32122 19116 32128 19168
rect 32180 19156 32186 19168
rect 32585 19159 32643 19165
rect 32585 19156 32597 19159
rect 32180 19128 32597 19156
rect 32180 19116 32186 19128
rect 32585 19125 32597 19128
rect 32631 19125 32643 19159
rect 32585 19119 32643 19125
rect 32858 19116 32864 19168
rect 32916 19156 32922 19168
rect 36998 19156 37004 19168
rect 32916 19128 37004 19156
rect 32916 19116 32922 19128
rect 36998 19116 37004 19128
rect 37056 19116 37062 19168
rect 42334 19116 42340 19168
rect 42392 19156 42398 19168
rect 42613 19159 42671 19165
rect 42613 19156 42625 19159
rect 42392 19128 42625 19156
rect 42392 19116 42398 19128
rect 42613 19125 42625 19128
rect 42659 19125 42671 19159
rect 42613 19119 42671 19125
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 22462 18912 22468 18964
rect 22520 18952 22526 18964
rect 24581 18955 24639 18961
rect 24581 18952 24593 18955
rect 22520 18924 24593 18952
rect 22520 18912 22526 18924
rect 24581 18921 24593 18924
rect 24627 18921 24639 18955
rect 24581 18915 24639 18921
rect 27157 18955 27215 18961
rect 27157 18921 27169 18955
rect 27203 18952 27215 18955
rect 35066 18952 35072 18964
rect 27203 18924 35072 18952
rect 27203 18921 27215 18924
rect 27157 18915 27215 18921
rect 35066 18912 35072 18924
rect 35124 18912 35130 18964
rect 35618 18952 35624 18964
rect 35452 18924 35624 18952
rect 29362 18844 29368 18896
rect 29420 18884 29426 18896
rect 32122 18884 32128 18896
rect 29420 18856 32128 18884
rect 29420 18844 29426 18856
rect 32122 18844 32128 18856
rect 32180 18844 32186 18896
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18816 25283 18819
rect 25498 18816 25504 18828
rect 25271 18788 25504 18816
rect 25271 18785 25283 18788
rect 25225 18779 25283 18785
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 26234 18776 26240 18828
rect 26292 18816 26298 18828
rect 27709 18819 27767 18825
rect 27709 18816 27721 18819
rect 26292 18788 27721 18816
rect 26292 18776 26298 18788
rect 27709 18785 27721 18788
rect 27755 18785 27767 18819
rect 27709 18779 27767 18785
rect 29730 18776 29736 18828
rect 29788 18816 29794 18828
rect 30653 18819 30711 18825
rect 30653 18816 30665 18819
rect 29788 18788 30665 18816
rect 29788 18776 29794 18788
rect 30653 18785 30665 18788
rect 30699 18816 30711 18819
rect 32582 18816 32588 18828
rect 30699 18788 32588 18816
rect 30699 18785 30711 18788
rect 30653 18779 30711 18785
rect 32582 18776 32588 18788
rect 32640 18776 32646 18828
rect 32858 18776 32864 18828
rect 32916 18776 32922 18828
rect 35250 18776 35256 18828
rect 35308 18816 35314 18828
rect 35452 18825 35480 18924
rect 35618 18912 35624 18924
rect 35676 18912 35682 18964
rect 41782 18912 41788 18964
rect 41840 18912 41846 18964
rect 36725 18887 36783 18893
rect 36725 18884 36737 18887
rect 35544 18856 36737 18884
rect 35345 18819 35403 18825
rect 35345 18816 35357 18819
rect 35308 18788 35357 18816
rect 35308 18776 35314 18788
rect 35345 18785 35357 18788
rect 35391 18785 35403 18819
rect 35345 18779 35403 18785
rect 35437 18819 35495 18825
rect 35437 18785 35449 18819
rect 35483 18785 35495 18819
rect 35437 18779 35495 18785
rect 27246 18708 27252 18760
rect 27304 18748 27310 18760
rect 27617 18751 27675 18757
rect 27617 18748 27629 18751
rect 27304 18720 27629 18748
rect 27304 18708 27310 18720
rect 27617 18717 27629 18720
rect 27663 18717 27675 18751
rect 27617 18711 27675 18717
rect 28718 18708 28724 18760
rect 28776 18708 28782 18760
rect 31662 18708 31668 18760
rect 31720 18748 31726 18760
rect 31720 18720 32536 18748
rect 31720 18708 31726 18720
rect 27430 18640 27436 18692
rect 27488 18680 27494 18692
rect 29917 18683 29975 18689
rect 29917 18680 29929 18683
rect 27488 18652 29929 18680
rect 27488 18640 27494 18652
rect 29917 18649 29929 18652
rect 29963 18680 29975 18683
rect 32398 18680 32404 18692
rect 29963 18652 32404 18680
rect 29963 18649 29975 18652
rect 29917 18643 29975 18649
rect 32398 18640 32404 18652
rect 32456 18640 32462 18692
rect 32508 18680 32536 18720
rect 34422 18708 34428 18760
rect 34480 18748 34486 18760
rect 35544 18748 35572 18856
rect 36725 18853 36737 18856
rect 36771 18853 36783 18887
rect 36725 18847 36783 18853
rect 37642 18816 37648 18828
rect 36280 18788 37648 18816
rect 36280 18757 36308 18788
rect 37642 18776 37648 18788
rect 37700 18776 37706 18828
rect 40862 18776 40868 18828
rect 40920 18816 40926 18828
rect 40957 18819 41015 18825
rect 40957 18816 40969 18819
rect 40920 18788 40969 18816
rect 40920 18776 40926 18788
rect 40957 18785 40969 18788
rect 41003 18785 41015 18819
rect 40957 18779 41015 18785
rect 41046 18776 41052 18828
rect 41104 18776 41110 18828
rect 41414 18776 41420 18828
rect 41472 18816 41478 18828
rect 41693 18819 41751 18825
rect 41693 18816 41705 18819
rect 41472 18788 41705 18816
rect 41472 18776 41478 18788
rect 41693 18785 41705 18788
rect 41739 18785 41751 18819
rect 41800 18816 41828 18912
rect 41969 18819 42027 18825
rect 41969 18816 41981 18819
rect 41800 18788 41981 18816
rect 41693 18779 41751 18785
rect 41969 18785 41981 18788
rect 42015 18785 42027 18819
rect 41969 18779 42027 18785
rect 34480 18720 35572 18748
rect 36265 18751 36323 18757
rect 34480 18708 34486 18720
rect 36265 18717 36277 18751
rect 36311 18717 36323 18751
rect 36265 18711 36323 18717
rect 36909 18751 36967 18757
rect 36909 18717 36921 18751
rect 36955 18748 36967 18751
rect 38286 18748 38292 18760
rect 36955 18720 38292 18748
rect 36955 18717 36967 18720
rect 36909 18711 36967 18717
rect 38286 18708 38292 18720
rect 38344 18708 38350 18760
rect 47946 18708 47952 18760
rect 48004 18708 48010 18760
rect 49142 18708 49148 18760
rect 49200 18708 49206 18760
rect 32858 18680 32864 18692
rect 32508 18652 32864 18680
rect 32858 18640 32864 18652
rect 32916 18640 32922 18692
rect 34146 18680 34152 18692
rect 34086 18652 34152 18680
rect 34146 18640 34152 18652
rect 34204 18640 34210 18692
rect 40402 18680 40408 18692
rect 34900 18652 40408 18680
rect 24946 18572 24952 18624
rect 25004 18572 25010 18624
rect 25041 18615 25099 18621
rect 25041 18581 25053 18615
rect 25087 18612 25099 18615
rect 26326 18612 26332 18624
rect 25087 18584 26332 18612
rect 25087 18581 25099 18584
rect 25041 18575 25099 18581
rect 26326 18572 26332 18584
rect 26384 18572 26390 18624
rect 26418 18572 26424 18624
rect 26476 18612 26482 18624
rect 27525 18615 27583 18621
rect 27525 18612 27537 18615
rect 26476 18584 27537 18612
rect 26476 18572 26482 18584
rect 27525 18581 27537 18584
rect 27571 18581 27583 18615
rect 27525 18575 27583 18581
rect 34330 18572 34336 18624
rect 34388 18572 34394 18624
rect 34900 18621 34928 18652
rect 40402 18640 40408 18652
rect 40460 18640 40466 18692
rect 43990 18680 43996 18692
rect 43194 18652 43996 18680
rect 43990 18640 43996 18652
rect 44048 18640 44054 18692
rect 34885 18615 34943 18621
rect 34885 18581 34897 18615
rect 34931 18581 34943 18615
rect 34885 18575 34943 18581
rect 35250 18572 35256 18624
rect 35308 18572 35314 18624
rect 35710 18572 35716 18624
rect 35768 18612 35774 18624
rect 36081 18615 36139 18621
rect 36081 18612 36093 18615
rect 35768 18584 36093 18612
rect 35768 18572 35774 18584
rect 36081 18581 36093 18584
rect 36127 18581 36139 18615
rect 36081 18575 36139 18581
rect 39482 18572 39488 18624
rect 39540 18612 39546 18624
rect 40497 18615 40555 18621
rect 40497 18612 40509 18615
rect 39540 18584 40509 18612
rect 39540 18572 39546 18584
rect 40497 18581 40509 18584
rect 40543 18581 40555 18615
rect 40497 18575 40555 18581
rect 40862 18572 40868 18624
rect 40920 18572 40926 18624
rect 42886 18572 42892 18624
rect 42944 18612 42950 18624
rect 43346 18612 43352 18624
rect 42944 18584 43352 18612
rect 42944 18572 42950 18584
rect 43346 18572 43352 18584
rect 43404 18612 43410 18624
rect 43441 18615 43499 18621
rect 43441 18612 43453 18615
rect 43404 18584 43453 18612
rect 43404 18572 43410 18584
rect 43441 18581 43453 18584
rect 43487 18581 43499 18615
rect 43441 18575 43499 18581
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 23385 18411 23443 18417
rect 23385 18377 23397 18411
rect 23431 18408 23443 18411
rect 26050 18408 26056 18420
rect 23431 18380 26056 18408
rect 23431 18377 23443 18380
rect 23385 18371 23443 18377
rect 26050 18368 26056 18380
rect 26108 18368 26114 18420
rect 28626 18368 28632 18420
rect 28684 18368 28690 18420
rect 32306 18368 32312 18420
rect 32364 18408 32370 18420
rect 35250 18408 35256 18420
rect 32364 18380 35256 18408
rect 32364 18368 32370 18380
rect 35250 18368 35256 18380
rect 35308 18368 35314 18420
rect 35526 18368 35532 18420
rect 35584 18368 35590 18420
rect 38378 18368 38384 18420
rect 38436 18408 38442 18420
rect 39669 18411 39727 18417
rect 39669 18408 39681 18411
rect 38436 18380 39681 18408
rect 38436 18368 38442 18380
rect 39669 18377 39681 18380
rect 39715 18377 39727 18411
rect 39669 18371 39727 18377
rect 44358 18368 44364 18420
rect 44416 18368 44422 18420
rect 25038 18340 25044 18352
rect 23768 18312 25044 18340
rect 23658 18232 23664 18284
rect 23716 18272 23722 18284
rect 23768 18281 23796 18312
rect 25038 18300 25044 18312
rect 25096 18300 25102 18352
rect 30190 18340 30196 18352
rect 28000 18312 30196 18340
rect 23753 18275 23811 18281
rect 23753 18272 23765 18275
rect 23716 18244 23765 18272
rect 23716 18232 23722 18244
rect 23753 18241 23765 18244
rect 23799 18241 23811 18275
rect 23753 18235 23811 18241
rect 23845 18275 23903 18281
rect 23845 18241 23857 18275
rect 23891 18272 23903 18275
rect 25958 18272 25964 18284
rect 23891 18244 25964 18272
rect 23891 18241 23903 18244
rect 23845 18235 23903 18241
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 26605 18275 26663 18281
rect 26605 18241 26617 18275
rect 26651 18272 26663 18275
rect 27709 18275 27767 18281
rect 27709 18272 27721 18275
rect 26651 18244 27721 18272
rect 26651 18241 26663 18244
rect 26605 18235 26663 18241
rect 27709 18241 27721 18244
rect 27755 18241 27767 18275
rect 27709 18235 27767 18241
rect 24029 18207 24087 18213
rect 24029 18173 24041 18207
rect 24075 18204 24087 18207
rect 25222 18204 25228 18216
rect 24075 18176 25228 18204
rect 24075 18173 24087 18176
rect 24029 18167 24087 18173
rect 25222 18164 25228 18176
rect 25280 18164 25286 18216
rect 27798 18164 27804 18216
rect 27856 18164 27862 18216
rect 28000 18213 28028 18312
rect 30190 18300 30196 18312
rect 30248 18300 30254 18352
rect 30285 18343 30343 18349
rect 30285 18309 30297 18343
rect 30331 18340 30343 18343
rect 30374 18340 30380 18352
rect 30331 18312 30380 18340
rect 30331 18309 30343 18312
rect 30285 18303 30343 18309
rect 30374 18300 30380 18312
rect 30432 18300 30438 18352
rect 31018 18300 31024 18352
rect 31076 18300 31082 18352
rect 31570 18300 31576 18352
rect 31628 18340 31634 18352
rect 35437 18343 35495 18349
rect 35437 18340 35449 18343
rect 31628 18312 35449 18340
rect 31628 18300 31634 18312
rect 35437 18309 35449 18312
rect 35483 18309 35495 18343
rect 35437 18303 35495 18309
rect 37642 18300 37648 18352
rect 37700 18340 37706 18352
rect 37737 18343 37795 18349
rect 37737 18340 37749 18343
rect 37700 18312 37749 18340
rect 37700 18300 37706 18312
rect 37737 18309 37749 18312
rect 37783 18309 37795 18343
rect 37737 18303 37795 18309
rect 42886 18300 42892 18352
rect 42944 18300 42950 18352
rect 28442 18232 28448 18284
rect 28500 18272 28506 18284
rect 28997 18275 29055 18281
rect 28997 18272 29009 18275
rect 28500 18244 29009 18272
rect 28500 18232 28506 18244
rect 28997 18241 29009 18244
rect 29043 18241 29055 18275
rect 28997 18235 29055 18241
rect 29089 18275 29147 18281
rect 29089 18241 29101 18275
rect 29135 18272 29147 18275
rect 29914 18272 29920 18284
rect 29135 18244 29920 18272
rect 29135 18241 29147 18244
rect 29089 18235 29147 18241
rect 29914 18232 29920 18244
rect 29972 18232 29978 18284
rect 34425 18275 34483 18281
rect 34425 18241 34437 18275
rect 34471 18272 34483 18275
rect 36262 18272 36268 18284
rect 34471 18244 36268 18272
rect 34471 18241 34483 18244
rect 34425 18235 34483 18241
rect 36262 18232 36268 18244
rect 36320 18232 36326 18284
rect 38838 18232 38844 18284
rect 38896 18232 38902 18284
rect 39853 18275 39911 18281
rect 39853 18241 39865 18275
rect 39899 18272 39911 18275
rect 41138 18272 41144 18284
rect 39899 18244 41144 18272
rect 39899 18241 39911 18244
rect 39853 18235 39911 18241
rect 41138 18232 41144 18244
rect 41196 18232 41202 18284
rect 41414 18232 41420 18284
rect 41472 18272 41478 18284
rect 42613 18275 42671 18281
rect 42613 18272 42625 18275
rect 41472 18244 42625 18272
rect 41472 18232 41478 18244
rect 42613 18241 42625 18244
rect 42659 18241 42671 18275
rect 42613 18235 42671 18241
rect 43990 18232 43996 18284
rect 44048 18232 44054 18284
rect 45189 18275 45247 18281
rect 45189 18241 45201 18275
rect 45235 18241 45247 18275
rect 45189 18235 45247 18241
rect 47949 18275 48007 18281
rect 47949 18241 47961 18275
rect 47995 18241 48007 18275
rect 47949 18235 48007 18241
rect 27985 18207 28043 18213
rect 27985 18173 27997 18207
rect 28031 18173 28043 18207
rect 27985 18167 28043 18173
rect 29178 18164 29184 18216
rect 29236 18164 29242 18216
rect 29730 18164 29736 18216
rect 29788 18204 29794 18216
rect 30009 18207 30067 18213
rect 30009 18204 30021 18207
rect 29788 18176 30021 18204
rect 29788 18164 29794 18176
rect 30009 18173 30021 18176
rect 30055 18173 30067 18207
rect 30009 18167 30067 18173
rect 34330 18164 34336 18216
rect 34388 18204 34394 18216
rect 35621 18207 35679 18213
rect 35621 18204 35633 18207
rect 34388 18176 35633 18204
rect 34388 18164 34394 18176
rect 35621 18173 35633 18176
rect 35667 18173 35679 18207
rect 35621 18167 35679 18173
rect 37458 18164 37464 18216
rect 37516 18164 37522 18216
rect 40770 18204 40776 18216
rect 39132 18176 40776 18204
rect 25590 18028 25596 18080
rect 25648 18028 25654 18080
rect 27341 18071 27399 18077
rect 27341 18037 27353 18071
rect 27387 18068 27399 18071
rect 30466 18068 30472 18080
rect 27387 18040 30472 18068
rect 27387 18037 27399 18040
rect 27341 18031 27399 18037
rect 30466 18028 30472 18040
rect 30524 18028 30530 18080
rect 31757 18071 31815 18077
rect 31757 18037 31769 18071
rect 31803 18068 31815 18071
rect 32122 18068 32128 18080
rect 31803 18040 32128 18068
rect 31803 18037 31815 18040
rect 31757 18031 31815 18037
rect 32122 18028 32128 18040
rect 32180 18028 32186 18080
rect 32582 18028 32588 18080
rect 32640 18068 32646 18080
rect 34517 18071 34575 18077
rect 34517 18068 34529 18071
rect 32640 18040 34529 18068
rect 32640 18028 32646 18040
rect 34517 18037 34529 18040
rect 34563 18037 34575 18071
rect 34517 18031 34575 18037
rect 35069 18071 35127 18077
rect 35069 18037 35081 18071
rect 35115 18068 35127 18071
rect 39132 18068 39160 18176
rect 40770 18164 40776 18176
rect 40828 18164 40834 18216
rect 40862 18164 40868 18216
rect 40920 18204 40926 18216
rect 42061 18207 42119 18213
rect 42061 18204 42073 18207
rect 40920 18176 42073 18204
rect 40920 18164 40926 18176
rect 42061 18173 42073 18176
rect 42107 18173 42119 18207
rect 42061 18167 42119 18173
rect 43438 18164 43444 18216
rect 43496 18204 43502 18216
rect 45204 18204 45232 18235
rect 43496 18176 45232 18204
rect 43496 18164 43502 18176
rect 39209 18139 39267 18145
rect 39209 18105 39221 18139
rect 39255 18136 39267 18139
rect 39942 18136 39948 18148
rect 39255 18108 39948 18136
rect 39255 18105 39267 18108
rect 39209 18099 39267 18105
rect 39942 18096 39948 18108
rect 40000 18096 40006 18148
rect 45005 18139 45063 18145
rect 45005 18105 45017 18139
rect 45051 18136 45063 18139
rect 47964 18136 47992 18235
rect 49142 18164 49148 18216
rect 49200 18164 49206 18216
rect 45051 18108 47992 18136
rect 45051 18105 45063 18108
rect 45005 18099 45063 18105
rect 35115 18040 39160 18068
rect 35115 18037 35127 18040
rect 35069 18031 35127 18037
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 25682 17824 25688 17876
rect 25740 17864 25746 17876
rect 27614 17864 27620 17876
rect 25740 17836 27620 17864
rect 25740 17824 25746 17836
rect 27614 17824 27620 17836
rect 27672 17864 27678 17876
rect 28902 17864 28908 17876
rect 27672 17836 28908 17864
rect 27672 17824 27678 17836
rect 28902 17824 28908 17836
rect 28960 17824 28966 17876
rect 37090 17824 37096 17876
rect 37148 17864 37154 17876
rect 37185 17867 37243 17873
rect 37185 17864 37197 17867
rect 37148 17836 37197 17864
rect 37148 17824 37154 17836
rect 37185 17833 37197 17836
rect 37231 17833 37243 17867
rect 37185 17827 37243 17833
rect 39209 17867 39267 17873
rect 39209 17833 39221 17867
rect 39255 17864 39267 17867
rect 43438 17864 43444 17876
rect 39255 17836 43444 17864
rect 39255 17833 39267 17836
rect 39209 17827 39267 17833
rect 43438 17824 43444 17836
rect 43496 17824 43502 17876
rect 25222 17756 25228 17808
rect 25280 17796 25286 17808
rect 25280 17768 25544 17796
rect 25280 17756 25286 17768
rect 25406 17688 25412 17740
rect 25464 17688 25470 17740
rect 25516 17728 25544 17768
rect 34146 17756 34152 17808
rect 34204 17756 34210 17808
rect 40313 17799 40371 17805
rect 34348 17768 35572 17796
rect 27433 17731 27491 17737
rect 27433 17728 27445 17731
rect 25516 17700 27445 17728
rect 27433 17697 27445 17700
rect 27479 17728 27491 17731
rect 27614 17728 27620 17740
rect 27479 17700 27620 17728
rect 27479 17697 27491 17700
rect 27433 17691 27491 17697
rect 27614 17688 27620 17700
rect 27672 17688 27678 17740
rect 28537 17731 28595 17737
rect 28537 17697 28549 17731
rect 28583 17728 28595 17731
rect 32030 17728 32036 17740
rect 28583 17700 32036 17728
rect 28583 17697 28595 17700
rect 28537 17691 28595 17697
rect 32030 17688 32036 17700
rect 32088 17688 32094 17740
rect 28261 17663 28319 17669
rect 28261 17629 28273 17663
rect 28307 17660 28319 17663
rect 28718 17660 28724 17672
rect 28307 17632 28724 17660
rect 28307 17629 28319 17632
rect 28261 17623 28319 17629
rect 28718 17620 28724 17632
rect 28776 17620 28782 17672
rect 28994 17620 29000 17672
rect 29052 17660 29058 17672
rect 29917 17663 29975 17669
rect 29917 17660 29929 17663
rect 29052 17632 29929 17660
rect 29052 17620 29058 17632
rect 29917 17629 29929 17632
rect 29963 17629 29975 17663
rect 29917 17623 29975 17629
rect 33410 17620 33416 17672
rect 33468 17660 33474 17672
rect 34348 17669 34376 17768
rect 34514 17688 34520 17740
rect 34572 17728 34578 17740
rect 35437 17731 35495 17737
rect 35437 17728 35449 17731
rect 34572 17700 35449 17728
rect 34572 17688 34578 17700
rect 35437 17697 35449 17700
rect 35483 17697 35495 17731
rect 35544 17728 35572 17768
rect 40313 17765 40325 17799
rect 40359 17796 40371 17799
rect 42518 17796 42524 17808
rect 40359 17768 42524 17796
rect 40359 17765 40371 17768
rect 40313 17759 40371 17765
rect 42518 17756 42524 17768
rect 42576 17756 42582 17808
rect 49786 17796 49792 17808
rect 44100 17768 49792 17796
rect 37366 17728 37372 17740
rect 35544 17700 37372 17728
rect 35437 17691 35495 17697
rect 37366 17688 37372 17700
rect 37424 17688 37430 17740
rect 38654 17688 38660 17740
rect 38712 17728 38718 17740
rect 38712 17700 41184 17728
rect 38712 17688 38718 17700
rect 33689 17663 33747 17669
rect 33689 17660 33701 17663
rect 33468 17632 33701 17660
rect 33468 17620 33474 17632
rect 33689 17629 33701 17632
rect 33735 17629 33747 17663
rect 33689 17623 33747 17629
rect 34333 17663 34391 17669
rect 34333 17629 34345 17663
rect 34379 17629 34391 17663
rect 34333 17623 34391 17629
rect 36998 17620 37004 17672
rect 37056 17660 37062 17672
rect 39393 17663 39451 17669
rect 39393 17660 39405 17663
rect 37056 17632 39405 17660
rect 37056 17620 37062 17632
rect 39393 17629 39405 17632
rect 39439 17629 39451 17663
rect 39393 17623 39451 17629
rect 40402 17620 40408 17672
rect 40460 17660 40466 17672
rect 40497 17663 40555 17669
rect 40497 17660 40509 17663
rect 40460 17632 40509 17660
rect 40460 17620 40466 17632
rect 40497 17629 40509 17632
rect 40543 17629 40555 17663
rect 40497 17623 40555 17629
rect 41156 17656 41184 17700
rect 41322 17688 41328 17740
rect 41380 17728 41386 17740
rect 44100 17728 44128 17768
rect 49786 17756 49792 17768
rect 49844 17756 49850 17808
rect 49694 17728 49700 17740
rect 41380 17700 44128 17728
rect 44192 17700 49700 17728
rect 41380 17688 41386 17700
rect 41233 17663 41291 17669
rect 41233 17656 41245 17663
rect 41156 17629 41245 17656
rect 41279 17629 41291 17663
rect 41156 17628 41291 17629
rect 41233 17623 41291 17628
rect 42794 17620 42800 17672
rect 42852 17660 42858 17672
rect 44192 17669 44220 17700
rect 49694 17688 49700 17700
rect 49752 17688 49758 17740
rect 42889 17663 42947 17669
rect 42889 17660 42901 17663
rect 42852 17632 42901 17660
rect 42852 17620 42858 17632
rect 42889 17629 42901 17632
rect 42935 17629 42947 17663
rect 42889 17623 42947 17629
rect 44177 17663 44235 17669
rect 44177 17629 44189 17663
rect 44223 17629 44235 17663
rect 44177 17623 44235 17629
rect 45281 17663 45339 17669
rect 45281 17629 45293 17663
rect 45327 17660 45339 17663
rect 50062 17660 50068 17672
rect 45327 17632 50068 17660
rect 45327 17629 45339 17632
rect 45281 17623 45339 17629
rect 50062 17620 50068 17632
rect 50120 17620 50126 17672
rect 25685 17595 25743 17601
rect 25685 17561 25697 17595
rect 25731 17561 25743 17595
rect 27338 17592 27344 17604
rect 26910 17564 27344 17592
rect 25685 17555 25743 17561
rect 25700 17524 25728 17555
rect 27338 17552 27344 17564
rect 27396 17552 27402 17604
rect 33318 17592 33324 17604
rect 27908 17564 33324 17592
rect 27706 17524 27712 17536
rect 25700 17496 27712 17524
rect 27706 17484 27712 17496
rect 27764 17484 27770 17536
rect 27908 17533 27936 17564
rect 33318 17552 33324 17564
rect 33376 17552 33382 17604
rect 34054 17552 34060 17604
rect 34112 17592 34118 17604
rect 35713 17595 35771 17601
rect 35713 17592 35725 17595
rect 34112 17564 35725 17592
rect 34112 17552 34118 17564
rect 35713 17561 35725 17564
rect 35759 17561 35771 17595
rect 35713 17555 35771 17561
rect 36170 17552 36176 17604
rect 36228 17552 36234 17604
rect 44361 17595 44419 17601
rect 37016 17564 44312 17592
rect 27893 17527 27951 17533
rect 27893 17493 27905 17527
rect 27939 17493 27951 17527
rect 27893 17487 27951 17493
rect 28350 17484 28356 17536
rect 28408 17484 28414 17536
rect 28534 17484 28540 17536
rect 28592 17524 28598 17536
rect 34882 17524 34888 17536
rect 28592 17496 34888 17524
rect 28592 17484 28598 17496
rect 34882 17484 34888 17496
rect 34940 17524 34946 17536
rect 37016 17524 37044 17564
rect 34940 17496 37044 17524
rect 41049 17527 41107 17533
rect 34940 17484 34946 17496
rect 41049 17493 41061 17527
rect 41095 17524 41107 17527
rect 43530 17524 43536 17536
rect 41095 17496 43536 17524
rect 41095 17493 41107 17496
rect 41049 17487 41107 17493
rect 43530 17484 43536 17496
rect 43588 17484 43594 17536
rect 44284 17524 44312 17564
rect 44361 17561 44373 17595
rect 44407 17592 44419 17595
rect 44542 17592 44548 17604
rect 44407 17564 44548 17592
rect 44407 17561 44419 17564
rect 44361 17555 44419 17561
rect 44542 17552 44548 17564
rect 44600 17552 44606 17604
rect 45462 17552 45468 17604
rect 45520 17552 45526 17604
rect 49418 17524 49424 17536
rect 44284 17496 49424 17524
rect 49418 17484 49424 17496
rect 49476 17484 49482 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 20349 17323 20407 17329
rect 20349 17289 20361 17323
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 25041 17323 25099 17329
rect 25041 17289 25053 17323
rect 25087 17320 25099 17323
rect 25130 17320 25136 17332
rect 25087 17292 25136 17320
rect 25087 17289 25099 17292
rect 25041 17283 25099 17289
rect 20364 17252 20392 17283
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 25409 17323 25467 17329
rect 25409 17289 25421 17323
rect 25455 17320 25467 17323
rect 25590 17320 25596 17332
rect 25455 17292 25596 17320
rect 25455 17289 25467 17292
rect 25409 17283 25467 17289
rect 25590 17280 25596 17292
rect 25648 17280 25654 17332
rect 25958 17280 25964 17332
rect 26016 17320 26022 17332
rect 27893 17323 27951 17329
rect 27893 17320 27905 17323
rect 26016 17292 27905 17320
rect 26016 17280 26022 17292
rect 27893 17289 27905 17292
rect 27939 17289 27951 17323
rect 27893 17283 27951 17289
rect 28261 17323 28319 17329
rect 28261 17289 28273 17323
rect 28307 17320 28319 17323
rect 28534 17320 28540 17332
rect 28307 17292 28540 17320
rect 28307 17289 28319 17292
rect 28261 17283 28319 17289
rect 27154 17252 27160 17264
rect 20364 17224 27160 17252
rect 27154 17212 27160 17224
rect 27212 17212 27218 17264
rect 27433 17255 27491 17261
rect 27433 17221 27445 17255
rect 27479 17252 27491 17255
rect 28276 17252 28304 17283
rect 28534 17280 28540 17292
rect 28592 17280 28598 17332
rect 29457 17323 29515 17329
rect 29457 17289 29469 17323
rect 29503 17320 29515 17323
rect 30377 17323 30435 17329
rect 30377 17320 30389 17323
rect 29503 17292 30389 17320
rect 29503 17289 29515 17292
rect 29457 17283 29515 17289
rect 30377 17289 30389 17292
rect 30423 17320 30435 17323
rect 31754 17320 31760 17332
rect 30423 17292 31760 17320
rect 30423 17289 30435 17292
rect 30377 17283 30435 17289
rect 31754 17280 31760 17292
rect 31812 17280 31818 17332
rect 32493 17323 32551 17329
rect 32493 17320 32505 17323
rect 31864 17292 32505 17320
rect 27479 17224 28304 17252
rect 27479 17221 27491 17224
rect 27433 17215 27491 17221
rect 29178 17212 29184 17264
rect 29236 17252 29242 17264
rect 31864 17252 31892 17292
rect 32493 17289 32505 17292
rect 32539 17289 32551 17323
rect 32493 17283 32551 17289
rect 33045 17323 33103 17329
rect 33045 17289 33057 17323
rect 33091 17289 33103 17323
rect 33045 17283 33103 17289
rect 29236 17224 31892 17252
rect 29236 17212 29242 17224
rect 32030 17212 32036 17264
rect 32088 17252 32094 17264
rect 32401 17255 32459 17261
rect 32401 17252 32413 17255
rect 32088 17224 32413 17252
rect 32088 17212 32094 17224
rect 32401 17221 32413 17224
rect 32447 17221 32459 17255
rect 33060 17252 33088 17283
rect 33410 17280 33416 17332
rect 33468 17280 33474 17332
rect 37458 17280 37464 17332
rect 37516 17320 37522 17332
rect 38562 17320 38568 17332
rect 37516 17292 38568 17320
rect 37516 17280 37522 17292
rect 38562 17280 38568 17292
rect 38620 17320 38626 17332
rect 39666 17320 39672 17332
rect 38620 17292 39672 17320
rect 38620 17280 38626 17292
rect 39666 17280 39672 17292
rect 39724 17320 39730 17332
rect 39724 17292 44036 17320
rect 39724 17280 39730 17292
rect 36998 17252 37004 17264
rect 33060 17224 37004 17252
rect 32401 17215 32459 17221
rect 36998 17212 37004 17224
rect 37056 17212 37062 17264
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17184 20775 17187
rect 20990 17184 20996 17196
rect 20763 17156 20996 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 26234 17184 26240 17196
rect 22066 17156 26240 17184
rect 19794 17076 19800 17128
rect 19852 17116 19858 17128
rect 19889 17119 19947 17125
rect 19889 17116 19901 17119
rect 19852 17088 19901 17116
rect 19852 17076 19858 17088
rect 19889 17085 19901 17088
rect 19935 17116 19947 17119
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 19935 17088 20821 17116
rect 19935 17085 19947 17088
rect 19889 17079 19947 17085
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 20901 17119 20959 17125
rect 20901 17085 20913 17119
rect 20947 17116 20959 17119
rect 22066 17116 22094 17156
rect 26234 17144 26240 17156
rect 26292 17144 26298 17196
rect 29454 17184 29460 17196
rect 27540 17156 29460 17184
rect 20947 17088 22094 17116
rect 20947 17085 20959 17088
rect 20901 17079 20959 17085
rect 24854 17076 24860 17128
rect 24912 17116 24918 17128
rect 25501 17119 25559 17125
rect 25501 17116 25513 17119
rect 24912 17088 25513 17116
rect 24912 17076 24918 17088
rect 25501 17085 25513 17088
rect 25547 17085 25559 17119
rect 25501 17079 25559 17085
rect 25685 17119 25743 17125
rect 25685 17085 25697 17119
rect 25731 17116 25743 17119
rect 27540 17116 27568 17156
rect 29454 17144 29460 17156
rect 29512 17144 29518 17196
rect 30742 17144 30748 17196
rect 30800 17184 30806 17196
rect 30837 17187 30895 17193
rect 30837 17184 30849 17187
rect 30800 17156 30849 17184
rect 30800 17144 30806 17156
rect 30837 17153 30849 17156
rect 30883 17153 30895 17187
rect 30837 17147 30895 17153
rect 30926 17144 30932 17196
rect 30984 17144 30990 17196
rect 32122 17144 32128 17196
rect 32180 17184 32186 17196
rect 37476 17193 37504 17280
rect 40402 17252 40408 17264
rect 39500 17224 40408 17252
rect 37461 17187 37519 17193
rect 32180 17156 33640 17184
rect 32180 17144 32186 17156
rect 25731 17088 27568 17116
rect 25731 17085 25743 17088
rect 25685 17079 25743 17085
rect 27798 17076 27804 17128
rect 27856 17116 27862 17128
rect 28353 17119 28411 17125
rect 28353 17116 28365 17119
rect 27856 17088 28365 17116
rect 27856 17076 27862 17088
rect 28353 17085 28365 17088
rect 28399 17085 28411 17119
rect 28353 17079 28411 17085
rect 28534 17076 28540 17128
rect 28592 17076 28598 17128
rect 28626 17076 28632 17128
rect 28684 17116 28690 17128
rect 29549 17119 29607 17125
rect 29549 17116 29561 17119
rect 28684 17088 29561 17116
rect 28684 17076 28690 17088
rect 29549 17085 29561 17088
rect 29595 17085 29607 17119
rect 29549 17079 29607 17085
rect 29641 17119 29699 17125
rect 29641 17085 29653 17119
rect 29687 17085 29699 17119
rect 29641 17079 29699 17085
rect 27706 17008 27712 17060
rect 27764 17048 27770 17060
rect 28552 17048 28580 17076
rect 27764 17020 28580 17048
rect 27764 17008 27770 17020
rect 28718 17008 28724 17060
rect 28776 17048 28782 17060
rect 29656 17048 29684 17079
rect 30374 17076 30380 17128
rect 30432 17116 30438 17128
rect 33612 17125 33640 17156
rect 37461 17153 37473 17187
rect 37507 17153 37519 17187
rect 37461 17147 37519 17153
rect 38838 17144 38844 17196
rect 38896 17184 38902 17196
rect 39500 17184 39528 17224
rect 40402 17212 40408 17224
rect 40460 17212 40466 17264
rect 42886 17212 42892 17264
rect 42944 17252 42950 17264
rect 43073 17255 43131 17261
rect 43073 17252 43085 17255
rect 42944 17224 43085 17252
rect 42944 17212 42950 17224
rect 43073 17221 43085 17224
rect 43119 17221 43131 17255
rect 43073 17215 43131 17221
rect 38896 17156 39528 17184
rect 38896 17144 38902 17156
rect 39666 17144 39672 17196
rect 39724 17144 39730 17196
rect 44008 17193 44036 17292
rect 44082 17280 44088 17332
rect 44140 17320 44146 17332
rect 44140 17292 44404 17320
rect 44140 17280 44146 17292
rect 44266 17212 44272 17264
rect 44324 17212 44330 17264
rect 44376 17252 44404 17292
rect 44376 17224 44758 17252
rect 42061 17187 42119 17193
rect 42061 17153 42073 17187
rect 42107 17184 42119 17187
rect 42981 17187 43039 17193
rect 42981 17184 42993 17187
rect 42107 17156 42993 17184
rect 42107 17153 42119 17156
rect 42061 17147 42119 17153
rect 42981 17153 42993 17156
rect 43027 17153 43039 17187
rect 42981 17147 43039 17153
rect 43993 17187 44051 17193
rect 43993 17153 44005 17187
rect 44039 17153 44051 17187
rect 43993 17147 44051 17153
rect 45554 17144 45560 17196
rect 45612 17184 45618 17196
rect 47949 17187 48007 17193
rect 47949 17184 47961 17187
rect 45612 17156 47961 17184
rect 45612 17144 45618 17156
rect 47949 17153 47961 17156
rect 47995 17153 48007 17187
rect 47949 17147 48007 17153
rect 31021 17119 31079 17125
rect 31021 17116 31033 17119
rect 30432 17088 31033 17116
rect 30432 17076 30438 17088
rect 31021 17085 31033 17088
rect 31067 17085 31079 17119
rect 33505 17119 33563 17125
rect 33505 17116 33517 17119
rect 31021 17079 31079 17085
rect 31956 17088 33517 17116
rect 28776 17020 29684 17048
rect 30469 17051 30527 17057
rect 28776 17008 28782 17020
rect 30469 17017 30481 17051
rect 30515 17048 30527 17051
rect 31956 17048 31984 17088
rect 33505 17085 33517 17088
rect 33551 17085 33563 17119
rect 33505 17079 33563 17085
rect 33597 17119 33655 17125
rect 33597 17085 33609 17119
rect 33643 17085 33655 17119
rect 33597 17079 33655 17085
rect 37734 17076 37740 17128
rect 37792 17076 37798 17128
rect 37826 17076 37832 17128
rect 37884 17116 37890 17128
rect 39209 17119 39267 17125
rect 39209 17116 39221 17119
rect 37884 17088 39221 17116
rect 37884 17076 37890 17088
rect 39209 17085 39221 17088
rect 39255 17085 39267 17119
rect 39209 17079 39267 17085
rect 39942 17076 39948 17128
rect 40000 17076 40006 17128
rect 40402 17076 40408 17128
rect 40460 17116 40466 17128
rect 43257 17119 43315 17125
rect 40460 17088 42748 17116
rect 40460 17076 40466 17088
rect 30515 17020 31984 17048
rect 30515 17017 30527 17020
rect 30469 17011 30527 17017
rect 39022 17008 39028 17060
rect 39080 17048 39086 17060
rect 39080 17020 39712 17048
rect 39080 17008 39086 17020
rect 29086 16940 29092 16992
rect 29144 16940 29150 16992
rect 31754 16940 31760 16992
rect 31812 16940 31818 16992
rect 39684 16980 39712 17020
rect 41046 17008 41052 17060
rect 41104 17048 41110 17060
rect 42613 17051 42671 17057
rect 42613 17048 42625 17051
rect 41104 17020 42625 17048
rect 41104 17008 41110 17020
rect 42613 17017 42625 17020
rect 42659 17017 42671 17051
rect 42720 17048 42748 17088
rect 43257 17085 43269 17119
rect 43303 17116 43315 17119
rect 43346 17116 43352 17128
rect 43303 17088 43352 17116
rect 43303 17085 43315 17088
rect 43257 17079 43315 17085
rect 43346 17076 43352 17088
rect 43404 17076 43410 17128
rect 49142 17076 49148 17128
rect 49200 17076 49206 17128
rect 43990 17048 43996 17060
rect 42720 17020 43996 17048
rect 42613 17011 42671 17017
rect 43990 17008 43996 17020
rect 44048 17008 44054 17060
rect 41417 16983 41475 16989
rect 41417 16980 41429 16983
rect 39684 16952 41429 16980
rect 41417 16949 41429 16952
rect 41463 16949 41475 16983
rect 41417 16943 41475 16949
rect 45741 16983 45799 16989
rect 45741 16949 45753 16983
rect 45787 16980 45799 16983
rect 46106 16980 46112 16992
rect 45787 16952 46112 16980
rect 45787 16949 45799 16952
rect 45741 16943 45799 16949
rect 46106 16940 46112 16952
rect 46164 16940 46170 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 20990 16736 20996 16788
rect 21048 16736 21054 16788
rect 22544 16779 22602 16785
rect 22544 16745 22556 16779
rect 22590 16776 22602 16779
rect 23842 16776 23848 16788
rect 22590 16748 23848 16776
rect 22590 16745 22602 16748
rect 22544 16739 22602 16745
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 25222 16736 25228 16788
rect 25280 16776 25286 16788
rect 29178 16776 29184 16788
rect 25280 16748 29184 16776
rect 25280 16736 25286 16748
rect 29178 16736 29184 16748
rect 29236 16736 29242 16788
rect 31938 16736 31944 16788
rect 31996 16776 32002 16788
rect 35802 16776 35808 16788
rect 31996 16748 35808 16776
rect 31996 16736 32002 16748
rect 35802 16736 35808 16748
rect 35860 16776 35866 16788
rect 41322 16776 41328 16788
rect 35860 16748 41328 16776
rect 35860 16736 35866 16748
rect 41322 16736 41328 16748
rect 41380 16736 41386 16788
rect 29086 16708 29092 16720
rect 25608 16680 29092 16708
rect 22281 16643 22339 16649
rect 22281 16609 22293 16643
rect 22327 16640 22339 16643
rect 23566 16640 23572 16652
rect 22327 16612 23572 16640
rect 22327 16609 22339 16612
rect 22281 16603 22339 16609
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 25608 16649 25636 16680
rect 29086 16668 29092 16680
rect 29144 16668 29150 16720
rect 33962 16668 33968 16720
rect 34020 16708 34026 16720
rect 37826 16708 37832 16720
rect 34020 16680 37832 16708
rect 34020 16668 34026 16680
rect 37826 16668 37832 16680
rect 37884 16668 37890 16720
rect 25593 16643 25651 16649
rect 25593 16609 25605 16643
rect 25639 16609 25651 16643
rect 25593 16603 25651 16609
rect 25682 16600 25688 16652
rect 25740 16600 25746 16652
rect 27154 16600 27160 16652
rect 27212 16600 27218 16652
rect 27341 16643 27399 16649
rect 27341 16609 27353 16643
rect 27387 16640 27399 16643
rect 27522 16640 27528 16652
rect 27387 16612 27528 16640
rect 27387 16609 27399 16612
rect 27341 16603 27399 16609
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 27614 16600 27620 16652
rect 27672 16640 27678 16652
rect 28626 16640 28632 16652
rect 27672 16612 28632 16640
rect 27672 16600 27678 16612
rect 28626 16600 28632 16612
rect 28684 16600 28690 16652
rect 28813 16643 28871 16649
rect 28813 16609 28825 16643
rect 28859 16640 28871 16643
rect 29638 16640 29644 16652
rect 28859 16612 29644 16640
rect 28859 16609 28871 16612
rect 28813 16603 28871 16609
rect 29638 16600 29644 16612
rect 29696 16600 29702 16652
rect 29730 16600 29736 16652
rect 29788 16600 29794 16652
rect 30009 16643 30067 16649
rect 30009 16609 30021 16643
rect 30055 16640 30067 16643
rect 30055 16612 31892 16640
rect 30055 16609 30067 16612
rect 30009 16603 30067 16609
rect 25501 16575 25559 16581
rect 25501 16541 25513 16575
rect 25547 16572 25559 16575
rect 25774 16572 25780 16584
rect 25547 16544 25780 16572
rect 25547 16541 25559 16544
rect 25501 16535 25559 16541
rect 25774 16532 25780 16544
rect 25832 16572 25838 16584
rect 26510 16572 26516 16584
rect 25832 16544 26516 16572
rect 25832 16532 25838 16544
rect 26510 16532 26516 16544
rect 26568 16532 26574 16584
rect 28537 16575 28595 16581
rect 28537 16541 28549 16575
rect 28583 16572 28595 16575
rect 28994 16572 29000 16584
rect 28583 16544 29000 16572
rect 28583 16541 28595 16544
rect 28537 16535 28595 16541
rect 28994 16532 29000 16544
rect 29052 16532 29058 16584
rect 31018 16532 31024 16584
rect 31076 16572 31082 16584
rect 31076 16544 31754 16572
rect 31076 16532 31082 16544
rect 24762 16504 24768 16516
rect 23782 16476 24768 16504
rect 24762 16464 24768 16476
rect 24820 16464 24826 16516
rect 26786 16504 26792 16516
rect 25148 16476 26792 16504
rect 24029 16439 24087 16445
rect 24029 16405 24041 16439
rect 24075 16436 24087 16439
rect 24118 16436 24124 16448
rect 24075 16408 24124 16436
rect 24075 16405 24087 16408
rect 24029 16399 24087 16405
rect 24118 16396 24124 16408
rect 24176 16396 24182 16448
rect 25148 16445 25176 16476
rect 26786 16464 26792 16476
rect 26844 16464 26850 16516
rect 27338 16464 27344 16516
rect 27396 16504 27402 16516
rect 29638 16504 29644 16516
rect 27396 16476 29644 16504
rect 27396 16464 27402 16476
rect 29638 16464 29644 16476
rect 29696 16464 29702 16516
rect 25133 16439 25191 16445
rect 25133 16405 25145 16439
rect 25179 16405 25191 16439
rect 25133 16399 25191 16405
rect 26694 16396 26700 16448
rect 26752 16396 26758 16448
rect 27062 16396 27068 16448
rect 27120 16396 27126 16448
rect 28169 16439 28227 16445
rect 28169 16405 28181 16439
rect 28215 16436 28227 16439
rect 29270 16436 29276 16448
rect 28215 16408 29276 16436
rect 28215 16405 28227 16408
rect 28169 16399 28227 16405
rect 29270 16396 29276 16408
rect 29328 16396 29334 16448
rect 30374 16396 30380 16448
rect 30432 16436 30438 16448
rect 31481 16439 31539 16445
rect 31481 16436 31493 16439
rect 30432 16408 31493 16436
rect 30432 16396 30438 16408
rect 31481 16405 31493 16408
rect 31527 16405 31539 16439
rect 31726 16436 31754 16544
rect 31864 16504 31892 16612
rect 31938 16600 31944 16652
rect 31996 16600 32002 16652
rect 32217 16643 32275 16649
rect 32217 16609 32229 16643
rect 32263 16640 32275 16643
rect 34330 16640 34336 16652
rect 32263 16612 34336 16640
rect 32263 16609 32275 16612
rect 32217 16603 32275 16609
rect 34330 16600 34336 16612
rect 34388 16600 34394 16652
rect 36541 16643 36599 16649
rect 36541 16609 36553 16643
rect 36587 16640 36599 16643
rect 36722 16640 36728 16652
rect 36587 16612 36728 16640
rect 36587 16609 36599 16612
rect 36541 16603 36599 16609
rect 36722 16600 36728 16612
rect 36780 16600 36786 16652
rect 38470 16600 38476 16652
rect 38528 16600 38534 16652
rect 38657 16643 38715 16649
rect 38657 16609 38669 16643
rect 38703 16640 38715 16643
rect 39942 16640 39948 16652
rect 38703 16612 39948 16640
rect 38703 16609 38715 16612
rect 38657 16603 38715 16609
rect 39942 16600 39948 16612
rect 40000 16600 40006 16652
rect 42610 16600 42616 16652
rect 42668 16640 42674 16652
rect 42705 16643 42763 16649
rect 42705 16640 42717 16643
rect 42668 16612 42717 16640
rect 42668 16600 42674 16612
rect 42705 16609 42717 16612
rect 42751 16609 42763 16643
rect 42705 16603 42763 16609
rect 42889 16643 42947 16649
rect 42889 16609 42901 16643
rect 42935 16640 42947 16643
rect 46106 16640 46112 16652
rect 42935 16612 46112 16640
rect 42935 16609 42947 16612
rect 42889 16603 42947 16609
rect 46106 16600 46112 16612
rect 46164 16600 46170 16652
rect 33318 16532 33324 16584
rect 33376 16572 33382 16584
rect 35066 16572 35072 16584
rect 33376 16544 35072 16572
rect 33376 16532 33382 16544
rect 35066 16532 35072 16544
rect 35124 16532 35130 16584
rect 35529 16575 35587 16581
rect 35529 16541 35541 16575
rect 35575 16541 35587 16575
rect 35529 16535 35587 16541
rect 36357 16575 36415 16581
rect 36357 16541 36369 16575
rect 36403 16572 36415 16575
rect 37182 16572 37188 16584
rect 36403 16544 37188 16572
rect 36403 16541 36415 16544
rect 36357 16535 36415 16541
rect 32122 16504 32128 16516
rect 31864 16476 32128 16504
rect 32122 16464 32128 16476
rect 32180 16464 32186 16516
rect 35434 16504 35440 16516
rect 33612 16476 35440 16504
rect 32858 16436 32864 16448
rect 31726 16408 32864 16436
rect 31481 16399 31539 16405
rect 32858 16396 32864 16408
rect 32916 16396 32922 16448
rect 32950 16396 32956 16448
rect 33008 16436 33014 16448
rect 33612 16436 33640 16476
rect 35434 16464 35440 16476
rect 35492 16464 35498 16516
rect 35544 16504 35572 16535
rect 37182 16532 37188 16544
rect 37240 16532 37246 16584
rect 40221 16575 40279 16581
rect 40221 16541 40233 16575
rect 40267 16572 40279 16575
rect 40310 16572 40316 16584
rect 40267 16544 40316 16572
rect 40267 16541 40279 16544
rect 40221 16535 40279 16541
rect 40310 16532 40316 16544
rect 40368 16532 40374 16584
rect 44450 16532 44456 16584
rect 44508 16572 44514 16584
rect 47949 16575 48007 16581
rect 47949 16572 47961 16575
rect 44508 16544 47961 16572
rect 44508 16532 44514 16544
rect 47949 16541 47961 16544
rect 47995 16541 48007 16575
rect 47949 16535 48007 16541
rect 36906 16504 36912 16516
rect 35544 16476 36912 16504
rect 36906 16464 36912 16476
rect 36964 16464 36970 16516
rect 37366 16464 37372 16516
rect 37424 16504 37430 16516
rect 38381 16507 38439 16513
rect 38381 16504 38393 16507
rect 37424 16476 38393 16504
rect 37424 16464 37430 16476
rect 38381 16473 38393 16476
rect 38427 16473 38439 16507
rect 40494 16504 40500 16516
rect 38381 16467 38439 16473
rect 39960 16476 40500 16504
rect 33008 16408 33640 16436
rect 33689 16439 33747 16445
rect 33008 16396 33014 16408
rect 33689 16405 33701 16439
rect 33735 16436 33747 16439
rect 33870 16436 33876 16448
rect 33735 16408 33876 16436
rect 33735 16405 33747 16408
rect 33689 16399 33747 16405
rect 33870 16396 33876 16408
rect 33928 16396 33934 16448
rect 35345 16439 35403 16445
rect 35345 16405 35357 16439
rect 35391 16436 35403 16439
rect 35526 16436 35532 16448
rect 35391 16408 35532 16436
rect 35391 16405 35403 16408
rect 35345 16399 35403 16405
rect 35526 16396 35532 16408
rect 35584 16396 35590 16448
rect 38013 16439 38071 16445
rect 38013 16405 38025 16439
rect 38059 16436 38071 16439
rect 39960 16436 39988 16476
rect 40494 16464 40500 16476
rect 40552 16464 40558 16516
rect 42613 16507 42671 16513
rect 42613 16473 42625 16507
rect 42659 16504 42671 16507
rect 42794 16504 42800 16516
rect 42659 16476 42800 16504
rect 42659 16473 42671 16476
rect 42613 16467 42671 16473
rect 42794 16464 42800 16476
rect 42852 16464 42858 16516
rect 49142 16464 49148 16516
rect 49200 16464 49206 16516
rect 38059 16408 39988 16436
rect 38059 16405 38071 16408
rect 38013 16399 38071 16405
rect 40034 16396 40040 16448
rect 40092 16396 40098 16448
rect 40218 16396 40224 16448
rect 40276 16436 40282 16448
rect 42245 16439 42303 16445
rect 42245 16436 42257 16439
rect 40276 16408 42257 16436
rect 40276 16396 40282 16408
rect 42245 16405 42257 16408
rect 42291 16405 42303 16439
rect 42245 16399 42303 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 27706 16192 27712 16244
rect 27764 16232 27770 16244
rect 28258 16232 28264 16244
rect 27764 16204 28264 16232
rect 27764 16192 27770 16204
rect 28258 16192 28264 16204
rect 28316 16192 28322 16244
rect 31754 16192 31760 16244
rect 31812 16232 31818 16244
rect 32677 16235 32735 16241
rect 32677 16232 32689 16235
rect 31812 16204 32689 16232
rect 31812 16192 31818 16204
rect 32677 16201 32689 16204
rect 32723 16201 32735 16235
rect 34514 16232 34520 16244
rect 32677 16195 32735 16201
rect 33612 16204 34520 16232
rect 24118 16124 24124 16176
rect 24176 16164 24182 16176
rect 24765 16167 24823 16173
rect 24765 16164 24777 16167
rect 24176 16136 24777 16164
rect 24176 16124 24182 16136
rect 24765 16133 24777 16136
rect 24811 16133 24823 16167
rect 27338 16164 27344 16176
rect 25990 16150 27344 16164
rect 24765 16127 24823 16133
rect 25976 16136 27344 16150
rect 23566 15988 23572 16040
rect 23624 16028 23630 16040
rect 24486 16028 24492 16040
rect 23624 16000 24492 16028
rect 23624 15988 23630 16000
rect 24486 15988 24492 16000
rect 24544 15988 24550 16040
rect 24762 15988 24768 16040
rect 24820 16028 24826 16040
rect 25976 16028 26004 16136
rect 27338 16124 27344 16136
rect 27396 16124 27402 16176
rect 29638 16164 29644 16176
rect 29578 16136 29644 16164
rect 29638 16124 29644 16136
rect 29696 16164 29702 16176
rect 31018 16164 31024 16176
rect 29696 16136 31024 16164
rect 29696 16124 29702 16136
rect 31018 16124 31024 16136
rect 31076 16124 31082 16176
rect 33612 16164 33640 16204
rect 34514 16192 34520 16204
rect 34572 16192 34578 16244
rect 34790 16192 34796 16244
rect 34848 16232 34854 16244
rect 35253 16235 35311 16241
rect 35253 16232 35265 16235
rect 34848 16204 35265 16232
rect 34848 16192 34854 16204
rect 35253 16201 35265 16204
rect 35299 16201 35311 16235
rect 35253 16195 35311 16201
rect 35066 16164 35072 16176
rect 33520 16136 33640 16164
rect 35006 16136 35072 16164
rect 33520 16105 33548 16136
rect 35066 16124 35072 16136
rect 35124 16164 35130 16176
rect 36170 16164 36176 16176
rect 35124 16136 36176 16164
rect 35124 16124 35130 16136
rect 36170 16124 36176 16136
rect 36228 16124 36234 16176
rect 33505 16099 33563 16105
rect 33505 16065 33517 16099
rect 33551 16065 33563 16099
rect 33505 16059 33563 16065
rect 37550 16056 37556 16108
rect 37608 16096 37614 16108
rect 37645 16099 37703 16105
rect 37645 16096 37657 16099
rect 37608 16068 37657 16096
rect 37608 16056 37614 16068
rect 37645 16065 37657 16068
rect 37691 16065 37703 16099
rect 37645 16059 37703 16065
rect 38933 16099 38991 16105
rect 38933 16065 38945 16099
rect 38979 16096 38991 16099
rect 39390 16096 39396 16108
rect 38979 16068 39396 16096
rect 38979 16065 38991 16068
rect 38933 16059 38991 16065
rect 39390 16056 39396 16068
rect 39448 16056 39454 16108
rect 40770 16056 40776 16108
rect 40828 16056 40834 16108
rect 24820 16000 26004 16028
rect 26513 16031 26571 16037
rect 24820 15988 24826 16000
rect 26513 15997 26525 16031
rect 26559 16028 26571 16031
rect 27522 16028 27528 16040
rect 26559 16000 27528 16028
rect 26559 15997 26571 16000
rect 26513 15991 26571 15997
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 27706 15988 27712 16040
rect 27764 16028 27770 16040
rect 28077 16031 28135 16037
rect 28077 16028 28089 16031
rect 27764 16000 28089 16028
rect 27764 15988 27770 16000
rect 28077 15997 28089 16000
rect 28123 15997 28135 16031
rect 28077 15991 28135 15997
rect 28353 16031 28411 16037
rect 28353 15997 28365 16031
rect 28399 16028 28411 16031
rect 28718 16028 28724 16040
rect 28399 16000 28724 16028
rect 28399 15997 28411 16000
rect 28353 15991 28411 15997
rect 28718 15988 28724 16000
rect 28776 15988 28782 16040
rect 28902 15988 28908 16040
rect 28960 16028 28966 16040
rect 30101 16031 30159 16037
rect 30101 16028 30113 16031
rect 28960 16000 30113 16028
rect 28960 15988 28966 16000
rect 30101 15997 30113 16000
rect 30147 16028 30159 16031
rect 30466 16028 30472 16040
rect 30147 16000 30472 16028
rect 30147 15997 30159 16000
rect 30101 15991 30159 15997
rect 30466 15988 30472 16000
rect 30524 15988 30530 16040
rect 32030 15988 32036 16040
rect 32088 16028 32094 16040
rect 32769 16031 32827 16037
rect 32769 16028 32781 16031
rect 32088 16000 32781 16028
rect 32088 15988 32094 16000
rect 32769 15997 32781 16000
rect 32815 15997 32827 16031
rect 32769 15991 32827 15997
rect 32950 15988 32956 16040
rect 33008 15988 33014 16040
rect 33781 16031 33839 16037
rect 33781 15997 33793 16031
rect 33827 16028 33839 16031
rect 34790 16028 34796 16040
rect 33827 16000 34796 16028
rect 33827 15997 33839 16000
rect 33781 15991 33839 15997
rect 34790 15988 34796 16000
rect 34848 15988 34854 16040
rect 35986 15960 35992 15972
rect 34808 15932 35992 15960
rect 32309 15895 32367 15901
rect 32309 15861 32321 15895
rect 32355 15892 32367 15895
rect 34808 15892 34836 15932
rect 35986 15920 35992 15932
rect 36044 15920 36050 15972
rect 32355 15864 34836 15892
rect 37461 15895 37519 15901
rect 32355 15861 32367 15864
rect 32309 15855 32367 15861
rect 37461 15861 37473 15895
rect 37507 15892 37519 15895
rect 37550 15892 37556 15904
rect 37507 15864 37556 15892
rect 37507 15861 37519 15864
rect 37461 15855 37519 15861
rect 37550 15852 37556 15864
rect 37608 15852 37614 15904
rect 38286 15852 38292 15904
rect 38344 15892 38350 15904
rect 38749 15895 38807 15901
rect 38749 15892 38761 15895
rect 38344 15864 38761 15892
rect 38344 15852 38350 15864
rect 38749 15861 38761 15864
rect 38795 15861 38807 15895
rect 38749 15855 38807 15861
rect 40589 15895 40647 15901
rect 40589 15861 40601 15895
rect 40635 15892 40647 15895
rect 42702 15892 42708 15904
rect 40635 15864 42708 15892
rect 40635 15861 40647 15864
rect 40589 15855 40647 15861
rect 42702 15852 42708 15864
rect 42760 15852 42766 15904
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 23290 15648 23296 15700
rect 23348 15648 23354 15700
rect 26970 15648 26976 15700
rect 27028 15688 27034 15700
rect 27801 15691 27859 15697
rect 27801 15688 27813 15691
rect 27028 15660 27813 15688
rect 27028 15648 27034 15660
rect 27801 15657 27813 15660
rect 27847 15657 27859 15691
rect 27801 15651 27859 15657
rect 31113 15691 31171 15697
rect 31113 15657 31125 15691
rect 31159 15688 31171 15691
rect 31570 15688 31576 15700
rect 31159 15660 31576 15688
rect 31159 15657 31171 15660
rect 31113 15651 31171 15657
rect 31570 15648 31576 15660
rect 31628 15648 31634 15700
rect 37369 15691 37427 15697
rect 37369 15657 37381 15691
rect 37415 15688 37427 15691
rect 37734 15688 37740 15700
rect 37415 15660 37740 15688
rect 37415 15657 37427 15660
rect 37369 15651 37427 15657
rect 37734 15648 37740 15660
rect 37792 15648 37798 15700
rect 23842 15512 23848 15564
rect 23900 15512 23906 15564
rect 24486 15512 24492 15564
rect 24544 15552 24550 15564
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 24544 15524 25237 15552
rect 24544 15512 24550 15524
rect 25225 15521 25237 15524
rect 25271 15552 25283 15555
rect 26234 15552 26240 15564
rect 25271 15524 26240 15552
rect 25271 15521 25283 15524
rect 25225 15515 25283 15521
rect 26234 15512 26240 15524
rect 26292 15512 26298 15564
rect 28258 15512 28264 15564
rect 28316 15552 28322 15564
rect 28353 15555 28411 15561
rect 28353 15552 28365 15555
rect 28316 15524 28365 15552
rect 28316 15512 28322 15524
rect 28353 15521 28365 15524
rect 28399 15521 28411 15555
rect 28353 15515 28411 15521
rect 31662 15512 31668 15564
rect 31720 15512 31726 15564
rect 34514 15512 34520 15564
rect 34572 15552 34578 15564
rect 35618 15552 35624 15564
rect 34572 15524 35624 15552
rect 34572 15512 34578 15524
rect 35618 15512 35624 15524
rect 35676 15512 35682 15564
rect 35894 15512 35900 15564
rect 35952 15512 35958 15564
rect 37752 15552 37780 15648
rect 37829 15623 37887 15629
rect 37829 15589 37841 15623
rect 37875 15620 37887 15623
rect 40862 15620 40868 15632
rect 37875 15592 40868 15620
rect 37875 15589 37887 15592
rect 37829 15583 37887 15589
rect 40862 15580 40868 15592
rect 40920 15580 40926 15632
rect 44453 15623 44511 15629
rect 44453 15589 44465 15623
rect 44499 15620 44511 15623
rect 45554 15620 45560 15632
rect 44499 15592 45560 15620
rect 44499 15589 44511 15592
rect 44453 15583 44511 15589
rect 45554 15580 45560 15592
rect 45612 15580 45618 15632
rect 38381 15555 38439 15561
rect 38381 15552 38393 15555
rect 37752 15524 38393 15552
rect 38381 15521 38393 15524
rect 38427 15521 38439 15555
rect 38381 15515 38439 15521
rect 27249 15487 27307 15493
rect 27249 15453 27261 15487
rect 27295 15484 27307 15487
rect 28718 15484 28724 15496
rect 27295 15456 28724 15484
rect 27295 15453 27307 15456
rect 27249 15447 27307 15453
rect 28718 15444 28724 15456
rect 28776 15444 28782 15496
rect 30650 15444 30656 15496
rect 30708 15444 30714 15496
rect 31481 15487 31539 15493
rect 31481 15453 31493 15487
rect 31527 15484 31539 15487
rect 32493 15487 32551 15493
rect 32493 15484 32505 15487
rect 31527 15456 32505 15484
rect 31527 15453 31539 15456
rect 31481 15447 31539 15453
rect 32493 15453 32505 15456
rect 32539 15453 32551 15487
rect 32493 15447 32551 15453
rect 33597 15487 33655 15493
rect 33597 15453 33609 15487
rect 33643 15484 33655 15487
rect 34238 15484 34244 15496
rect 33643 15456 34244 15484
rect 33643 15453 33655 15456
rect 33597 15447 33655 15453
rect 34238 15444 34244 15456
rect 34296 15444 34302 15496
rect 37274 15444 37280 15496
rect 37332 15484 37338 15496
rect 38289 15487 38347 15493
rect 38289 15484 38301 15487
rect 37332 15456 38301 15484
rect 37332 15444 37338 15456
rect 38289 15453 38301 15456
rect 38335 15453 38347 15487
rect 38289 15447 38347 15453
rect 39117 15487 39175 15493
rect 39117 15453 39129 15487
rect 39163 15484 39175 15487
rect 43622 15484 43628 15496
rect 39163 15456 43628 15484
rect 39163 15453 39175 15456
rect 39117 15447 39175 15453
rect 43622 15444 43628 15456
rect 43680 15444 43686 15496
rect 44726 15444 44732 15496
rect 44784 15484 44790 15496
rect 47949 15487 48007 15493
rect 47949 15484 47961 15487
rect 44784 15456 47961 15484
rect 44784 15444 44790 15456
rect 47949 15453 47961 15456
rect 47995 15453 48007 15487
rect 47949 15447 48007 15453
rect 49142 15444 49148 15496
rect 49200 15444 49206 15496
rect 23382 15376 23388 15428
rect 23440 15416 23446 15428
rect 23753 15419 23811 15425
rect 23753 15416 23765 15419
rect 23440 15388 23765 15416
rect 23440 15376 23446 15388
rect 23753 15385 23765 15388
rect 23799 15385 23811 15419
rect 23753 15379 23811 15385
rect 25498 15376 25504 15428
rect 25556 15376 25562 15428
rect 27338 15416 27344 15428
rect 26726 15388 27344 15416
rect 27338 15376 27344 15388
rect 27396 15376 27402 15428
rect 28169 15419 28227 15425
rect 28169 15385 28181 15419
rect 28215 15416 28227 15419
rect 29546 15416 29552 15428
rect 28215 15388 29552 15416
rect 28215 15385 28227 15388
rect 28169 15379 28227 15385
rect 29546 15376 29552 15388
rect 29604 15376 29610 15428
rect 30834 15376 30840 15428
rect 30892 15416 30898 15428
rect 31573 15419 31631 15425
rect 31573 15416 31585 15419
rect 30892 15388 31585 15416
rect 30892 15376 30898 15388
rect 31573 15385 31585 15388
rect 31619 15385 31631 15419
rect 31573 15379 31631 15385
rect 33502 15376 33508 15428
rect 33560 15416 33566 15428
rect 33560 15388 33824 15416
rect 33560 15376 33566 15388
rect 23661 15351 23719 15357
rect 23661 15317 23673 15351
rect 23707 15348 23719 15351
rect 25866 15348 25872 15360
rect 23707 15320 25872 15348
rect 23707 15317 23719 15320
rect 23661 15311 23719 15317
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 28261 15351 28319 15357
rect 28261 15317 28273 15351
rect 28307 15348 28319 15351
rect 29822 15348 29828 15360
rect 28307 15320 29828 15348
rect 28307 15317 28319 15320
rect 28261 15311 28319 15317
rect 29822 15308 29828 15320
rect 29880 15308 29886 15360
rect 33686 15308 33692 15360
rect 33744 15308 33750 15360
rect 33796 15348 33824 15388
rect 36354 15376 36360 15428
rect 36412 15376 36418 15428
rect 37458 15376 37464 15428
rect 37516 15416 37522 15428
rect 37516 15388 38424 15416
rect 37516 15376 37522 15388
rect 38197 15351 38255 15357
rect 38197 15348 38209 15351
rect 33796 15320 38209 15348
rect 38197 15317 38209 15320
rect 38243 15317 38255 15351
rect 38396 15348 38424 15388
rect 38654 15376 38660 15428
rect 38712 15416 38718 15428
rect 44269 15419 44327 15425
rect 44269 15416 44281 15419
rect 38712 15388 44281 15416
rect 38712 15376 38718 15388
rect 44269 15385 44281 15388
rect 44315 15385 44327 15419
rect 44269 15379 44327 15385
rect 45557 15419 45615 15425
rect 45557 15385 45569 15419
rect 45603 15385 45615 15419
rect 45557 15379 45615 15385
rect 45741 15419 45799 15425
rect 45741 15385 45753 15419
rect 45787 15416 45799 15419
rect 47762 15416 47768 15428
rect 45787 15388 47768 15416
rect 45787 15385 45799 15388
rect 45741 15379 45799 15385
rect 39209 15351 39267 15357
rect 39209 15348 39221 15351
rect 38396 15320 39221 15348
rect 38197 15311 38255 15317
rect 39209 15317 39221 15320
rect 39255 15317 39267 15351
rect 39209 15311 39267 15317
rect 42518 15308 42524 15360
rect 42576 15348 42582 15360
rect 45572 15348 45600 15379
rect 47762 15376 47768 15388
rect 47820 15376 47826 15428
rect 42576 15320 45600 15348
rect 42576 15308 42582 15320
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 25133 15147 25191 15153
rect 25133 15113 25145 15147
rect 25179 15144 25191 15147
rect 25498 15144 25504 15156
rect 25179 15116 25504 15144
rect 25179 15113 25191 15116
rect 25133 15107 25191 15113
rect 25498 15104 25504 15116
rect 25556 15104 25562 15156
rect 27801 15147 27859 15153
rect 27801 15113 27813 15147
rect 27847 15144 27859 15147
rect 29181 15147 29239 15153
rect 29181 15144 29193 15147
rect 27847 15116 29193 15144
rect 27847 15113 27859 15116
rect 27801 15107 27859 15113
rect 29181 15113 29193 15116
rect 29227 15144 29239 15147
rect 30469 15147 30527 15153
rect 29227 15116 29684 15144
rect 29227 15113 29239 15116
rect 29181 15107 29239 15113
rect 23566 15076 23572 15088
rect 23400 15048 23572 15076
rect 23400 15017 23428 15048
rect 23566 15036 23572 15048
rect 23624 15036 23630 15088
rect 26234 15036 26240 15088
rect 26292 15076 26298 15088
rect 26421 15079 26479 15085
rect 26421 15076 26433 15079
rect 26292 15048 26433 15076
rect 26292 15036 26298 15048
rect 26421 15045 26433 15048
rect 26467 15045 26479 15079
rect 29656 15076 29684 15116
rect 30469 15113 30481 15147
rect 30515 15144 30527 15147
rect 30650 15144 30656 15156
rect 30515 15116 30656 15144
rect 30515 15113 30527 15116
rect 30469 15107 30527 15113
rect 30650 15104 30656 15116
rect 30708 15104 30714 15156
rect 32858 15144 32864 15156
rect 32416 15116 32864 15144
rect 29656 15048 30604 15076
rect 26421 15039 26479 15045
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 14977 23443 15011
rect 23385 14971 23443 14977
rect 24762 14968 24768 15020
rect 24820 14968 24826 15020
rect 25685 15011 25743 15017
rect 25685 14977 25697 15011
rect 25731 15008 25743 15011
rect 27430 15008 27436 15020
rect 25731 14980 27436 15008
rect 25731 14977 25743 14980
rect 25685 14971 25743 14977
rect 27430 14968 27436 14980
rect 27488 14968 27494 15020
rect 27522 14968 27528 15020
rect 27580 15008 27586 15020
rect 30576 15008 30604 15048
rect 31938 15036 31944 15088
rect 31996 15076 32002 15088
rect 32416 15076 32444 15116
rect 32858 15104 32864 15116
rect 32916 15144 32922 15156
rect 34514 15144 34520 15156
rect 32916 15116 34520 15144
rect 32916 15104 32922 15116
rect 34514 15104 34520 15116
rect 34572 15104 34578 15156
rect 37645 15147 37703 15153
rect 37645 15113 37657 15147
rect 37691 15144 37703 15147
rect 38654 15144 38660 15156
rect 37691 15116 38660 15144
rect 37691 15113 37703 15116
rect 37645 15107 37703 15113
rect 38654 15104 38660 15116
rect 38712 15104 38718 15156
rect 31996 15048 32444 15076
rect 31996 15036 32002 15048
rect 32122 15008 32128 15020
rect 27580 14980 29408 15008
rect 30576 14980 32128 15008
rect 27580 14968 27586 14980
rect 23661 14943 23719 14949
rect 23661 14909 23673 14943
rect 23707 14940 23719 14943
rect 25498 14940 25504 14952
rect 23707 14912 25504 14940
rect 23707 14909 23719 14912
rect 23661 14903 23719 14909
rect 25498 14900 25504 14912
rect 25556 14900 25562 14952
rect 29380 14949 29408 14980
rect 32122 14968 32128 14980
rect 32180 14968 32186 15020
rect 32324 15017 32352 15048
rect 33318 15036 33324 15088
rect 33376 15036 33382 15088
rect 34974 15076 34980 15088
rect 33888 15048 34980 15076
rect 32309 15011 32367 15017
rect 32309 14977 32321 15011
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 29273 14943 29331 14949
rect 29273 14909 29285 14943
rect 29319 14909 29331 14943
rect 29273 14903 29331 14909
rect 29365 14943 29423 14949
rect 29365 14909 29377 14943
rect 29411 14940 29423 14943
rect 30282 14940 30288 14952
rect 29411 14912 30288 14940
rect 29411 14909 29423 14912
rect 29365 14903 29423 14909
rect 25038 14832 25044 14884
rect 25096 14872 25102 14884
rect 28813 14875 28871 14881
rect 28813 14872 28825 14875
rect 25096 14844 28825 14872
rect 25096 14832 25102 14844
rect 28813 14841 28825 14844
rect 28859 14841 28871 14875
rect 28813 14835 28871 14841
rect 28258 14764 28264 14816
rect 28316 14804 28322 14816
rect 29288 14804 29316 14903
rect 30282 14900 30288 14912
rect 30340 14900 30346 14952
rect 30558 14900 30564 14952
rect 30616 14900 30622 14952
rect 30745 14943 30803 14949
rect 30745 14909 30757 14943
rect 30791 14940 30803 14943
rect 31846 14940 31852 14952
rect 30791 14912 31852 14940
rect 30791 14909 30803 14912
rect 30745 14903 30803 14909
rect 31846 14900 31852 14912
rect 31904 14900 31910 14952
rect 32585 14943 32643 14949
rect 32585 14909 32597 14943
rect 32631 14940 32643 14943
rect 33888 14940 33916 15048
rect 34974 15036 34980 15048
rect 35032 15076 35038 15088
rect 35342 15076 35348 15088
rect 35032 15048 35348 15076
rect 35032 15036 35038 15048
rect 35342 15036 35348 15048
rect 35400 15036 35406 15088
rect 35618 15036 35624 15088
rect 35676 15036 35682 15088
rect 36357 15079 36415 15085
rect 36357 15045 36369 15079
rect 36403 15076 36415 15079
rect 36538 15076 36544 15088
rect 36403 15048 36544 15076
rect 36403 15045 36415 15048
rect 36357 15039 36415 15045
rect 36538 15036 36544 15048
rect 36596 15036 36602 15088
rect 39022 15036 39028 15088
rect 39080 15036 39086 15088
rect 40402 15076 40408 15088
rect 40250 15048 40408 15076
rect 40402 15036 40408 15048
rect 40460 15036 40466 15088
rect 34885 15011 34943 15017
rect 34885 15008 34897 15011
rect 32631 14912 33916 14940
rect 33980 14980 34897 15008
rect 32631 14909 32643 14912
rect 32585 14903 32643 14909
rect 30101 14875 30159 14881
rect 30101 14841 30113 14875
rect 30147 14872 30159 14875
rect 32306 14872 32312 14884
rect 30147 14844 32312 14872
rect 30147 14841 30159 14844
rect 30101 14835 30159 14841
rect 32306 14832 32312 14844
rect 32364 14832 32370 14884
rect 30742 14804 30748 14816
rect 28316 14776 30748 14804
rect 28316 14764 28322 14776
rect 30742 14764 30748 14776
rect 30800 14764 30806 14816
rect 32398 14764 32404 14816
rect 32456 14804 32462 14816
rect 33980 14804 34008 14980
rect 34885 14977 34897 14980
rect 34931 15008 34943 15011
rect 36262 15008 36268 15020
rect 34931 14980 36268 15008
rect 34931 14977 34943 14980
rect 34885 14971 34943 14977
rect 36262 14968 36268 14980
rect 36320 14968 36326 15020
rect 37274 14968 37280 15020
rect 37332 15008 37338 15020
rect 37829 15011 37887 15017
rect 37829 15008 37841 15011
rect 37332 14980 37841 15008
rect 37332 14968 37338 14980
rect 37829 14977 37841 14980
rect 37875 14977 37887 15011
rect 37829 14971 37887 14977
rect 38562 14968 38568 15020
rect 38620 15008 38626 15020
rect 38749 15011 38807 15017
rect 38749 15008 38761 15011
rect 38620 14980 38761 15008
rect 38620 14968 38626 14980
rect 38749 14977 38761 14980
rect 38795 14977 38807 15011
rect 38749 14971 38807 14977
rect 43530 14968 43536 15020
rect 43588 15008 43594 15020
rect 46017 15011 46075 15017
rect 46017 15008 46029 15011
rect 43588 14980 46029 15008
rect 43588 14968 43594 14980
rect 46017 14977 46029 14980
rect 46063 14977 46075 15011
rect 46017 14971 46075 14977
rect 47946 14968 47952 15020
rect 48004 14968 48010 15020
rect 34054 14900 34060 14952
rect 34112 14900 34118 14952
rect 49142 14900 49148 14952
rect 49200 14900 49206 14952
rect 32456 14776 34008 14804
rect 32456 14764 32462 14776
rect 36446 14764 36452 14816
rect 36504 14764 36510 14816
rect 39390 14764 39396 14816
rect 39448 14804 39454 14816
rect 40497 14807 40555 14813
rect 40497 14804 40509 14807
rect 39448 14776 40509 14804
rect 39448 14764 39454 14776
rect 40497 14773 40509 14776
rect 40543 14773 40555 14807
rect 40497 14767 40555 14773
rect 45833 14807 45891 14813
rect 45833 14773 45845 14807
rect 45879 14804 45891 14807
rect 47854 14804 47860 14816
rect 45879 14776 47860 14804
rect 45879 14773 45891 14776
rect 45833 14767 45891 14773
rect 47854 14764 47860 14776
rect 47912 14764 47918 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 25314 14560 25320 14612
rect 25372 14600 25378 14612
rect 25593 14603 25651 14609
rect 25593 14600 25605 14603
rect 25372 14572 25605 14600
rect 25372 14560 25378 14572
rect 25593 14569 25605 14572
rect 25639 14569 25651 14603
rect 25593 14563 25651 14569
rect 28442 14560 28448 14612
rect 28500 14560 28506 14612
rect 30282 14560 30288 14612
rect 30340 14600 30346 14612
rect 31478 14600 31484 14612
rect 30340 14572 31484 14600
rect 30340 14560 30346 14572
rect 31478 14560 31484 14572
rect 31536 14560 31542 14612
rect 32122 14560 32128 14612
rect 32180 14600 32186 14612
rect 35342 14600 35348 14612
rect 32180 14572 35348 14600
rect 32180 14560 32186 14572
rect 35342 14560 35348 14572
rect 35400 14600 35406 14612
rect 45649 14603 45707 14609
rect 35400 14572 41414 14600
rect 35400 14560 35406 14572
rect 30190 14492 30196 14544
rect 30248 14532 30254 14544
rect 35066 14532 35072 14544
rect 30248 14504 35072 14532
rect 30248 14492 30254 14504
rect 35066 14492 35072 14504
rect 35124 14492 35130 14544
rect 35161 14535 35219 14541
rect 35161 14501 35173 14535
rect 35207 14532 35219 14535
rect 41230 14532 41236 14544
rect 35207 14504 41236 14532
rect 35207 14501 35219 14504
rect 35161 14495 35219 14501
rect 41230 14492 41236 14504
rect 41288 14492 41294 14544
rect 41386 14532 41414 14572
rect 45649 14569 45661 14603
rect 45695 14600 45707 14603
rect 47946 14600 47952 14612
rect 45695 14572 47952 14600
rect 45695 14569 45707 14572
rect 45649 14563 45707 14569
rect 47946 14560 47952 14572
rect 48004 14560 48010 14612
rect 49234 14532 49240 14544
rect 41386 14504 49240 14532
rect 49234 14492 49240 14504
rect 49292 14492 49298 14544
rect 23842 14424 23848 14476
rect 23900 14464 23906 14476
rect 26145 14467 26203 14473
rect 26145 14464 26157 14467
rect 23900 14436 26157 14464
rect 23900 14424 23906 14436
rect 26145 14433 26157 14436
rect 26191 14433 26203 14467
rect 26145 14427 26203 14433
rect 26786 14424 26792 14476
rect 26844 14464 26850 14476
rect 27157 14467 27215 14473
rect 27157 14464 27169 14467
rect 26844 14436 27169 14464
rect 26844 14424 26850 14436
rect 27157 14433 27169 14436
rect 27203 14433 27215 14467
rect 27157 14427 27215 14433
rect 27706 14424 27712 14476
rect 27764 14464 27770 14476
rect 28169 14467 28227 14473
rect 28169 14464 28181 14467
rect 27764 14436 28181 14464
rect 27764 14424 27770 14436
rect 28169 14433 28181 14436
rect 28215 14433 28227 14467
rect 28169 14427 28227 14433
rect 28902 14424 28908 14476
rect 28960 14464 28966 14476
rect 28997 14467 29055 14473
rect 28997 14464 29009 14467
rect 28960 14436 29009 14464
rect 28960 14424 28966 14436
rect 28997 14433 29009 14436
rect 29043 14433 29055 14467
rect 28997 14427 29055 14433
rect 31478 14424 31484 14476
rect 31536 14464 31542 14476
rect 32125 14467 32183 14473
rect 32125 14464 32137 14467
rect 31536 14436 32137 14464
rect 31536 14424 31542 14436
rect 32125 14433 32137 14436
rect 32171 14433 32183 14467
rect 32125 14427 32183 14433
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 35713 14467 35771 14473
rect 35713 14464 35725 14467
rect 34848 14436 35725 14464
rect 34848 14424 34854 14436
rect 35713 14433 35725 14436
rect 35759 14433 35771 14467
rect 35713 14427 35771 14433
rect 38105 14467 38163 14473
rect 38105 14433 38117 14467
rect 38151 14464 38163 14467
rect 38562 14464 38568 14476
rect 38151 14436 38568 14464
rect 38151 14433 38163 14436
rect 38105 14427 38163 14433
rect 38562 14424 38568 14436
rect 38620 14424 38626 14476
rect 39206 14424 39212 14476
rect 39264 14424 39270 14476
rect 39390 14424 39396 14476
rect 39448 14424 39454 14476
rect 41138 14464 41144 14476
rect 40512 14436 41144 14464
rect 25133 14399 25191 14405
rect 25133 14365 25145 14399
rect 25179 14396 25191 14399
rect 26234 14396 26240 14408
rect 25179 14368 26240 14396
rect 25179 14365 25191 14368
rect 25133 14359 25191 14365
rect 26234 14356 26240 14368
rect 26292 14356 26298 14408
rect 26970 14356 26976 14408
rect 27028 14356 27034 14408
rect 27430 14356 27436 14408
rect 27488 14356 27494 14408
rect 28442 14356 28448 14408
rect 28500 14396 28506 14408
rect 28810 14396 28816 14408
rect 28500 14368 28816 14396
rect 28500 14356 28506 14368
rect 28810 14356 28816 14368
rect 28868 14356 28874 14408
rect 30926 14356 30932 14408
rect 30984 14396 30990 14408
rect 32030 14396 32036 14408
rect 30984 14368 32036 14396
rect 30984 14356 30990 14368
rect 32030 14356 32036 14368
rect 32088 14356 32094 14408
rect 35529 14399 35587 14405
rect 35529 14365 35541 14399
rect 35575 14396 35587 14399
rect 36541 14399 36599 14405
rect 36541 14396 36553 14399
rect 35575 14368 36553 14396
rect 35575 14365 35587 14368
rect 35529 14359 35587 14365
rect 36541 14365 36553 14368
rect 36587 14365 36599 14399
rect 36541 14359 36599 14365
rect 39114 14356 39120 14408
rect 39172 14356 39178 14408
rect 25961 14331 26019 14337
rect 25961 14297 25973 14331
rect 26007 14328 26019 14331
rect 27338 14328 27344 14340
rect 26007 14300 27344 14328
rect 26007 14297 26019 14300
rect 25961 14291 26019 14297
rect 27338 14288 27344 14300
rect 27396 14288 27402 14340
rect 30561 14331 30619 14337
rect 30561 14297 30573 14331
rect 30607 14328 30619 14331
rect 30607 14300 31754 14328
rect 30607 14297 30619 14300
rect 30561 14291 30619 14297
rect 26053 14263 26111 14269
rect 26053 14229 26065 14263
rect 26099 14260 26111 14263
rect 26510 14260 26516 14272
rect 26099 14232 26516 14260
rect 26099 14229 26111 14232
rect 26053 14223 26111 14229
rect 26510 14220 26516 14232
rect 26568 14220 26574 14272
rect 26602 14220 26608 14272
rect 26660 14220 26666 14272
rect 26878 14220 26884 14272
rect 26936 14260 26942 14272
rect 27065 14263 27123 14269
rect 27065 14260 27077 14263
rect 26936 14232 27077 14260
rect 26936 14220 26942 14232
rect 27065 14229 27077 14232
rect 27111 14229 27123 14263
rect 27065 14223 27123 14229
rect 28810 14220 28816 14272
rect 28868 14220 28874 14272
rect 28902 14220 28908 14272
rect 28960 14220 28966 14272
rect 30926 14220 30932 14272
rect 30984 14260 30990 14272
rect 31021 14263 31079 14269
rect 31021 14260 31033 14263
rect 30984 14232 31033 14260
rect 30984 14220 30990 14232
rect 31021 14229 31033 14232
rect 31067 14229 31079 14263
rect 31021 14223 31079 14229
rect 31570 14220 31576 14272
rect 31628 14220 31634 14272
rect 31726 14260 31754 14300
rect 31846 14288 31852 14340
rect 31904 14328 31910 14340
rect 34698 14328 34704 14340
rect 31904 14300 34704 14328
rect 31904 14288 31910 14300
rect 34698 14288 34704 14300
rect 34756 14288 34762 14340
rect 34808 14300 35848 14328
rect 31941 14263 31999 14269
rect 31941 14260 31953 14263
rect 31726 14232 31953 14260
rect 31941 14229 31953 14232
rect 31987 14260 31999 14263
rect 34808 14260 34836 14300
rect 31987 14232 34836 14260
rect 31987 14229 31999 14232
rect 31941 14223 31999 14229
rect 35618 14220 35624 14272
rect 35676 14220 35682 14272
rect 35820 14260 35848 14300
rect 35894 14288 35900 14340
rect 35952 14328 35958 14340
rect 36262 14328 36268 14340
rect 35952 14300 36268 14328
rect 35952 14288 35958 14300
rect 36262 14288 36268 14300
rect 36320 14328 36326 14340
rect 37277 14331 37335 14337
rect 37277 14328 37289 14331
rect 36320 14300 37289 14328
rect 36320 14288 36326 14300
rect 37277 14297 37289 14300
rect 37323 14297 37335 14331
rect 39132 14328 39160 14356
rect 40512 14328 40540 14436
rect 41138 14424 41144 14436
rect 41196 14424 41202 14476
rect 41322 14424 41328 14476
rect 41380 14464 41386 14476
rect 50522 14464 50528 14476
rect 41380 14436 50528 14464
rect 41380 14424 41386 14436
rect 50522 14424 50528 14436
rect 50580 14424 50586 14476
rect 40589 14399 40647 14405
rect 40589 14365 40601 14399
rect 40635 14396 40647 14399
rect 40635 14368 41184 14396
rect 40635 14365 40647 14368
rect 40589 14359 40647 14365
rect 37277 14291 37335 14297
rect 37384 14300 40540 14328
rect 41156 14328 41184 14368
rect 41230 14356 41236 14408
rect 41288 14356 41294 14408
rect 45833 14399 45891 14405
rect 45833 14365 45845 14399
rect 45879 14365 45891 14399
rect 45833 14359 45891 14365
rect 42150 14328 42156 14340
rect 41156 14300 42156 14328
rect 37384 14260 37412 14300
rect 42150 14288 42156 14300
rect 42208 14288 42214 14340
rect 45848 14328 45876 14359
rect 43640 14300 45876 14328
rect 35820 14232 37412 14260
rect 38746 14220 38752 14272
rect 38804 14220 38810 14272
rect 38838 14220 38844 14272
rect 38896 14260 38902 14272
rect 39117 14263 39175 14269
rect 39117 14260 39129 14263
rect 38896 14232 39129 14260
rect 38896 14220 38902 14232
rect 39117 14229 39129 14232
rect 39163 14229 39175 14263
rect 39117 14223 39175 14229
rect 40405 14263 40463 14269
rect 40405 14229 40417 14263
rect 40451 14260 40463 14263
rect 40954 14260 40960 14272
rect 40451 14232 40960 14260
rect 40451 14229 40463 14232
rect 40405 14223 40463 14229
rect 40954 14220 40960 14232
rect 41012 14220 41018 14272
rect 41049 14263 41107 14269
rect 41049 14229 41061 14263
rect 41095 14260 41107 14263
rect 43640 14260 43668 14300
rect 41095 14232 43668 14260
rect 41095 14229 41107 14232
rect 41049 14223 41107 14229
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 23750 14056 23756 14068
rect 23532 14028 23756 14056
rect 23532 14016 23538 14028
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 23842 14016 23848 14068
rect 23900 14056 23906 14068
rect 24581 14059 24639 14065
rect 24581 14056 24593 14059
rect 23900 14028 24593 14056
rect 23900 14016 23906 14028
rect 24581 14025 24593 14028
rect 24627 14025 24639 14059
rect 24581 14019 24639 14025
rect 25866 14016 25872 14068
rect 25924 14016 25930 14068
rect 26234 14016 26240 14068
rect 26292 14016 26298 14068
rect 26329 14059 26387 14065
rect 26329 14025 26341 14059
rect 26375 14056 26387 14059
rect 28166 14056 28172 14068
rect 26375 14028 28172 14056
rect 26375 14025 26387 14028
rect 26329 14019 26387 14025
rect 28166 14016 28172 14028
rect 28224 14016 28230 14068
rect 29914 14016 29920 14068
rect 29972 14056 29978 14068
rect 30285 14059 30343 14065
rect 30285 14056 30297 14059
rect 29972 14028 30297 14056
rect 29972 14016 29978 14028
rect 30285 14025 30297 14028
rect 30331 14025 30343 14059
rect 30285 14019 30343 14025
rect 30653 14059 30711 14065
rect 30653 14025 30665 14059
rect 30699 14056 30711 14059
rect 32122 14056 32128 14068
rect 30699 14028 32128 14056
rect 30699 14025 30711 14028
rect 30653 14019 30711 14025
rect 32122 14016 32128 14028
rect 32180 14016 32186 14068
rect 33318 14016 33324 14068
rect 33376 14056 33382 14068
rect 34609 14059 34667 14065
rect 33376 14028 33548 14056
rect 33376 14016 33382 14028
rect 23492 13988 23520 14016
rect 24762 13988 24768 14000
rect 22848 13960 23520 13988
rect 24334 13960 24768 13988
rect 22848 13929 22876 13960
rect 24762 13948 24768 13960
rect 24820 13948 24826 14000
rect 25314 13948 25320 14000
rect 25372 13988 25378 14000
rect 29638 13988 29644 14000
rect 25372 13960 27660 13988
rect 29210 13960 29644 13988
rect 25372 13948 25378 13960
rect 22833 13923 22891 13929
rect 22833 13889 22845 13923
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 27522 13920 27528 13932
rect 26292 13892 27528 13920
rect 26292 13880 26298 13892
rect 27522 13880 27528 13892
rect 27580 13880 27586 13932
rect 27632 13920 27660 13960
rect 29638 13948 29644 13960
rect 29696 13948 29702 14000
rect 33410 13988 33416 14000
rect 31772 13960 33416 13988
rect 27706 13920 27712 13932
rect 27764 13929 27770 13932
rect 31772 13929 31800 13960
rect 33410 13948 33416 13960
rect 33468 13948 33474 14000
rect 33520 13988 33548 14028
rect 34609 14025 34621 14059
rect 34655 14056 34667 14059
rect 34790 14056 34796 14068
rect 34655 14028 34796 14056
rect 34655 14025 34667 14028
rect 34609 14019 34667 14025
rect 34790 14016 34796 14028
rect 34848 14016 34854 14068
rect 35066 14016 35072 14068
rect 35124 14056 35130 14068
rect 37829 14059 37887 14065
rect 37829 14056 37841 14059
rect 35124 14028 37841 14056
rect 35124 14016 35130 14028
rect 37829 14025 37841 14028
rect 37875 14025 37887 14059
rect 37829 14019 37887 14025
rect 37918 14016 37924 14068
rect 37976 14016 37982 14068
rect 38746 14016 38752 14068
rect 38804 14056 38810 14068
rect 42426 14056 42432 14068
rect 38804 14028 42432 14056
rect 38804 14016 38810 14028
rect 42426 14016 42432 14028
rect 42484 14016 42490 14068
rect 43441 14059 43499 14065
rect 43441 14025 43453 14059
rect 43487 14056 43499 14059
rect 44450 14056 44456 14068
rect 43487 14028 44456 14056
rect 43487 14025 43499 14028
rect 43441 14019 43499 14025
rect 44450 14016 44456 14028
rect 44508 14016 44514 14068
rect 33520 13960 33626 13988
rect 34514 13948 34520 14000
rect 34572 13988 34578 14000
rect 35250 13988 35256 14000
rect 34572 13960 35256 13988
rect 34572 13948 34578 13960
rect 35250 13948 35256 13960
rect 35308 13948 35314 14000
rect 37366 13988 37372 14000
rect 35360 13960 37372 13988
rect 27632 13892 27712 13920
rect 27706 13880 27712 13892
rect 27764 13883 27774 13929
rect 30745 13923 30803 13929
rect 30745 13889 30757 13923
rect 30791 13920 30803 13923
rect 31757 13923 31815 13929
rect 30791 13892 31248 13920
rect 30791 13889 30803 13892
rect 30745 13883 30803 13889
rect 27764 13880 27770 13883
rect 26513 13855 26571 13861
rect 22940 13824 24164 13852
rect 20070 13676 20076 13728
rect 20128 13716 20134 13728
rect 20257 13719 20315 13725
rect 20257 13716 20269 13719
rect 20128 13688 20269 13716
rect 20128 13676 20134 13688
rect 20257 13685 20269 13688
rect 20303 13685 20315 13719
rect 20257 13679 20315 13685
rect 20346 13676 20352 13728
rect 20404 13716 20410 13728
rect 22940 13716 22968 13824
rect 24136 13784 24164 13824
rect 26513 13821 26525 13855
rect 26559 13821 26571 13855
rect 26513 13815 26571 13821
rect 26418 13784 26424 13796
rect 24136 13756 26424 13784
rect 26418 13744 26424 13756
rect 26476 13744 26482 13796
rect 26528 13784 26556 13815
rect 28534 13812 28540 13864
rect 28592 13852 28598 13864
rect 28718 13852 28724 13864
rect 28592 13824 28724 13852
rect 28592 13812 28598 13824
rect 28718 13812 28724 13824
rect 28776 13812 28782 13864
rect 30466 13812 30472 13864
rect 30524 13852 30530 13864
rect 30837 13855 30895 13861
rect 30837 13852 30849 13855
rect 30524 13824 30849 13852
rect 30524 13812 30530 13824
rect 30837 13821 30849 13824
rect 30883 13821 30895 13855
rect 31220 13852 31248 13892
rect 31757 13889 31769 13923
rect 31803 13889 31815 13923
rect 31757 13883 31815 13889
rect 32858 13880 32864 13932
rect 32916 13880 32922 13932
rect 35360 13920 35388 13960
rect 37366 13948 37372 13960
rect 37424 13948 37430 14000
rect 39301 13991 39359 13997
rect 39301 13957 39313 13991
rect 39347 13988 39359 13991
rect 39390 13988 39396 14000
rect 39347 13960 39396 13988
rect 39347 13957 39359 13960
rect 39301 13951 39359 13957
rect 39390 13948 39396 13960
rect 39448 13948 39454 14000
rect 42702 13948 42708 14000
rect 42760 13988 42766 14000
rect 45741 13991 45799 13997
rect 45741 13988 45753 13991
rect 42760 13960 45753 13988
rect 42760 13948 42766 13960
rect 45741 13957 45753 13960
rect 45787 13957 45799 13991
rect 45741 13951 45799 13957
rect 35084 13892 35388 13920
rect 35437 13923 35495 13929
rect 32674 13852 32680 13864
rect 31220 13824 32680 13852
rect 30837 13815 30895 13821
rect 32674 13812 32680 13824
rect 32732 13812 32738 13864
rect 27246 13784 27252 13796
rect 26528 13756 27252 13784
rect 27246 13744 27252 13756
rect 27304 13744 27310 13796
rect 32858 13784 32864 13796
rect 32324 13756 32864 13784
rect 20404 13688 22968 13716
rect 23096 13719 23154 13725
rect 20404 13676 20410 13688
rect 23096 13685 23108 13719
rect 23142 13716 23154 13719
rect 23474 13716 23480 13728
rect 23142 13688 23480 13716
rect 23142 13685 23154 13688
rect 23096 13679 23154 13685
rect 23474 13676 23480 13688
rect 23532 13676 23538 13728
rect 24670 13676 24676 13728
rect 24728 13716 24734 13728
rect 26786 13716 26792 13728
rect 24728 13688 26792 13716
rect 24728 13676 24734 13688
rect 26786 13676 26792 13688
rect 26844 13716 26850 13728
rect 27522 13716 27528 13728
rect 26844 13688 27528 13716
rect 26844 13676 26850 13688
rect 27522 13676 27528 13688
rect 27580 13676 27586 13728
rect 27972 13719 28030 13725
rect 27972 13685 27984 13719
rect 28018 13716 28030 13719
rect 28074 13716 28080 13728
rect 28018 13688 28080 13716
rect 28018 13685 28030 13688
rect 27972 13679 28030 13685
rect 28074 13676 28080 13688
rect 28132 13676 28138 13728
rect 28166 13676 28172 13728
rect 28224 13716 28230 13728
rect 28534 13716 28540 13728
rect 28224 13688 28540 13716
rect 28224 13676 28230 13688
rect 28534 13676 28540 13688
rect 28592 13716 28598 13728
rect 29362 13716 29368 13728
rect 28592 13688 29368 13716
rect 28592 13676 28598 13688
rect 29362 13676 29368 13688
rect 29420 13676 29426 13728
rect 29454 13676 29460 13728
rect 29512 13716 29518 13728
rect 32324 13716 32352 13756
rect 32858 13744 32864 13756
rect 32916 13744 32922 13796
rect 35084 13793 35112 13892
rect 35437 13889 35449 13923
rect 35483 13920 35495 13923
rect 36449 13923 36507 13929
rect 36449 13920 36461 13923
rect 35483 13892 36461 13920
rect 35483 13889 35495 13892
rect 35437 13883 35495 13889
rect 36449 13889 36461 13892
rect 36495 13889 36507 13923
rect 36449 13883 36507 13889
rect 37476 13892 38516 13920
rect 35250 13812 35256 13864
rect 35308 13852 35314 13864
rect 35529 13855 35587 13861
rect 35529 13852 35541 13855
rect 35308 13824 35541 13852
rect 35308 13812 35314 13824
rect 35529 13821 35541 13824
rect 35575 13821 35587 13855
rect 35529 13815 35587 13821
rect 35621 13855 35679 13861
rect 35621 13821 35633 13855
rect 35667 13821 35679 13855
rect 35621 13815 35679 13821
rect 35069 13787 35127 13793
rect 35069 13753 35081 13787
rect 35115 13753 35127 13787
rect 35069 13747 35127 13753
rect 29512 13688 32352 13716
rect 29512 13676 29518 13688
rect 32398 13676 32404 13728
rect 32456 13716 32462 13728
rect 33118 13719 33176 13725
rect 33118 13716 33130 13719
rect 32456 13688 33130 13716
rect 32456 13676 32462 13688
rect 33118 13685 33130 13688
rect 33164 13685 33176 13719
rect 35636 13716 35664 13815
rect 37476 13793 37504 13892
rect 38105 13855 38163 13861
rect 38105 13821 38117 13855
rect 38151 13821 38163 13855
rect 38488 13852 38516 13892
rect 38562 13880 38568 13932
rect 38620 13920 38626 13932
rect 39022 13920 39028 13932
rect 38620 13892 39028 13920
rect 38620 13880 38626 13892
rect 39022 13880 39028 13892
rect 39080 13880 39086 13932
rect 40402 13880 40408 13932
rect 40460 13920 40466 13932
rect 40586 13920 40592 13932
rect 40460 13892 40592 13920
rect 40460 13880 40466 13892
rect 40586 13880 40592 13892
rect 40644 13880 40650 13932
rect 43346 13880 43352 13932
rect 43404 13880 43410 13932
rect 47762 13880 47768 13932
rect 47820 13920 47826 13932
rect 47949 13923 48007 13929
rect 47949 13920 47961 13923
rect 47820 13892 47961 13920
rect 47820 13880 47826 13892
rect 47949 13889 47961 13892
rect 47995 13889 48007 13923
rect 47949 13883 48007 13889
rect 40678 13852 40684 13864
rect 38488 13824 40684 13852
rect 38105 13815 38163 13821
rect 37461 13787 37519 13793
rect 37461 13753 37473 13787
rect 37507 13753 37519 13787
rect 38120 13784 38148 13815
rect 40678 13812 40684 13824
rect 40736 13812 40742 13864
rect 45922 13812 45928 13864
rect 45980 13812 45986 13864
rect 49142 13812 49148 13864
rect 49200 13812 49206 13864
rect 38120 13756 38240 13784
rect 37461 13747 37519 13753
rect 37642 13716 37648 13728
rect 35636 13688 37648 13716
rect 33118 13679 33176 13685
rect 37642 13676 37648 13688
rect 37700 13676 37706 13728
rect 38212 13716 38240 13756
rect 40770 13716 40776 13728
rect 38212 13688 40776 13716
rect 40770 13676 40776 13688
rect 40828 13676 40834 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 19705 13515 19763 13521
rect 19705 13481 19717 13515
rect 19751 13512 19763 13515
rect 20346 13512 20352 13524
rect 19751 13484 20352 13512
rect 19751 13481 19763 13484
rect 19705 13475 19763 13481
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 20993 13515 21051 13521
rect 20993 13481 21005 13515
rect 21039 13481 21051 13515
rect 22189 13515 22247 13521
rect 22189 13512 22201 13515
rect 20993 13475 21051 13481
rect 21468 13484 22201 13512
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 20395 13348 20944 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 20070 13268 20076 13320
rect 20128 13268 20134 13320
rect 20165 13243 20223 13249
rect 20165 13240 20177 13243
rect 18616 13212 20177 13240
rect 18616 13184 18644 13212
rect 20165 13209 20177 13212
rect 20211 13209 20223 13243
rect 20165 13203 20223 13209
rect 18598 13132 18604 13184
rect 18656 13132 18662 13184
rect 20916 13172 20944 13348
rect 21008 13240 21036 13475
rect 21468 13388 21496 13484
rect 22189 13481 22201 13484
rect 22235 13481 22247 13515
rect 22189 13475 22247 13481
rect 24946 13472 24952 13524
rect 25004 13472 25010 13524
rect 26326 13472 26332 13524
rect 26384 13512 26390 13524
rect 26605 13515 26663 13521
rect 26605 13512 26617 13515
rect 26384 13484 26617 13512
rect 26384 13472 26390 13484
rect 26605 13481 26617 13484
rect 26651 13481 26663 13515
rect 26605 13475 26663 13481
rect 26786 13472 26792 13524
rect 26844 13512 26850 13524
rect 28442 13512 28448 13524
rect 26844 13484 28448 13512
rect 26844 13472 26850 13484
rect 28442 13472 28448 13484
rect 28500 13472 28506 13524
rect 29638 13472 29644 13524
rect 29696 13512 29702 13524
rect 31018 13512 31024 13524
rect 29696 13484 31024 13512
rect 29696 13472 29702 13484
rect 31018 13472 31024 13484
rect 31076 13472 31082 13524
rect 32306 13512 32312 13524
rect 31588 13484 32312 13512
rect 26418 13444 26424 13456
rect 21652 13416 26424 13444
rect 21450 13336 21456 13388
rect 21508 13336 21514 13388
rect 21652 13385 21680 13416
rect 26418 13404 26424 13416
rect 26476 13404 26482 13456
rect 27522 13404 27528 13456
rect 27580 13444 27586 13456
rect 30006 13444 30012 13456
rect 27580 13416 30012 13444
rect 27580 13404 27586 13416
rect 30006 13404 30012 13416
rect 30064 13444 30070 13456
rect 30064 13416 30972 13444
rect 30064 13404 30070 13416
rect 21637 13379 21695 13385
rect 21637 13345 21649 13379
rect 21683 13345 21695 13379
rect 21637 13339 21695 13345
rect 25498 13336 25504 13388
rect 25556 13376 25562 13388
rect 27157 13379 27215 13385
rect 27157 13376 27169 13379
rect 25556 13348 27169 13376
rect 25556 13336 25562 13348
rect 27157 13345 27169 13348
rect 27203 13345 27215 13379
rect 27157 13339 27215 13345
rect 28074 13336 28080 13388
rect 28132 13376 28138 13388
rect 28813 13379 28871 13385
rect 28813 13376 28825 13379
rect 28132 13348 28825 13376
rect 28132 13336 28138 13348
rect 28813 13345 28825 13348
rect 28859 13376 28871 13379
rect 30374 13376 30380 13388
rect 28859 13348 30380 13376
rect 28859 13345 28871 13348
rect 28813 13339 28871 13345
rect 30374 13336 30380 13348
rect 30432 13336 30438 13388
rect 30834 13336 30840 13388
rect 30892 13336 30898 13388
rect 30944 13385 30972 13416
rect 30929 13379 30987 13385
rect 30929 13345 30941 13379
rect 30975 13345 30987 13379
rect 30929 13339 30987 13345
rect 21361 13311 21419 13317
rect 21361 13277 21373 13311
rect 21407 13308 21419 13311
rect 22557 13311 22615 13317
rect 22557 13308 22569 13311
rect 21407 13280 22569 13308
rect 21407 13277 21419 13280
rect 21361 13271 21419 13277
rect 22557 13277 22569 13280
rect 22603 13277 22615 13311
rect 26786 13308 26792 13320
rect 22557 13271 22615 13277
rect 23216 13280 26792 13308
rect 23216 13240 23244 13280
rect 26786 13268 26792 13280
rect 26844 13268 26850 13320
rect 26878 13268 26884 13320
rect 26936 13308 26942 13320
rect 28537 13311 28595 13317
rect 28537 13308 28549 13311
rect 26936 13280 28549 13308
rect 26936 13268 26942 13280
rect 28537 13277 28549 13280
rect 28583 13277 28595 13311
rect 28537 13271 28595 13277
rect 28629 13311 28687 13317
rect 28629 13277 28641 13311
rect 28675 13308 28687 13311
rect 30650 13308 30656 13320
rect 28675 13280 30656 13308
rect 28675 13277 28687 13280
rect 28629 13271 28687 13277
rect 30650 13268 30656 13280
rect 30708 13268 30714 13320
rect 31588 13317 31616 13484
rect 32306 13472 32312 13484
rect 32364 13472 32370 13524
rect 32769 13515 32827 13521
rect 32769 13481 32781 13515
rect 32815 13512 32827 13515
rect 37090 13512 37096 13524
rect 32815 13484 37096 13512
rect 32815 13481 32827 13484
rect 32769 13475 32827 13481
rect 37090 13472 37096 13484
rect 37148 13472 37154 13524
rect 37182 13472 37188 13524
rect 37240 13512 37246 13524
rect 38197 13515 38255 13521
rect 38197 13512 38209 13515
rect 37240 13484 38209 13512
rect 37240 13472 37246 13484
rect 38197 13481 38209 13484
rect 38243 13481 38255 13515
rect 38197 13475 38255 13481
rect 38654 13472 38660 13524
rect 38712 13512 38718 13524
rect 48774 13512 48780 13524
rect 38712 13484 48780 13512
rect 38712 13472 38718 13484
rect 48774 13472 48780 13484
rect 48832 13472 48838 13524
rect 31757 13447 31815 13453
rect 31757 13413 31769 13447
rect 31803 13444 31815 13447
rect 35618 13444 35624 13456
rect 31803 13416 35624 13444
rect 31803 13413 31815 13416
rect 31757 13407 31815 13413
rect 35618 13404 35624 13416
rect 35676 13404 35682 13456
rect 42245 13447 42303 13453
rect 42245 13413 42257 13447
rect 42291 13444 42303 13447
rect 44634 13444 44640 13456
rect 42291 13416 44640 13444
rect 42291 13413 42303 13416
rect 42245 13407 42303 13413
rect 44634 13404 44640 13416
rect 44692 13404 44698 13456
rect 31680 13348 32352 13376
rect 30745 13311 30803 13317
rect 30745 13277 30757 13311
rect 30791 13308 30803 13311
rect 31573 13311 31631 13317
rect 31573 13308 31585 13311
rect 30791 13280 31585 13308
rect 30791 13277 30803 13280
rect 30745 13271 30803 13277
rect 31573 13277 31585 13280
rect 31619 13277 31631 13311
rect 31573 13271 31631 13277
rect 21008 13212 23244 13240
rect 23290 13200 23296 13252
rect 23348 13240 23354 13252
rect 24854 13240 24860 13252
rect 23348 13212 24860 13240
rect 23348 13200 23354 13212
rect 24854 13200 24860 13212
rect 24912 13200 24918 13252
rect 25317 13243 25375 13249
rect 25317 13209 25329 13243
rect 25363 13240 25375 13243
rect 27798 13240 27804 13252
rect 25363 13212 27804 13240
rect 25363 13209 25375 13212
rect 25317 13203 25375 13209
rect 27798 13200 27804 13212
rect 27856 13200 27862 13252
rect 31680 13240 31708 13348
rect 31754 13268 31760 13320
rect 31812 13308 31818 13320
rect 32125 13311 32183 13317
rect 32125 13308 32137 13311
rect 31812 13280 32137 13308
rect 31812 13268 31818 13280
rect 32125 13277 32137 13280
rect 32171 13277 32183 13311
rect 32125 13271 32183 13277
rect 28184 13212 31708 13240
rect 32324 13240 32352 13348
rect 32398 13336 32404 13388
rect 32456 13336 32462 13388
rect 32858 13336 32864 13388
rect 32916 13376 32922 13388
rect 33321 13379 33379 13385
rect 33321 13376 33333 13379
rect 32916 13348 33333 13376
rect 32916 13336 32922 13348
rect 33321 13345 33333 13348
rect 33367 13345 33379 13379
rect 33321 13339 33379 13345
rect 36262 13336 36268 13388
rect 36320 13376 36326 13388
rect 36449 13379 36507 13385
rect 36449 13376 36461 13379
rect 36320 13348 36461 13376
rect 36320 13336 36326 13348
rect 36449 13345 36461 13348
rect 36495 13376 36507 13379
rect 39022 13376 39028 13388
rect 36495 13348 39028 13376
rect 36495 13345 36507 13348
rect 36449 13339 36507 13345
rect 39022 13336 39028 13348
rect 39080 13336 39086 13388
rect 42334 13376 42340 13388
rect 40236 13348 42340 13376
rect 33137 13311 33195 13317
rect 33137 13277 33149 13311
rect 33183 13308 33195 13311
rect 33410 13308 33416 13320
rect 33183 13280 33416 13308
rect 33183 13277 33195 13280
rect 33137 13271 33195 13277
rect 33410 13268 33416 13280
rect 33468 13268 33474 13320
rect 35158 13308 35164 13320
rect 34440 13280 35164 13308
rect 33229 13243 33287 13249
rect 33229 13240 33241 13243
rect 32324 13212 33241 13240
rect 24026 13172 24032 13184
rect 20916 13144 24032 13172
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 25406 13132 25412 13184
rect 25464 13132 25470 13184
rect 26418 13132 26424 13184
rect 26476 13172 26482 13184
rect 26694 13172 26700 13184
rect 26476 13144 26700 13172
rect 26476 13132 26482 13144
rect 26694 13132 26700 13144
rect 26752 13132 26758 13184
rect 26970 13132 26976 13184
rect 27028 13132 27034 13184
rect 27065 13175 27123 13181
rect 27065 13141 27077 13175
rect 27111 13172 27123 13175
rect 28074 13172 28080 13184
rect 27111 13144 28080 13172
rect 27111 13141 27123 13144
rect 27065 13135 27123 13141
rect 28074 13132 28080 13144
rect 28132 13132 28138 13184
rect 28184 13181 28212 13212
rect 33229 13209 33241 13212
rect 33275 13209 33287 13243
rect 34440 13240 34468 13280
rect 35158 13268 35164 13280
rect 35216 13268 35222 13320
rect 35713 13311 35771 13317
rect 35713 13277 35725 13311
rect 35759 13308 35771 13311
rect 35802 13308 35808 13320
rect 35759 13280 35808 13308
rect 35759 13277 35771 13280
rect 35713 13271 35771 13277
rect 35802 13268 35808 13280
rect 35860 13268 35866 13320
rect 39482 13268 39488 13320
rect 39540 13268 39546 13320
rect 40236 13317 40264 13348
rect 42334 13336 42340 13348
rect 42392 13336 42398 13388
rect 44453 13379 44511 13385
rect 44453 13345 44465 13379
rect 44499 13376 44511 13379
rect 44726 13376 44732 13388
rect 44499 13348 44732 13376
rect 44499 13345 44511 13348
rect 44453 13339 44511 13345
rect 44726 13336 44732 13348
rect 44784 13336 44790 13388
rect 40221 13311 40279 13317
rect 40221 13277 40233 13311
rect 40267 13277 40279 13311
rect 40221 13271 40279 13277
rect 40494 13268 40500 13320
rect 40552 13308 40558 13320
rect 42429 13311 42487 13317
rect 42429 13308 42441 13311
rect 40552 13280 42441 13308
rect 40552 13268 40558 13280
rect 42429 13277 42441 13280
rect 42475 13277 42487 13311
rect 42429 13271 42487 13277
rect 44269 13311 44327 13317
rect 44269 13277 44281 13311
rect 44315 13308 44327 13311
rect 44358 13308 44364 13320
rect 44315 13280 44364 13308
rect 44315 13277 44327 13280
rect 44269 13271 44327 13277
rect 44358 13268 44364 13280
rect 44416 13268 44422 13320
rect 47854 13268 47860 13320
rect 47912 13308 47918 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 47912 13280 47961 13308
rect 47912 13268 47918 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 33229 13203 33287 13209
rect 33704 13212 34468 13240
rect 28169 13175 28227 13181
rect 28169 13141 28181 13175
rect 28215 13141 28227 13175
rect 28169 13135 28227 13141
rect 28258 13132 28264 13184
rect 28316 13172 28322 13184
rect 29638 13172 29644 13184
rect 28316 13144 29644 13172
rect 28316 13132 28322 13144
rect 29638 13132 29644 13144
rect 29696 13132 29702 13184
rect 30374 13132 30380 13184
rect 30432 13132 30438 13184
rect 32217 13175 32275 13181
rect 32217 13141 32229 13175
rect 32263 13172 32275 13175
rect 33704 13172 33732 13212
rect 34882 13200 34888 13252
rect 34940 13240 34946 13252
rect 34977 13243 35035 13249
rect 34977 13240 34989 13243
rect 34940 13212 34989 13240
rect 34940 13200 34946 13212
rect 34977 13209 34989 13212
rect 35023 13209 35035 13243
rect 34977 13203 35035 13209
rect 35897 13243 35955 13249
rect 35897 13209 35909 13243
rect 35943 13240 35955 13243
rect 35986 13240 35992 13252
rect 35943 13212 35992 13240
rect 35943 13209 35955 13212
rect 35897 13203 35955 13209
rect 35986 13200 35992 13212
rect 36044 13200 36050 13252
rect 36725 13243 36783 13249
rect 36725 13209 36737 13243
rect 36771 13209 36783 13243
rect 36725 13203 36783 13209
rect 32263 13144 33732 13172
rect 32263 13141 32275 13144
rect 32217 13135 32275 13141
rect 33778 13132 33784 13184
rect 33836 13172 33842 13184
rect 35069 13175 35127 13181
rect 35069 13172 35081 13175
rect 33836 13144 35081 13172
rect 33836 13132 33842 13144
rect 35069 13141 35081 13144
rect 35115 13141 35127 13175
rect 36740 13172 36768 13203
rect 37274 13200 37280 13252
rect 37332 13200 37338 13252
rect 49142 13200 49148 13252
rect 49200 13200 49206 13252
rect 37734 13172 37740 13184
rect 36740 13144 37740 13172
rect 35069 13135 35127 13141
rect 37734 13132 37740 13144
rect 37792 13132 37798 13184
rect 39206 13132 39212 13184
rect 39264 13172 39270 13184
rect 39301 13175 39359 13181
rect 39301 13172 39313 13175
rect 39264 13144 39313 13172
rect 39264 13132 39270 13144
rect 39301 13141 39313 13144
rect 39347 13141 39359 13175
rect 39301 13135 39359 13141
rect 40037 13175 40095 13181
rect 40037 13141 40049 13175
rect 40083 13172 40095 13175
rect 40494 13172 40500 13184
rect 40083 13144 40500 13172
rect 40083 13141 40095 13144
rect 40037 13135 40095 13141
rect 40494 13132 40500 13144
rect 40552 13132 40558 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 17218 12928 17224 12980
rect 17276 12968 17282 12980
rect 21450 12968 21456 12980
rect 17276 12940 21456 12968
rect 17276 12928 17282 12940
rect 21450 12928 21456 12940
rect 21508 12928 21514 12980
rect 22925 12971 22983 12977
rect 22925 12937 22937 12971
rect 22971 12968 22983 12971
rect 23382 12968 23388 12980
rect 22971 12940 23388 12968
rect 22971 12937 22983 12940
rect 22925 12931 22983 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 25314 12968 25320 12980
rect 24136 12940 25320 12968
rect 23290 12860 23296 12912
rect 23348 12860 23354 12912
rect 24136 12841 24164 12940
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 27338 12928 27344 12980
rect 27396 12968 27402 12980
rect 27433 12971 27491 12977
rect 27433 12968 27445 12971
rect 27396 12940 27445 12968
rect 27396 12928 27402 12940
rect 27433 12937 27445 12940
rect 27479 12937 27491 12971
rect 27433 12931 27491 12937
rect 27801 12971 27859 12977
rect 27801 12937 27813 12971
rect 27847 12968 27859 12971
rect 30374 12968 30380 12980
rect 27847 12940 30380 12968
rect 27847 12937 27859 12940
rect 27801 12931 27859 12937
rect 30374 12928 30380 12940
rect 30432 12928 30438 12980
rect 31570 12968 31576 12980
rect 30484 12940 31576 12968
rect 24854 12860 24860 12912
rect 24912 12860 24918 12912
rect 27893 12903 27951 12909
rect 27893 12869 27905 12903
rect 27939 12900 27951 12903
rect 29086 12900 29092 12912
rect 27939 12872 29092 12900
rect 27939 12869 27951 12872
rect 27893 12863 27951 12869
rect 29086 12860 29092 12872
rect 29144 12860 29150 12912
rect 29181 12903 29239 12909
rect 29181 12869 29193 12903
rect 29227 12900 29239 12903
rect 30484 12900 30512 12940
rect 31570 12928 31576 12940
rect 31628 12928 31634 12980
rect 32766 12928 32772 12980
rect 32824 12928 32830 12980
rect 48590 12968 48596 12980
rect 35268 12940 37504 12968
rect 29227 12872 30512 12900
rect 29227 12869 29239 12872
rect 29181 12863 29239 12869
rect 31018 12860 31024 12912
rect 31076 12860 31082 12912
rect 32306 12860 32312 12912
rect 32364 12900 32370 12912
rect 35268 12900 35296 12940
rect 32364 12872 35296 12900
rect 32364 12860 32370 12872
rect 35342 12860 35348 12912
rect 35400 12860 35406 12912
rect 36081 12903 36139 12909
rect 36081 12869 36093 12903
rect 36127 12900 36139 12903
rect 36814 12900 36820 12912
rect 36127 12872 36820 12900
rect 36127 12869 36139 12872
rect 36081 12863 36139 12869
rect 36814 12860 36820 12872
rect 36872 12860 36878 12912
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 27246 12792 27252 12844
rect 27304 12832 27310 12844
rect 29273 12835 29331 12841
rect 27304 12804 28028 12832
rect 27304 12792 27310 12804
rect 23385 12767 23443 12773
rect 23385 12733 23397 12767
rect 23431 12733 23443 12767
rect 23385 12727 23443 12733
rect 23400 12696 23428 12727
rect 23474 12724 23480 12776
rect 23532 12724 23538 12776
rect 24397 12767 24455 12773
rect 24397 12733 24409 12767
rect 24443 12764 24455 12767
rect 24762 12764 24768 12776
rect 24443 12736 24768 12764
rect 24443 12733 24455 12736
rect 24397 12727 24455 12733
rect 24762 12724 24768 12736
rect 24820 12724 24826 12776
rect 24854 12724 24860 12776
rect 24912 12764 24918 12776
rect 25130 12764 25136 12776
rect 24912 12736 25136 12764
rect 24912 12724 24918 12736
rect 25130 12724 25136 12736
rect 25188 12724 25194 12776
rect 26694 12724 26700 12776
rect 26752 12764 26758 12776
rect 27890 12764 27896 12776
rect 26752 12736 27896 12764
rect 26752 12724 26758 12736
rect 27890 12724 27896 12736
rect 27948 12724 27954 12776
rect 28000 12773 28028 12804
rect 29273 12801 29285 12835
rect 29319 12832 29331 12835
rect 29914 12832 29920 12844
rect 29319 12804 29920 12832
rect 29319 12801 29331 12804
rect 29273 12795 29331 12801
rect 29914 12792 29920 12804
rect 29972 12792 29978 12844
rect 32677 12835 32735 12841
rect 32677 12832 32689 12835
rect 31726 12804 32689 12832
rect 27985 12767 28043 12773
rect 27985 12733 27997 12767
rect 28031 12733 28043 12767
rect 27985 12727 28043 12733
rect 28074 12724 28080 12776
rect 28132 12764 28138 12776
rect 28132 12736 29316 12764
rect 28132 12724 28138 12736
rect 26602 12696 26608 12708
rect 23400 12668 23520 12696
rect 23492 12628 23520 12668
rect 25424 12668 26608 12696
rect 25424 12628 25452 12668
rect 26602 12656 26608 12668
rect 26660 12656 26666 12708
rect 26970 12656 26976 12708
rect 27028 12696 27034 12708
rect 28813 12699 28871 12705
rect 28813 12696 28825 12699
rect 27028 12668 28825 12696
rect 27028 12656 27034 12668
rect 28813 12665 28825 12668
rect 28859 12665 28871 12699
rect 29288 12696 29316 12736
rect 29362 12724 29368 12776
rect 29420 12724 29426 12776
rect 29730 12724 29736 12776
rect 29788 12764 29794 12776
rect 30009 12767 30067 12773
rect 30009 12764 30021 12767
rect 29788 12736 30021 12764
rect 29788 12724 29794 12736
rect 30009 12733 30021 12736
rect 30055 12733 30067 12767
rect 30285 12767 30343 12773
rect 30285 12764 30297 12767
rect 30009 12727 30067 12733
rect 30116 12736 30297 12764
rect 30116 12696 30144 12736
rect 30285 12733 30297 12736
rect 30331 12733 30343 12767
rect 30285 12727 30343 12733
rect 30374 12724 30380 12776
rect 30432 12764 30438 12776
rect 31726 12764 31754 12804
rect 32677 12801 32689 12804
rect 32723 12801 32735 12835
rect 34054 12832 34060 12844
rect 32677 12795 32735 12801
rect 32968 12804 34060 12832
rect 32968 12773 32996 12804
rect 34054 12792 34060 12804
rect 34112 12792 34118 12844
rect 36909 12835 36967 12841
rect 36909 12801 36921 12835
rect 36955 12801 36967 12835
rect 37476 12832 37504 12940
rect 37568 12940 48596 12968
rect 37568 12909 37596 12940
rect 48590 12928 48596 12940
rect 48648 12928 48654 12980
rect 37553 12903 37611 12909
rect 37553 12869 37565 12903
rect 37599 12869 37611 12903
rect 37553 12863 37611 12869
rect 38654 12832 38660 12844
rect 37476 12804 38660 12832
rect 36909 12795 36967 12801
rect 30432 12736 31754 12764
rect 32953 12767 33011 12773
rect 30432 12724 30438 12736
rect 32953 12733 32965 12767
rect 32999 12733 33011 12767
rect 32953 12727 33011 12733
rect 33962 12724 33968 12776
rect 34020 12764 34026 12776
rect 35529 12767 35587 12773
rect 35529 12764 35541 12767
rect 34020 12736 35541 12764
rect 34020 12724 34026 12736
rect 35529 12733 35541 12736
rect 35575 12733 35587 12767
rect 35529 12727 35587 12733
rect 33870 12696 33876 12708
rect 29288 12668 30144 12696
rect 28813 12659 28871 12665
rect 23492 12600 25452 12628
rect 25498 12588 25504 12640
rect 25556 12628 25562 12640
rect 25869 12631 25927 12637
rect 25869 12628 25881 12631
rect 25556 12600 25881 12628
rect 25556 12588 25562 12600
rect 25869 12597 25881 12600
rect 25915 12597 25927 12631
rect 25869 12591 25927 12597
rect 27798 12588 27804 12640
rect 27856 12628 27862 12640
rect 28350 12628 28356 12640
rect 27856 12600 28356 12628
rect 27856 12588 27862 12600
rect 28350 12588 28356 12600
rect 28408 12588 28414 12640
rect 28626 12588 28632 12640
rect 28684 12628 28690 12640
rect 28994 12628 29000 12640
rect 28684 12600 29000 12628
rect 28684 12588 28690 12600
rect 28994 12588 29000 12600
rect 29052 12588 29058 12640
rect 30116 12628 30144 12668
rect 31312 12668 33876 12696
rect 31312 12628 31340 12668
rect 33870 12656 33876 12668
rect 33928 12656 33934 12708
rect 34698 12656 34704 12708
rect 34756 12696 34762 12708
rect 34756 12668 34928 12696
rect 34756 12656 34762 12668
rect 30116 12600 31340 12628
rect 31754 12588 31760 12640
rect 31812 12588 31818 12640
rect 32306 12588 32312 12640
rect 32364 12588 32370 12640
rect 33686 12588 33692 12640
rect 33744 12588 33750 12640
rect 34790 12588 34796 12640
rect 34848 12588 34854 12640
rect 34900 12628 34928 12668
rect 34974 12656 34980 12708
rect 35032 12696 35038 12708
rect 36265 12699 36323 12705
rect 36265 12696 36277 12699
rect 35032 12668 36277 12696
rect 35032 12656 35038 12668
rect 36265 12665 36277 12668
rect 36311 12665 36323 12699
rect 36924 12696 36952 12795
rect 38654 12792 38660 12804
rect 38712 12792 38718 12844
rect 39022 12792 39028 12844
rect 39080 12832 39086 12844
rect 39209 12835 39267 12841
rect 39209 12832 39221 12835
rect 39080 12804 39221 12832
rect 39080 12792 39086 12804
rect 39209 12801 39221 12804
rect 39255 12801 39267 12835
rect 39209 12795 39267 12801
rect 40586 12792 40592 12844
rect 40644 12792 40650 12844
rect 40862 12792 40868 12844
rect 40920 12832 40926 12844
rect 41693 12835 41751 12841
rect 41693 12832 41705 12835
rect 40920 12804 41705 12832
rect 40920 12792 40926 12804
rect 41693 12801 41705 12804
rect 41739 12801 41751 12835
rect 41693 12795 41751 12801
rect 39485 12767 39543 12773
rect 39485 12733 39497 12767
rect 39531 12764 39543 12767
rect 40770 12764 40776 12776
rect 39531 12736 40776 12764
rect 39531 12733 39543 12736
rect 39485 12727 39543 12733
rect 40770 12724 40776 12736
rect 40828 12724 40834 12776
rect 36924 12668 39344 12696
rect 36265 12659 36323 12665
rect 36725 12631 36783 12637
rect 36725 12628 36737 12631
rect 34900 12600 36737 12628
rect 36725 12597 36737 12600
rect 36771 12597 36783 12631
rect 36725 12591 36783 12597
rect 37642 12588 37648 12640
rect 37700 12588 37706 12640
rect 39316 12628 39344 12668
rect 40218 12628 40224 12640
rect 39316 12600 40224 12628
rect 40218 12588 40224 12600
rect 40276 12588 40282 12640
rect 40678 12588 40684 12640
rect 40736 12628 40742 12640
rect 40957 12631 41015 12637
rect 40957 12628 40969 12631
rect 40736 12600 40969 12628
rect 40736 12588 40742 12600
rect 40957 12597 40969 12600
rect 41003 12597 41015 12631
rect 40957 12591 41015 12597
rect 41509 12631 41567 12637
rect 41509 12597 41521 12631
rect 41555 12628 41567 12631
rect 44174 12628 44180 12640
rect 41555 12600 44180 12628
rect 41555 12597 41567 12600
rect 41509 12591 41567 12597
rect 44174 12588 44180 12600
rect 44232 12588 44238 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 24581 12427 24639 12433
rect 24581 12393 24593 12427
rect 24627 12424 24639 12427
rect 25406 12424 25412 12436
rect 24627 12396 25412 12424
rect 24627 12393 24639 12396
rect 24581 12387 24639 12393
rect 25406 12384 25412 12396
rect 25464 12384 25470 12436
rect 27062 12384 27068 12436
rect 27120 12424 27126 12436
rect 27249 12427 27307 12433
rect 27249 12424 27261 12427
rect 27120 12396 27261 12424
rect 27120 12384 27126 12396
rect 27249 12393 27261 12396
rect 27295 12393 27307 12427
rect 27249 12387 27307 12393
rect 27540 12396 27752 12424
rect 24762 12316 24768 12368
rect 24820 12356 24826 12368
rect 24820 12328 25176 12356
rect 24820 12316 24826 12328
rect 25038 12248 25044 12300
rect 25096 12248 25102 12300
rect 25148 12297 25176 12328
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12257 25191 12291
rect 25133 12251 25191 12257
rect 24578 12180 24584 12232
rect 24636 12220 24642 12232
rect 26697 12223 26755 12229
rect 26697 12220 26709 12223
rect 24636 12192 26709 12220
rect 24636 12180 24642 12192
rect 26697 12189 26709 12192
rect 26743 12220 26755 12223
rect 27540 12220 27568 12396
rect 27614 12316 27620 12368
rect 27672 12316 27678 12368
rect 27724 12356 27752 12396
rect 29546 12384 29552 12436
rect 29604 12424 29610 12436
rect 29733 12427 29791 12433
rect 29733 12424 29745 12427
rect 29604 12396 29745 12424
rect 29604 12384 29610 12396
rect 29733 12393 29745 12396
rect 29779 12393 29791 12427
rect 29733 12387 29791 12393
rect 31846 12384 31852 12436
rect 31904 12424 31910 12436
rect 32490 12424 32496 12436
rect 31904 12396 32496 12424
rect 31904 12384 31910 12396
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 33137 12427 33195 12433
rect 33137 12393 33149 12427
rect 33183 12424 33195 12427
rect 33502 12424 33508 12436
rect 33183 12396 33508 12424
rect 33183 12393 33195 12396
rect 33137 12387 33195 12393
rect 33502 12384 33508 12396
rect 33560 12384 33566 12436
rect 36170 12424 36176 12436
rect 33796 12396 36176 12424
rect 28166 12356 28172 12368
rect 27724 12328 28172 12356
rect 27632 12229 27660 12316
rect 27724 12229 27752 12328
rect 28166 12316 28172 12328
rect 28224 12316 28230 12368
rect 28718 12316 28724 12368
rect 28776 12316 28782 12368
rect 31754 12356 31760 12368
rect 31726 12316 31760 12356
rect 31812 12316 31818 12368
rect 31941 12359 31999 12365
rect 31941 12325 31953 12359
rect 31987 12325 31999 12359
rect 31941 12319 31999 12325
rect 27893 12291 27951 12297
rect 27893 12257 27905 12291
rect 27939 12288 27951 12291
rect 28442 12288 28448 12300
rect 27939 12260 28448 12288
rect 27939 12257 27951 12260
rect 27893 12251 27951 12257
rect 28442 12248 28448 12260
rect 28500 12288 28506 12300
rect 28736 12288 28764 12316
rect 30282 12288 30288 12300
rect 28500 12260 30288 12288
rect 28500 12248 28506 12260
rect 30282 12248 30288 12260
rect 30340 12248 30346 12300
rect 26743 12192 27568 12220
rect 27617 12223 27675 12229
rect 26743 12189 26755 12192
rect 26697 12183 26755 12189
rect 27617 12189 27629 12223
rect 27663 12189 27675 12223
rect 27617 12183 27675 12189
rect 27709 12223 27767 12229
rect 27709 12189 27721 12223
rect 27755 12189 27767 12223
rect 27709 12183 27767 12189
rect 28629 12223 28687 12229
rect 28629 12189 28641 12223
rect 28675 12220 28687 12223
rect 28718 12220 28724 12232
rect 28675 12192 28724 12220
rect 28675 12189 28687 12192
rect 28629 12183 28687 12189
rect 28718 12180 28724 12192
rect 28776 12180 28782 12232
rect 30098 12180 30104 12232
rect 30156 12220 30162 12232
rect 31726 12220 31754 12316
rect 30156 12192 31754 12220
rect 31956 12220 31984 12319
rect 32214 12248 32220 12300
rect 32272 12288 32278 12300
rect 32401 12291 32459 12297
rect 32401 12288 32413 12291
rect 32272 12260 32413 12288
rect 32272 12248 32278 12260
rect 32401 12257 32413 12260
rect 32447 12257 32459 12291
rect 32401 12251 32459 12257
rect 32490 12248 32496 12300
rect 32548 12248 32554 12300
rect 33796 12297 33824 12396
rect 36170 12384 36176 12396
rect 36228 12424 36234 12436
rect 37182 12424 37188 12436
rect 36228 12396 37188 12424
rect 36228 12384 36234 12396
rect 37182 12384 37188 12396
rect 37240 12384 37246 12436
rect 37734 12384 37740 12436
rect 37792 12424 37798 12436
rect 38013 12427 38071 12433
rect 38013 12424 38025 12427
rect 37792 12396 38025 12424
rect 37792 12384 37798 12396
rect 38013 12393 38025 12396
rect 38059 12393 38071 12427
rect 38013 12387 38071 12393
rect 35452 12328 36400 12356
rect 33781 12291 33839 12297
rect 33781 12257 33793 12291
rect 33827 12257 33839 12291
rect 33781 12251 33839 12257
rect 35158 12248 35164 12300
rect 35216 12288 35222 12300
rect 35345 12291 35403 12297
rect 35345 12288 35357 12291
rect 35216 12260 35357 12288
rect 35216 12248 35222 12260
rect 35345 12257 35357 12260
rect 35391 12257 35403 12291
rect 35345 12251 35403 12257
rect 35452 12220 35480 12328
rect 35529 12291 35587 12297
rect 35529 12257 35541 12291
rect 35575 12257 35587 12291
rect 35529 12251 35587 12257
rect 31956 12192 35480 12220
rect 30156 12180 30162 12192
rect 28258 12152 28264 12164
rect 24964 12124 28264 12152
rect 24964 12096 24992 12124
rect 28258 12112 28264 12124
rect 28316 12112 28322 12164
rect 32309 12155 32367 12161
rect 32309 12152 32321 12155
rect 28368 12124 32321 12152
rect 24946 12044 24952 12096
rect 25004 12044 25010 12096
rect 26142 12044 26148 12096
rect 26200 12084 26206 12096
rect 28368 12084 28396 12124
rect 32309 12121 32321 12124
rect 32355 12121 32367 12155
rect 32309 12115 32367 12121
rect 33505 12155 33563 12161
rect 33505 12121 33517 12155
rect 33551 12152 33563 12155
rect 33686 12152 33692 12164
rect 33551 12124 33692 12152
rect 33551 12121 33563 12124
rect 33505 12115 33563 12121
rect 33686 12112 33692 12124
rect 33744 12112 33750 12164
rect 33870 12112 33876 12164
rect 33928 12152 33934 12164
rect 35253 12155 35311 12161
rect 35253 12152 35265 12155
rect 33928 12124 35265 12152
rect 33928 12112 33934 12124
rect 35253 12121 35265 12124
rect 35299 12121 35311 12155
rect 35544 12152 35572 12251
rect 36262 12248 36268 12300
rect 36320 12248 36326 12300
rect 36372 12288 36400 12328
rect 36372 12260 38700 12288
rect 38672 12229 38700 12260
rect 38657 12223 38715 12229
rect 38657 12189 38669 12223
rect 38703 12189 38715 12223
rect 38657 12183 38715 12189
rect 39298 12180 39304 12232
rect 39356 12180 39362 12232
rect 40221 12223 40279 12229
rect 40221 12189 40233 12223
rect 40267 12220 40279 12223
rect 41046 12220 41052 12232
rect 40267 12192 41052 12220
rect 40267 12189 40279 12192
rect 40221 12183 40279 12189
rect 41046 12180 41052 12192
rect 41104 12180 41110 12232
rect 45922 12180 45928 12232
rect 45980 12220 45986 12232
rect 47949 12223 48007 12229
rect 47949 12220 47961 12223
rect 45980 12192 47961 12220
rect 45980 12180 45986 12192
rect 47949 12189 47961 12192
rect 47995 12189 48007 12223
rect 47949 12183 48007 12189
rect 49142 12180 49148 12232
rect 49200 12180 49206 12232
rect 36541 12155 36599 12161
rect 36541 12152 36553 12155
rect 35544 12124 36553 12152
rect 35253 12115 35311 12121
rect 36541 12121 36553 12124
rect 36587 12152 36599 12155
rect 36630 12152 36636 12164
rect 36587 12124 36636 12152
rect 36587 12121 36599 12124
rect 36541 12115 36599 12121
rect 36630 12112 36636 12124
rect 36688 12112 36694 12164
rect 37274 12112 37280 12164
rect 37332 12112 37338 12164
rect 37826 12112 37832 12164
rect 37884 12152 37890 12164
rect 43346 12152 43352 12164
rect 37884 12124 43352 12152
rect 37884 12112 37890 12124
rect 43346 12112 43352 12124
rect 43404 12112 43410 12164
rect 26200 12056 28396 12084
rect 26200 12044 26206 12056
rect 30190 12044 30196 12096
rect 30248 12044 30254 12096
rect 30374 12044 30380 12096
rect 30432 12084 30438 12096
rect 30650 12084 30656 12096
rect 30432 12056 30656 12084
rect 30432 12044 30438 12056
rect 30650 12044 30656 12056
rect 30708 12044 30714 12096
rect 31110 12044 31116 12096
rect 31168 12084 31174 12096
rect 33597 12087 33655 12093
rect 33597 12084 33609 12087
rect 31168 12056 33609 12084
rect 31168 12044 31174 12056
rect 33597 12053 33609 12056
rect 33643 12053 33655 12087
rect 33597 12047 33655 12053
rect 34885 12087 34943 12093
rect 34885 12053 34897 12087
rect 34931 12084 34943 12087
rect 38286 12084 38292 12096
rect 34931 12056 38292 12084
rect 34931 12053 34943 12056
rect 34885 12047 34943 12053
rect 38286 12044 38292 12056
rect 38344 12044 38350 12096
rect 38470 12044 38476 12096
rect 38528 12044 38534 12096
rect 40037 12087 40095 12093
rect 40037 12053 40049 12087
rect 40083 12084 40095 12087
rect 40862 12084 40868 12096
rect 40083 12056 40868 12084
rect 40083 12053 40095 12056
rect 40037 12047 40095 12053
rect 40862 12044 40868 12056
rect 40920 12044 40926 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 23474 11840 23480 11892
rect 23532 11880 23538 11892
rect 25501 11883 25559 11889
rect 25501 11880 25513 11883
rect 23532 11852 25513 11880
rect 23532 11840 23538 11852
rect 25501 11849 25513 11852
rect 25547 11849 25559 11883
rect 25501 11843 25559 11849
rect 25516 11812 25544 11843
rect 26510 11840 26516 11892
rect 26568 11880 26574 11892
rect 27157 11883 27215 11889
rect 27157 11880 27169 11883
rect 26568 11852 27169 11880
rect 26568 11840 26574 11852
rect 27157 11849 27169 11852
rect 27203 11849 27215 11883
rect 27157 11843 27215 11849
rect 28350 11840 28356 11892
rect 28408 11840 28414 11892
rect 28718 11840 28724 11892
rect 28776 11840 28782 11892
rect 29822 11840 29828 11892
rect 29880 11880 29886 11892
rect 29917 11883 29975 11889
rect 29917 11880 29929 11883
rect 29880 11852 29929 11880
rect 29880 11840 29886 11852
rect 29917 11849 29929 11852
rect 29963 11849 29975 11883
rect 29917 11843 29975 11849
rect 30208 11852 30604 11880
rect 27246 11812 27252 11824
rect 25516 11784 27252 11812
rect 27246 11772 27252 11784
rect 27304 11772 27310 11824
rect 27525 11815 27583 11821
rect 27525 11781 27537 11815
rect 27571 11812 27583 11815
rect 29546 11812 29552 11824
rect 27571 11784 29552 11812
rect 27571 11781 27583 11784
rect 27525 11775 27583 11781
rect 29546 11772 29552 11784
rect 29604 11772 29610 11824
rect 30208 11812 30236 11852
rect 29748 11784 30236 11812
rect 25130 11704 25136 11756
rect 25188 11744 25194 11756
rect 26602 11744 26608 11756
rect 25188 11716 26608 11744
rect 25188 11704 25194 11716
rect 26602 11704 26608 11716
rect 26660 11704 26666 11756
rect 23750 11636 23756 11688
rect 23808 11636 23814 11688
rect 24026 11636 24032 11688
rect 24084 11676 24090 11688
rect 24670 11676 24676 11688
rect 24084 11648 24676 11676
rect 24084 11636 24090 11648
rect 24670 11636 24676 11648
rect 24728 11636 24734 11688
rect 27264 11676 27292 11772
rect 27617 11747 27675 11753
rect 27617 11713 27629 11747
rect 27663 11744 27675 11747
rect 29270 11744 29276 11756
rect 27663 11716 29276 11744
rect 27663 11713 27675 11716
rect 27617 11707 27675 11713
rect 29270 11704 29276 11716
rect 29328 11704 29334 11756
rect 27709 11679 27767 11685
rect 27709 11676 27721 11679
rect 27264 11648 27721 11676
rect 27709 11645 27721 11648
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 28813 11679 28871 11685
rect 28813 11645 28825 11679
rect 28859 11645 28871 11679
rect 28813 11639 28871 11645
rect 28997 11679 29055 11685
rect 28997 11645 29009 11679
rect 29043 11676 29055 11679
rect 29086 11676 29092 11688
rect 29043 11648 29092 11676
rect 29043 11645 29055 11648
rect 28997 11639 29055 11645
rect 23768 11540 23796 11636
rect 28828 11608 28856 11639
rect 29086 11636 29092 11648
rect 29144 11676 29150 11688
rect 29362 11676 29368 11688
rect 29144 11648 29368 11676
rect 29144 11636 29150 11648
rect 29362 11636 29368 11648
rect 29420 11636 29426 11688
rect 29178 11608 29184 11620
rect 28828 11580 29184 11608
rect 29178 11568 29184 11580
rect 29236 11608 29242 11620
rect 29748 11608 29776 11784
rect 30374 11772 30380 11824
rect 30432 11772 30438 11824
rect 30576 11812 30604 11852
rect 31662 11840 31668 11892
rect 31720 11880 31726 11892
rect 33870 11880 33876 11892
rect 31720 11852 33876 11880
rect 31720 11840 31726 11852
rect 33870 11840 33876 11852
rect 33928 11840 33934 11892
rect 34790 11840 34796 11892
rect 34848 11880 34854 11892
rect 35253 11883 35311 11889
rect 35253 11880 35265 11883
rect 34848 11852 35265 11880
rect 34848 11840 34854 11852
rect 35253 11849 35265 11852
rect 35299 11849 35311 11883
rect 35253 11843 35311 11849
rect 36081 11883 36139 11889
rect 36081 11849 36093 11883
rect 36127 11880 36139 11883
rect 37826 11880 37832 11892
rect 36127 11852 37832 11880
rect 36127 11849 36139 11852
rect 36081 11843 36139 11849
rect 37826 11840 37832 11852
rect 37884 11840 37890 11892
rect 38197 11883 38255 11889
rect 38197 11849 38209 11883
rect 38243 11880 38255 11883
rect 39298 11880 39304 11892
rect 38243 11852 39304 11880
rect 38243 11849 38255 11852
rect 38197 11843 38255 11849
rect 39298 11840 39304 11852
rect 39356 11840 39362 11892
rect 40586 11840 40592 11892
rect 40644 11840 40650 11892
rect 34698 11812 34704 11824
rect 30576 11784 34704 11812
rect 34698 11772 34704 11784
rect 34756 11772 34762 11824
rect 36814 11812 36820 11824
rect 34808 11784 36820 11812
rect 30282 11704 30288 11756
rect 30340 11704 30346 11756
rect 30392 11744 30420 11772
rect 30392 11716 30604 11744
rect 30374 11636 30380 11688
rect 30432 11676 30438 11688
rect 30576 11685 30604 11716
rect 31754 11704 31760 11756
rect 31812 11744 31818 11756
rect 34808 11744 34836 11784
rect 36814 11772 36820 11784
rect 36872 11772 36878 11824
rect 38286 11772 38292 11824
rect 38344 11772 38350 11824
rect 38470 11772 38476 11824
rect 38528 11812 38534 11824
rect 38528 11784 44772 11812
rect 38528 11772 38534 11784
rect 31812 11716 34836 11744
rect 35452 11716 36216 11744
rect 31812 11704 31818 11716
rect 30561 11679 30619 11685
rect 30432 11648 30512 11676
rect 30432 11636 30438 11648
rect 29236 11580 29776 11608
rect 30484 11608 30512 11648
rect 30561 11645 30573 11679
rect 30607 11645 30619 11679
rect 30561 11639 30619 11645
rect 33502 11636 33508 11688
rect 33560 11676 33566 11688
rect 35345 11679 35403 11685
rect 35345 11676 35357 11679
rect 33560 11648 35357 11676
rect 33560 11636 33566 11648
rect 35345 11645 35357 11648
rect 35391 11645 35403 11679
rect 35345 11639 35403 11645
rect 35250 11608 35256 11620
rect 30484 11580 35256 11608
rect 29236 11568 29242 11580
rect 35250 11568 35256 11580
rect 35308 11568 35314 11620
rect 24762 11540 24768 11552
rect 23768 11512 24768 11540
rect 24762 11500 24768 11512
rect 24820 11500 24826 11552
rect 27614 11500 27620 11552
rect 27672 11540 27678 11552
rect 32490 11540 32496 11552
rect 27672 11512 32496 11540
rect 27672 11500 27678 11512
rect 32490 11500 32496 11512
rect 32548 11500 32554 11552
rect 34885 11543 34943 11549
rect 34885 11509 34897 11543
rect 34931 11540 34943 11543
rect 35452 11540 35480 11716
rect 35529 11679 35587 11685
rect 35529 11645 35541 11679
rect 35575 11645 35587 11679
rect 36188 11676 36216 11716
rect 36262 11704 36268 11756
rect 36320 11704 36326 11756
rect 37734 11704 37740 11756
rect 37792 11744 37798 11756
rect 37792 11716 38516 11744
rect 37792 11704 37798 11716
rect 37918 11676 37924 11688
rect 36188 11648 37924 11676
rect 35529 11639 35587 11645
rect 34931 11512 35480 11540
rect 35544 11540 35572 11639
rect 37918 11636 37924 11648
rect 37976 11636 37982 11688
rect 38488 11685 38516 11716
rect 38562 11704 38568 11756
rect 38620 11744 38626 11756
rect 38620 11716 38976 11744
rect 38620 11704 38626 11716
rect 38473 11679 38531 11685
rect 38473 11645 38485 11679
rect 38519 11645 38531 11679
rect 38948 11676 38976 11716
rect 39114 11704 39120 11756
rect 39172 11704 39178 11756
rect 40497 11747 40555 11753
rect 40497 11713 40509 11747
rect 40543 11744 40555 11747
rect 41509 11747 41567 11753
rect 41509 11744 41521 11747
rect 40543 11716 41521 11744
rect 40543 11713 40555 11716
rect 40497 11707 40555 11713
rect 41509 11713 41521 11716
rect 41555 11713 41567 11747
rect 41509 11707 41567 11713
rect 42426 11704 42432 11756
rect 42484 11744 42490 11756
rect 44744 11753 44772 11784
rect 42797 11747 42855 11753
rect 42797 11744 42809 11747
rect 42484 11716 42809 11744
rect 42484 11704 42490 11716
rect 42797 11713 42809 11716
rect 42843 11713 42855 11747
rect 42797 11707 42855 11713
rect 44729 11747 44787 11753
rect 44729 11713 44741 11747
rect 44775 11713 44787 11747
rect 44729 11707 44787 11713
rect 47949 11747 48007 11753
rect 47949 11713 47961 11747
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 39301 11679 39359 11685
rect 39301 11676 39313 11679
rect 38948 11648 39313 11676
rect 38473 11639 38531 11645
rect 39301 11645 39313 11648
rect 39347 11645 39359 11679
rect 39301 11639 39359 11645
rect 40678 11636 40684 11688
rect 40736 11636 40742 11688
rect 43714 11676 43720 11688
rect 41386 11648 43720 11676
rect 37829 11611 37887 11617
rect 37829 11577 37841 11611
rect 37875 11608 37887 11611
rect 40129 11611 40187 11617
rect 37875 11580 39620 11608
rect 37875 11577 37887 11580
rect 37829 11571 37887 11577
rect 38930 11540 38936 11552
rect 35544 11512 38936 11540
rect 34931 11509 34943 11512
rect 34885 11503 34943 11509
rect 38930 11500 38936 11512
rect 38988 11500 38994 11552
rect 39592 11540 39620 11580
rect 40129 11577 40141 11611
rect 40175 11608 40187 11611
rect 41386 11608 41414 11648
rect 43714 11636 43720 11648
rect 43772 11636 43778 11688
rect 42794 11608 42800 11620
rect 40175 11580 41414 11608
rect 42076 11580 42800 11608
rect 40175 11577 40187 11580
rect 40129 11571 40187 11577
rect 42076 11540 42104 11580
rect 42794 11568 42800 11580
rect 42852 11568 42858 11620
rect 44545 11611 44603 11617
rect 44545 11577 44557 11611
rect 44591 11608 44603 11611
rect 47964 11608 47992 11707
rect 49142 11636 49148 11688
rect 49200 11636 49206 11688
rect 44591 11580 47992 11608
rect 44591 11577 44603 11580
rect 44545 11571 44603 11577
rect 39592 11512 42104 11540
rect 42613 11543 42671 11549
rect 42613 11509 42625 11543
rect 42659 11540 42671 11543
rect 45186 11540 45192 11552
rect 42659 11512 45192 11540
rect 42659 11509 42671 11512
rect 42613 11503 42671 11509
rect 45186 11500 45192 11512
rect 45244 11500 45250 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 24578 11336 24584 11348
rect 13412 11308 24584 11336
rect 13412 11296 13418 11308
rect 24578 11296 24584 11308
rect 24636 11296 24642 11348
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 27065 11339 27123 11345
rect 27065 11336 27077 11339
rect 24912 11308 27077 11336
rect 24912 11296 24918 11308
rect 27065 11305 27077 11308
rect 27111 11305 27123 11339
rect 27065 11299 27123 11305
rect 28169 11339 28227 11345
rect 28169 11305 28181 11339
rect 28215 11336 28227 11339
rect 28810 11336 28816 11348
rect 28215 11308 28816 11336
rect 28215 11305 28227 11308
rect 28169 11299 28227 11305
rect 19978 11228 19984 11280
rect 20036 11268 20042 11280
rect 27080 11268 27108 11299
rect 28810 11296 28816 11308
rect 28868 11296 28874 11348
rect 29638 11296 29644 11348
rect 29696 11336 29702 11348
rect 29733 11339 29791 11345
rect 29733 11336 29745 11339
rect 29696 11308 29745 11336
rect 29696 11296 29702 11308
rect 29733 11305 29745 11308
rect 29779 11305 29791 11339
rect 29733 11299 29791 11305
rect 29914 11296 29920 11348
rect 29972 11336 29978 11348
rect 30929 11339 30987 11345
rect 30929 11336 30941 11339
rect 29972 11308 30941 11336
rect 29972 11296 29978 11308
rect 30929 11305 30941 11308
rect 30975 11305 30987 11339
rect 30929 11299 30987 11305
rect 32122 11296 32128 11348
rect 32180 11296 32186 11348
rect 37645 11339 37703 11345
rect 32324 11308 37504 11336
rect 32324 11280 32352 11308
rect 29086 11268 29092 11280
rect 20036 11240 22094 11268
rect 27080 11240 29092 11268
rect 20036 11228 20042 11240
rect 22066 11064 22094 11240
rect 29086 11228 29092 11240
rect 29144 11268 29150 11280
rect 29144 11240 30328 11268
rect 29144 11228 29150 11240
rect 25314 11160 25320 11212
rect 25372 11160 25378 11212
rect 25593 11203 25651 11209
rect 25593 11169 25605 11203
rect 25639 11200 25651 11203
rect 26234 11200 26240 11212
rect 25639 11172 26240 11200
rect 25639 11169 25651 11172
rect 25593 11163 25651 11169
rect 26234 11160 26240 11172
rect 26292 11160 26298 11212
rect 28626 11160 28632 11212
rect 28684 11200 28690 11212
rect 28721 11203 28779 11209
rect 28721 11200 28733 11203
rect 28684 11172 28733 11200
rect 28684 11160 28690 11172
rect 28721 11169 28733 11172
rect 28767 11169 28779 11203
rect 28721 11163 28779 11169
rect 29822 11160 29828 11212
rect 29880 11200 29886 11212
rect 30300 11209 30328 11240
rect 32306 11228 32312 11280
rect 32364 11228 32370 11280
rect 32582 11228 32588 11280
rect 32640 11268 32646 11280
rect 34514 11268 34520 11280
rect 32640 11240 34520 11268
rect 32640 11228 32646 11240
rect 34514 11228 34520 11240
rect 34572 11228 34578 11280
rect 34885 11271 34943 11277
rect 34885 11237 34897 11271
rect 34931 11268 34943 11271
rect 34931 11240 37136 11268
rect 34931 11237 34943 11240
rect 34885 11231 34943 11237
rect 30193 11203 30251 11209
rect 30193 11200 30205 11203
rect 29880 11172 30205 11200
rect 29880 11160 29886 11172
rect 30193 11169 30205 11172
rect 30239 11169 30251 11203
rect 30193 11163 30251 11169
rect 30285 11203 30343 11209
rect 30285 11169 30297 11203
rect 30331 11169 30343 11203
rect 30285 11163 30343 11169
rect 31570 11160 31576 11212
rect 31628 11160 31634 11212
rect 32766 11160 32772 11212
rect 32824 11160 32830 11212
rect 35158 11160 35164 11212
rect 35216 11200 35222 11212
rect 35437 11203 35495 11209
rect 35437 11200 35449 11203
rect 35216 11172 35449 11200
rect 35216 11160 35222 11172
rect 35437 11169 35449 11172
rect 35483 11169 35495 11203
rect 35437 11163 35495 11169
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11132 28595 11135
rect 29638 11132 29644 11144
rect 28583 11104 29644 11132
rect 28583 11101 28595 11104
rect 28537 11095 28595 11101
rect 29638 11092 29644 11104
rect 29696 11092 29702 11144
rect 30558 11092 30564 11144
rect 30616 11132 30622 11144
rect 31110 11132 31116 11144
rect 30616 11104 31116 11132
rect 30616 11092 30622 11104
rect 31110 11092 31116 11104
rect 31168 11092 31174 11144
rect 31297 11135 31355 11141
rect 31297 11101 31309 11135
rect 31343 11132 31355 11135
rect 31386 11132 31392 11144
rect 31343 11104 31392 11132
rect 31343 11101 31355 11104
rect 31297 11095 31355 11101
rect 31386 11092 31392 11104
rect 31444 11092 31450 11144
rect 32306 11092 32312 11144
rect 32364 11132 32370 11144
rect 32493 11135 32551 11141
rect 32493 11132 32505 11135
rect 32364 11104 32505 11132
rect 32364 11092 32370 11104
rect 32493 11101 32505 11104
rect 32539 11101 32551 11135
rect 32493 11095 32551 11101
rect 33413 11135 33471 11141
rect 33413 11101 33425 11135
rect 33459 11132 33471 11135
rect 35894 11132 35900 11144
rect 33459 11104 35900 11132
rect 33459 11101 33471 11104
rect 33413 11095 33471 11101
rect 35894 11092 35900 11104
rect 35952 11132 35958 11144
rect 36265 11135 36323 11141
rect 36265 11132 36277 11135
rect 35952 11104 36277 11132
rect 35952 11092 35958 11104
rect 36265 11101 36277 11104
rect 36311 11101 36323 11135
rect 36265 11095 36323 11101
rect 22066 11036 26004 11064
rect 25976 10996 26004 11036
rect 26602 11024 26608 11076
rect 26660 11024 26666 11076
rect 27617 11067 27675 11073
rect 27617 11064 27629 11067
rect 26896 11036 27629 11064
rect 26896 10996 26924 11036
rect 27617 11033 27629 11036
rect 27663 11064 27675 11067
rect 28629 11067 28687 11073
rect 28629 11064 28641 11067
rect 27663 11036 28641 11064
rect 27663 11033 27675 11036
rect 27617 11027 27675 11033
rect 28629 11033 28641 11036
rect 28675 11064 28687 11067
rect 29914 11064 29920 11076
rect 28675 11036 29920 11064
rect 28675 11033 28687 11036
rect 28629 11027 28687 11033
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 30101 11067 30159 11073
rect 30101 11033 30113 11067
rect 30147 11064 30159 11067
rect 31938 11064 31944 11076
rect 30147 11036 31944 11064
rect 30147 11033 30159 11036
rect 30101 11027 30159 11033
rect 31938 11024 31944 11036
rect 31996 11024 32002 11076
rect 32582 11024 32588 11076
rect 32640 11024 32646 11076
rect 34054 11024 34060 11076
rect 34112 11064 34118 11076
rect 34149 11067 34207 11073
rect 34149 11064 34161 11067
rect 34112 11036 34161 11064
rect 34112 11024 34118 11036
rect 34149 11033 34161 11036
rect 34195 11033 34207 11067
rect 34149 11027 34207 11033
rect 35250 11024 35256 11076
rect 35308 11024 35314 11076
rect 35342 11024 35348 11076
rect 35400 11024 35406 11076
rect 36998 11024 37004 11076
rect 37056 11024 37062 11076
rect 37108 11064 37136 11240
rect 37476 11200 37504 11308
rect 37645 11305 37657 11339
rect 37691 11336 37703 11339
rect 44358 11336 44364 11348
rect 37691 11308 44364 11336
rect 37691 11305 37703 11308
rect 37645 11299 37703 11305
rect 44358 11296 44364 11308
rect 44416 11296 44422 11348
rect 37918 11228 37924 11280
rect 37976 11268 37982 11280
rect 38838 11268 38844 11280
rect 37976 11240 38844 11268
rect 37976 11228 37982 11240
rect 38838 11228 38844 11240
rect 38896 11228 38902 11280
rect 39482 11200 39488 11212
rect 37476 11172 39488 11200
rect 39482 11160 39488 11172
rect 39540 11200 39546 11212
rect 40954 11200 40960 11212
rect 39540 11172 40960 11200
rect 39540 11160 39546 11172
rect 40954 11160 40960 11172
rect 41012 11160 41018 11212
rect 37826 11092 37832 11144
rect 37884 11092 37890 11144
rect 38654 11092 38660 11144
rect 38712 11092 38718 11144
rect 38930 11132 38936 11144
rect 38764 11104 38936 11132
rect 38764 11064 38792 11104
rect 38930 11092 38936 11104
rect 38988 11092 38994 11144
rect 37108 11036 38792 11064
rect 38838 11024 38844 11076
rect 38896 11024 38902 11076
rect 25976 10968 26924 10996
rect 28994 10956 29000 11008
rect 29052 10996 29058 11008
rect 31110 10996 31116 11008
rect 29052 10968 31116 10996
rect 29052 10956 29058 10968
rect 31110 10956 31116 10968
rect 31168 10956 31174 11008
rect 31389 10999 31447 11005
rect 31389 10965 31401 10999
rect 31435 10996 31447 10999
rect 31570 10996 31576 11008
rect 31435 10968 31576 10996
rect 31435 10965 31447 10968
rect 31389 10959 31447 10965
rect 31570 10956 31576 10968
rect 31628 10956 31634 11008
rect 32122 10956 32128 11008
rect 32180 10996 32186 11008
rect 37550 10996 37556 11008
rect 32180 10968 37556 10996
rect 32180 10956 32186 10968
rect 37550 10956 37556 10968
rect 37608 10956 37614 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 27154 10752 27160 10804
rect 27212 10792 27218 10804
rect 28353 10795 28411 10801
rect 28353 10792 28365 10795
rect 27212 10764 28365 10792
rect 27212 10752 27218 10764
rect 28353 10761 28365 10764
rect 28399 10761 28411 10795
rect 28353 10755 28411 10761
rect 29546 10752 29552 10804
rect 29604 10752 29610 10804
rect 29917 10795 29975 10801
rect 29917 10761 29929 10795
rect 29963 10792 29975 10795
rect 30098 10792 30104 10804
rect 29963 10764 30104 10792
rect 29963 10761 29975 10764
rect 29917 10755 29975 10761
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 31018 10752 31024 10804
rect 31076 10792 31082 10804
rect 31386 10792 31392 10804
rect 31076 10764 31392 10792
rect 31076 10752 31082 10764
rect 31386 10752 31392 10764
rect 31444 10792 31450 10804
rect 35621 10795 35679 10801
rect 31444 10764 32352 10792
rect 31444 10752 31450 10764
rect 30006 10684 30012 10736
rect 30064 10684 30070 10736
rect 28718 10616 28724 10668
rect 28776 10616 28782 10668
rect 30024 10656 30052 10684
rect 31113 10659 31171 10665
rect 30024 10628 30144 10656
rect 28810 10548 28816 10600
rect 28868 10548 28874 10600
rect 28905 10591 28963 10597
rect 28905 10557 28917 10591
rect 28951 10557 28963 10591
rect 28905 10551 28963 10557
rect 28442 10480 28448 10532
rect 28500 10520 28506 10532
rect 28920 10520 28948 10551
rect 29362 10548 29368 10600
rect 29420 10588 29426 10600
rect 30116 10597 30144 10628
rect 31113 10625 31125 10659
rect 31159 10656 31171 10659
rect 32122 10656 32128 10668
rect 31159 10628 32128 10656
rect 31159 10625 31171 10628
rect 31113 10619 31171 10625
rect 32122 10616 32128 10628
rect 32180 10616 32186 10668
rect 32324 10656 32352 10764
rect 32416 10764 35572 10792
rect 32416 10733 32444 10764
rect 32401 10727 32459 10733
rect 32401 10693 32413 10727
rect 32447 10693 32459 10727
rect 35544 10724 35572 10764
rect 35621 10761 35633 10795
rect 35667 10792 35679 10795
rect 40126 10792 40132 10804
rect 35667 10764 40132 10792
rect 35667 10761 35679 10764
rect 35621 10755 35679 10761
rect 40126 10752 40132 10764
rect 40184 10752 40190 10804
rect 35710 10724 35716 10736
rect 32401 10687 32459 10693
rect 32508 10696 33902 10724
rect 35544 10696 35716 10724
rect 32508 10656 32536 10696
rect 35710 10684 35716 10696
rect 35768 10684 35774 10736
rect 36078 10684 36084 10736
rect 36136 10684 36142 10736
rect 32324 10628 32536 10656
rect 35989 10659 36047 10665
rect 35989 10625 36001 10659
rect 36035 10625 36047 10659
rect 35989 10619 36047 10625
rect 30009 10591 30067 10597
rect 30009 10588 30021 10591
rect 29420 10560 30021 10588
rect 29420 10548 29426 10560
rect 30009 10557 30021 10560
rect 30055 10557 30067 10591
rect 30009 10551 30067 10557
rect 30101 10591 30159 10597
rect 30101 10557 30113 10591
rect 30147 10557 30159 10591
rect 30101 10551 30159 10557
rect 28500 10492 28948 10520
rect 30024 10520 30052 10551
rect 30742 10548 30748 10600
rect 30800 10588 30806 10600
rect 30926 10588 30932 10600
rect 30800 10560 30932 10588
rect 30800 10548 30806 10560
rect 30926 10548 30932 10560
rect 30984 10548 30990 10600
rect 31202 10548 31208 10600
rect 31260 10548 31266 10600
rect 31297 10591 31355 10597
rect 31297 10557 31309 10591
rect 31343 10588 31355 10591
rect 32766 10588 32772 10600
rect 31343 10560 32772 10588
rect 31343 10557 31355 10560
rect 31297 10551 31355 10557
rect 30190 10520 30196 10532
rect 30024 10492 30196 10520
rect 28500 10480 28506 10492
rect 30190 10480 30196 10492
rect 30248 10480 30254 10532
rect 31110 10480 31116 10532
rect 31168 10520 31174 10532
rect 31312 10520 31340 10551
rect 32766 10548 32772 10560
rect 32824 10548 32830 10600
rect 33137 10591 33195 10597
rect 33137 10557 33149 10591
rect 33183 10588 33195 10591
rect 33183 10560 33272 10588
rect 33183 10557 33195 10560
rect 33137 10551 33195 10557
rect 31168 10492 31340 10520
rect 31168 10480 31174 10492
rect 28902 10412 28908 10464
rect 28960 10452 28966 10464
rect 30745 10455 30803 10461
rect 30745 10452 30757 10455
rect 28960 10424 30757 10452
rect 28960 10412 28966 10424
rect 30745 10421 30757 10424
rect 30791 10421 30803 10455
rect 30745 10415 30803 10421
rect 31018 10412 31024 10464
rect 31076 10452 31082 10464
rect 32493 10455 32551 10461
rect 32493 10452 32505 10455
rect 31076 10424 32505 10452
rect 31076 10412 31082 10424
rect 32493 10421 32505 10424
rect 32539 10421 32551 10455
rect 33244 10452 33272 10560
rect 33410 10548 33416 10600
rect 33468 10548 33474 10600
rect 34146 10548 34152 10600
rect 34204 10588 34210 10600
rect 36004 10588 36032 10619
rect 40310 10616 40316 10668
rect 40368 10616 40374 10668
rect 42794 10616 42800 10668
rect 42852 10616 42858 10668
rect 45554 10616 45560 10668
rect 45612 10656 45618 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 45612 10628 47961 10656
rect 45612 10616 45618 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 34204 10560 36032 10588
rect 36265 10591 36323 10597
rect 34204 10548 34210 10560
rect 36265 10557 36277 10591
rect 36311 10557 36323 10591
rect 36265 10551 36323 10557
rect 34698 10480 34704 10532
rect 34756 10520 34762 10532
rect 34885 10523 34943 10529
rect 34885 10520 34897 10523
rect 34756 10492 34897 10520
rect 34756 10480 34762 10492
rect 34885 10489 34897 10492
rect 34931 10520 34943 10523
rect 35066 10520 35072 10532
rect 34931 10492 35072 10520
rect 34931 10489 34943 10492
rect 34885 10483 34943 10489
rect 35066 10480 35072 10492
rect 35124 10480 35130 10532
rect 36280 10520 36308 10551
rect 36998 10548 37004 10600
rect 37056 10588 37062 10600
rect 38933 10591 38991 10597
rect 38933 10588 38945 10591
rect 37056 10560 38945 10588
rect 37056 10548 37062 10560
rect 38933 10557 38945 10560
rect 38979 10557 38991 10591
rect 38933 10551 38991 10557
rect 39209 10591 39267 10597
rect 39209 10557 39221 10591
rect 39255 10588 39267 10591
rect 40678 10588 40684 10600
rect 39255 10560 40684 10588
rect 39255 10557 39267 10560
rect 39209 10551 39267 10557
rect 40678 10548 40684 10560
rect 40736 10548 40742 10600
rect 49142 10548 49148 10600
rect 49200 10548 49206 10600
rect 38746 10520 38752 10532
rect 36280 10492 38752 10520
rect 38746 10480 38752 10492
rect 38804 10480 38810 10532
rect 34790 10452 34796 10464
rect 33244 10424 34796 10452
rect 32493 10415 32551 10421
rect 34790 10412 34796 10424
rect 34848 10412 34854 10464
rect 36354 10412 36360 10464
rect 36412 10452 36418 10464
rect 37826 10452 37832 10464
rect 36412 10424 37832 10452
rect 36412 10412 36418 10424
rect 37826 10412 37832 10424
rect 37884 10412 37890 10464
rect 38764 10452 38792 10480
rect 40681 10455 40739 10461
rect 40681 10452 40693 10455
rect 38764 10424 40693 10452
rect 40681 10421 40693 10424
rect 40727 10421 40739 10455
rect 40681 10415 40739 10421
rect 42613 10455 42671 10461
rect 42613 10421 42625 10455
rect 42659 10452 42671 10455
rect 44082 10452 44088 10464
rect 42659 10424 44088 10452
rect 42659 10421 42671 10424
rect 42613 10415 42671 10421
rect 44082 10412 44088 10424
rect 44140 10412 44146 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 28718 10208 28724 10260
rect 28776 10248 28782 10260
rect 28776 10220 32352 10248
rect 28776 10208 28782 10220
rect 29822 10140 29828 10192
rect 29880 10180 29886 10192
rect 32324 10180 32352 10220
rect 32398 10208 32404 10260
rect 32456 10208 32462 10260
rect 32674 10208 32680 10260
rect 32732 10248 32738 10260
rect 32861 10251 32919 10257
rect 32861 10248 32873 10251
rect 32732 10220 32873 10248
rect 32732 10208 32738 10220
rect 32861 10217 32873 10220
rect 32907 10217 32919 10251
rect 32861 10211 32919 10217
rect 33318 10208 33324 10260
rect 33376 10248 33382 10260
rect 34146 10248 34152 10260
rect 33376 10220 34152 10248
rect 33376 10208 33382 10220
rect 34146 10208 34152 10220
rect 34204 10208 34210 10260
rect 36630 10208 36636 10260
rect 36688 10248 36694 10260
rect 37093 10251 37151 10257
rect 37093 10248 37105 10251
rect 36688 10220 37105 10248
rect 36688 10208 36694 10220
rect 37093 10217 37105 10220
rect 37139 10217 37151 10251
rect 37093 10211 37151 10217
rect 35342 10180 35348 10192
rect 29880 10152 30788 10180
rect 32324 10152 35348 10180
rect 29880 10140 29886 10152
rect 25314 10072 25320 10124
rect 25372 10112 25378 10124
rect 25774 10112 25780 10124
rect 25372 10084 25780 10112
rect 25372 10072 25378 10084
rect 25774 10072 25780 10084
rect 25832 10072 25838 10124
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10112 26111 10115
rect 29454 10112 29460 10124
rect 26099 10084 29460 10112
rect 26099 10081 26111 10084
rect 26053 10075 26111 10081
rect 29454 10072 29460 10084
rect 29512 10072 29518 10124
rect 29730 10072 29736 10124
rect 29788 10112 29794 10124
rect 30653 10115 30711 10121
rect 30653 10112 30665 10115
rect 29788 10084 30665 10112
rect 29788 10072 29794 10084
rect 30653 10081 30665 10084
rect 30699 10081 30711 10115
rect 30760 10112 30788 10152
rect 35342 10140 35348 10152
rect 35400 10140 35406 10192
rect 32306 10112 32312 10124
rect 30760 10084 32312 10112
rect 30653 10075 30711 10081
rect 32306 10072 32312 10084
rect 32364 10072 32370 10124
rect 32766 10072 32772 10124
rect 32824 10112 32830 10124
rect 33413 10115 33471 10121
rect 33413 10112 33425 10115
rect 32824 10084 33425 10112
rect 32824 10072 32830 10084
rect 33413 10081 33425 10084
rect 33459 10081 33471 10115
rect 36998 10112 37004 10124
rect 33413 10075 33471 10081
rect 35360 10084 37004 10112
rect 34882 10004 34888 10056
rect 34940 10044 34946 10056
rect 35360 10053 35388 10084
rect 36998 10072 37004 10084
rect 37056 10072 37062 10124
rect 35345 10047 35403 10053
rect 35345 10044 35357 10047
rect 34940 10016 35357 10044
rect 34940 10004 34946 10016
rect 35345 10013 35357 10016
rect 35391 10013 35403 10047
rect 37182 10044 37188 10056
rect 36754 10016 37188 10044
rect 35345 10007 35403 10013
rect 37182 10004 37188 10016
rect 37240 10004 37246 10056
rect 37737 10047 37795 10053
rect 37737 10013 37749 10047
rect 37783 10044 37795 10047
rect 38654 10044 38660 10056
rect 37783 10016 38660 10044
rect 37783 10013 37795 10016
rect 37737 10007 37795 10013
rect 38654 10004 38660 10016
rect 38712 10004 38718 10056
rect 38749 10047 38807 10053
rect 38749 10013 38761 10047
rect 38795 10013 38807 10047
rect 38749 10007 38807 10013
rect 26602 9936 26608 9988
rect 26660 9936 26666 9988
rect 30926 9936 30932 9988
rect 30984 9936 30990 9988
rect 31386 9936 31392 9988
rect 31444 9936 31450 9988
rect 32214 9936 32220 9988
rect 32272 9976 32278 9988
rect 32272 9948 33456 9976
rect 32272 9936 32278 9948
rect 27522 9868 27528 9920
rect 27580 9868 27586 9920
rect 29546 9868 29552 9920
rect 29604 9908 29610 9920
rect 31018 9908 31024 9920
rect 29604 9880 31024 9908
rect 29604 9868 29610 9880
rect 31018 9868 31024 9880
rect 31076 9868 31082 9920
rect 33226 9868 33232 9920
rect 33284 9868 33290 9920
rect 33318 9868 33324 9920
rect 33376 9868 33382 9920
rect 33428 9908 33456 9948
rect 34606 9936 34612 9988
rect 34664 9976 34670 9988
rect 35066 9976 35072 9988
rect 34664 9948 35072 9976
rect 34664 9936 34670 9948
rect 35066 9936 35072 9948
rect 35124 9936 35130 9988
rect 35621 9979 35679 9985
rect 35621 9945 35633 9979
rect 35667 9976 35679 9979
rect 35710 9976 35716 9988
rect 35667 9948 35716 9976
rect 35667 9945 35679 9948
rect 35621 9939 35679 9945
rect 35710 9936 35716 9948
rect 35768 9936 35774 9988
rect 38764 9976 38792 10007
rect 44634 10004 44640 10056
rect 44692 10044 44698 10056
rect 46845 10047 46903 10053
rect 46845 10044 46857 10047
rect 44692 10016 46857 10044
rect 44692 10004 44698 10016
rect 46845 10013 46857 10016
rect 46891 10013 46903 10047
rect 46845 10007 46903 10013
rect 46934 10004 46940 10056
rect 46992 10044 46998 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 46992 10016 47961 10044
rect 46992 10004 46998 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 36924 9948 38792 9976
rect 36924 9908 36952 9948
rect 44174 9936 44180 9988
rect 44232 9976 44238 9988
rect 46109 9979 46167 9985
rect 46109 9976 46121 9979
rect 44232 9948 46121 9976
rect 44232 9936 44238 9948
rect 46109 9945 46121 9948
rect 46155 9945 46167 9979
rect 46109 9939 46167 9945
rect 46290 9936 46296 9988
rect 46348 9936 46354 9988
rect 47026 9936 47032 9988
rect 47084 9936 47090 9988
rect 49142 9936 49148 9988
rect 49200 9936 49206 9988
rect 33428 9880 36952 9908
rect 38565 9911 38623 9917
rect 38565 9877 38577 9911
rect 38611 9908 38623 9911
rect 40402 9908 40408 9920
rect 38611 9880 40408 9908
rect 38611 9877 38623 9880
rect 38565 9871 38623 9877
rect 40402 9868 40408 9880
rect 40460 9868 40466 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 29564 9676 30420 9704
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 24394 9636 24400 9648
rect 3476 9608 24400 9636
rect 3476 9596 3482 9608
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 29564 9636 29592 9676
rect 24504 9608 29592 9636
rect 29641 9639 29699 9645
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 24504 9568 24532 9608
rect 29641 9605 29653 9639
rect 29687 9636 29699 9639
rect 30282 9636 30288 9648
rect 29687 9608 30288 9636
rect 29687 9605 29699 9608
rect 29641 9599 29699 9605
rect 30282 9596 30288 9608
rect 30340 9596 30346 9648
rect 30392 9636 30420 9676
rect 31478 9664 31484 9716
rect 31536 9704 31542 9716
rect 32582 9704 32588 9716
rect 31536 9676 32588 9704
rect 31536 9664 31542 9676
rect 32582 9664 32588 9676
rect 32640 9664 32646 9716
rect 33226 9664 33232 9716
rect 33284 9704 33290 9716
rect 39114 9704 39120 9716
rect 33284 9676 39120 9704
rect 33284 9664 33290 9676
rect 39114 9664 39120 9676
rect 39172 9664 39178 9716
rect 30650 9636 30656 9648
rect 30392 9608 30656 9636
rect 30650 9596 30656 9608
rect 30708 9596 30714 9648
rect 30837 9639 30895 9645
rect 30837 9605 30849 9639
rect 30883 9636 30895 9639
rect 34790 9636 34796 9648
rect 30883 9608 34796 9636
rect 30883 9605 30895 9608
rect 30837 9599 30895 9605
rect 34790 9596 34796 9608
rect 34848 9596 34854 9648
rect 36173 9639 36231 9645
rect 36173 9605 36185 9639
rect 36219 9636 36231 9639
rect 38378 9636 38384 9648
rect 36219 9608 38384 9636
rect 36219 9605 36231 9608
rect 36173 9599 36231 9605
rect 38378 9596 38384 9608
rect 38436 9596 38442 9648
rect 38746 9596 38752 9648
rect 38804 9596 38810 9648
rect 39022 9596 39028 9648
rect 39080 9636 39086 9648
rect 39080 9608 39238 9636
rect 39080 9596 39086 9608
rect 22796 9540 24532 9568
rect 22796 9528 22802 9540
rect 29086 9528 29092 9580
rect 29144 9568 29150 9580
rect 29733 9571 29791 9577
rect 29733 9568 29745 9571
rect 29144 9540 29745 9568
rect 29144 9528 29150 9540
rect 29733 9537 29745 9540
rect 29779 9537 29791 9571
rect 29733 9531 29791 9537
rect 30024 9540 31064 9568
rect 25130 9460 25136 9512
rect 25188 9500 25194 9512
rect 25188 9472 29132 9500
rect 25188 9460 25194 9472
rect 23934 9392 23940 9444
rect 23992 9432 23998 9444
rect 28994 9432 29000 9444
rect 23992 9404 29000 9432
rect 23992 9392 23998 9404
rect 28994 9392 29000 9404
rect 29052 9392 29058 9444
rect 23290 9324 23296 9376
rect 23348 9324 23354 9376
rect 26418 9324 26424 9376
rect 26476 9324 26482 9376
rect 28810 9324 28816 9376
rect 28868 9324 28874 9376
rect 29104 9364 29132 9472
rect 29270 9392 29276 9444
rect 29328 9392 29334 9444
rect 29748 9432 29776 9531
rect 30024 9512 30052 9540
rect 29917 9503 29975 9509
rect 29917 9469 29929 9503
rect 29963 9500 29975 9503
rect 30006 9500 30012 9512
rect 29963 9472 30012 9500
rect 29963 9469 29975 9472
rect 29917 9463 29975 9469
rect 30006 9460 30012 9472
rect 30064 9460 30070 9512
rect 30558 9460 30564 9512
rect 30616 9500 30622 9512
rect 31036 9509 31064 9540
rect 31110 9528 31116 9580
rect 31168 9568 31174 9580
rect 33137 9571 33195 9577
rect 33137 9568 33149 9571
rect 31168 9540 33149 9568
rect 31168 9528 31174 9540
rect 33137 9537 33149 9540
rect 33183 9537 33195 9571
rect 33137 9531 33195 9537
rect 34977 9571 35035 9577
rect 34977 9537 34989 9571
rect 35023 9537 35035 9571
rect 34977 9531 35035 9537
rect 30929 9503 30987 9509
rect 30929 9500 30941 9503
rect 30616 9472 30941 9500
rect 30616 9460 30622 9472
rect 30929 9469 30941 9472
rect 30975 9469 30987 9503
rect 30929 9463 30987 9469
rect 31021 9503 31079 9509
rect 31021 9469 31033 9503
rect 31067 9469 31079 9503
rect 33226 9500 33232 9512
rect 31021 9463 31079 9469
rect 31128 9472 33232 9500
rect 30374 9432 30380 9444
rect 29748 9404 30380 9432
rect 30374 9392 30380 9404
rect 30432 9392 30438 9444
rect 30466 9392 30472 9444
rect 30524 9392 30530 9444
rect 31128 9364 31156 9472
rect 33226 9460 33232 9472
rect 33284 9460 33290 9512
rect 33413 9503 33471 9509
rect 33413 9469 33425 9503
rect 33459 9500 33471 9503
rect 34514 9500 34520 9512
rect 33459 9472 34520 9500
rect 33459 9469 33471 9472
rect 33413 9463 33471 9469
rect 34514 9460 34520 9472
rect 34572 9460 34578 9512
rect 31662 9392 31668 9444
rect 31720 9432 31726 9444
rect 34992 9432 35020 9531
rect 35066 9528 35072 9580
rect 35124 9528 35130 9580
rect 36998 9528 37004 9580
rect 37056 9568 37062 9580
rect 38473 9571 38531 9577
rect 38473 9568 38485 9571
rect 37056 9540 38485 9568
rect 37056 9528 37062 9540
rect 38473 9537 38485 9540
rect 38519 9537 38531 9571
rect 38473 9531 38531 9537
rect 43714 9528 43720 9580
rect 43772 9528 43778 9580
rect 44082 9528 44088 9580
rect 44140 9568 44146 9580
rect 46477 9571 46535 9577
rect 46477 9568 46489 9571
rect 44140 9540 46489 9568
rect 44140 9528 44146 9540
rect 46477 9537 46489 9540
rect 46523 9537 46535 9571
rect 46477 9531 46535 9537
rect 35253 9503 35311 9509
rect 35253 9469 35265 9503
rect 35299 9500 35311 9503
rect 36446 9500 36452 9512
rect 35299 9472 36452 9500
rect 35299 9469 35311 9472
rect 35253 9463 35311 9469
rect 36446 9460 36452 9472
rect 36504 9460 36510 9512
rect 36722 9460 36728 9512
rect 36780 9500 36786 9512
rect 40034 9500 40040 9512
rect 36780 9472 40040 9500
rect 36780 9460 36786 9472
rect 40034 9460 40040 9472
rect 40092 9460 40098 9512
rect 31720 9404 35020 9432
rect 36188 9404 36492 9432
rect 31720 9392 31726 9404
rect 29104 9336 31156 9364
rect 32766 9324 32772 9376
rect 32824 9324 32830 9376
rect 34609 9367 34667 9373
rect 34609 9333 34621 9367
rect 34655 9364 34667 9367
rect 36188 9364 36216 9404
rect 34655 9336 36216 9364
rect 34655 9333 34667 9336
rect 34609 9327 34667 9333
rect 36262 9324 36268 9376
rect 36320 9324 36326 9376
rect 36464 9364 36492 9404
rect 36740 9404 38608 9432
rect 36740 9364 36768 9404
rect 36464 9336 36768 9364
rect 37458 9324 37464 9376
rect 37516 9364 37522 9376
rect 37645 9367 37703 9373
rect 37645 9364 37657 9367
rect 37516 9336 37657 9364
rect 37516 9324 37522 9336
rect 37645 9333 37657 9336
rect 37691 9333 37703 9367
rect 38580 9364 38608 9404
rect 39114 9364 39120 9376
rect 38580 9336 39120 9364
rect 37645 9327 37703 9333
rect 39114 9324 39120 9336
rect 39172 9324 39178 9376
rect 40218 9324 40224 9376
rect 40276 9324 40282 9376
rect 43533 9367 43591 9373
rect 43533 9333 43545 9367
rect 43579 9364 43591 9367
rect 45462 9364 45468 9376
rect 43579 9336 45468 9364
rect 43579 9333 43591 9336
rect 43533 9327 43591 9333
rect 45462 9324 45468 9336
rect 45520 9324 45526 9376
rect 46293 9367 46351 9373
rect 46293 9333 46305 9367
rect 46339 9364 46351 9367
rect 47854 9364 47860 9376
rect 46339 9336 47860 9364
rect 46339 9333 46351 9336
rect 46293 9327 46351 9333
rect 47854 9324 47860 9336
rect 47912 9324 47918 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 22738 9120 22744 9172
rect 22796 9120 22802 9172
rect 34698 9160 34704 9172
rect 23400 9132 34704 9160
rect 23400 9033 23428 9132
rect 34698 9120 34704 9132
rect 34756 9120 34762 9172
rect 35710 9120 35716 9172
rect 35768 9160 35774 9172
rect 45373 9163 45431 9169
rect 35768 9132 37688 9160
rect 35768 9120 35774 9132
rect 27062 9052 27068 9104
rect 27120 9092 27126 9104
rect 27120 9064 27660 9092
rect 27120 9052 27126 9064
rect 23385 9027 23443 9033
rect 23385 8993 23397 9027
rect 23431 8993 23443 9027
rect 23385 8987 23443 8993
rect 24118 8984 24124 9036
rect 24176 9024 24182 9036
rect 25593 9027 25651 9033
rect 25593 9024 25605 9027
rect 24176 8996 25605 9024
rect 24176 8984 24182 8996
rect 25593 8993 25605 8996
rect 25639 9024 25651 9027
rect 27522 9024 27528 9036
rect 25639 8996 27528 9024
rect 25639 8993 25651 8996
rect 25593 8987 25651 8993
rect 27522 8984 27528 8996
rect 27580 8984 27586 9036
rect 27632 9024 27660 9064
rect 28350 9052 28356 9104
rect 28408 9092 28414 9104
rect 28445 9095 28503 9101
rect 28445 9092 28457 9095
rect 28408 9064 28457 9092
rect 28408 9052 28414 9064
rect 28445 9061 28457 9064
rect 28491 9061 28503 9095
rect 28445 9055 28503 9061
rect 31938 9052 31944 9104
rect 31996 9052 32002 9104
rect 37093 9095 37151 9101
rect 37093 9061 37105 9095
rect 37139 9092 37151 9095
rect 37274 9092 37280 9104
rect 37139 9064 37280 9092
rect 37139 9061 37151 9064
rect 37093 9055 37151 9061
rect 37274 9052 37280 9064
rect 37332 9052 37338 9104
rect 28997 9027 29055 9033
rect 28997 9024 29009 9027
rect 27632 8996 29009 9024
rect 28997 8993 29009 8996
rect 29043 8993 29055 9027
rect 28997 8987 29055 8993
rect 29730 8984 29736 9036
rect 29788 8984 29794 9036
rect 30009 9027 30067 9033
rect 30009 8993 30021 9027
rect 30055 9024 30067 9027
rect 31846 9024 31852 9036
rect 30055 8996 31852 9024
rect 30055 8993 30067 8996
rect 30009 8987 30067 8993
rect 31846 8984 31852 8996
rect 31904 8984 31910 9036
rect 32122 8984 32128 9036
rect 32180 9024 32186 9036
rect 32401 9027 32459 9033
rect 32401 9024 32413 9027
rect 32180 8996 32413 9024
rect 32180 8984 32186 8996
rect 32401 8993 32413 8996
rect 32447 8993 32459 9027
rect 32401 8987 32459 8993
rect 32582 8984 32588 9036
rect 32640 8984 32646 9036
rect 32766 8984 32772 9036
rect 32824 9024 32830 9036
rect 37660 9033 37688 9132
rect 45373 9129 45385 9163
rect 45419 9160 45431 9163
rect 45554 9160 45560 9172
rect 45419 9132 45560 9160
rect 45419 9129 45431 9132
rect 45373 9123 45431 9129
rect 45554 9120 45560 9132
rect 45612 9120 45618 9172
rect 45925 9163 45983 9169
rect 45925 9129 45937 9163
rect 45971 9160 45983 9163
rect 46934 9160 46940 9172
rect 45971 9132 46940 9160
rect 45971 9129 45983 9132
rect 45925 9123 45983 9129
rect 46934 9120 46940 9132
rect 46992 9120 46998 9172
rect 38289 9095 38347 9101
rect 38289 9061 38301 9095
rect 38335 9092 38347 9095
rect 40034 9092 40040 9104
rect 38335 9064 40040 9092
rect 38335 9061 38347 9064
rect 38289 9055 38347 9061
rect 40034 9052 40040 9064
rect 40092 9052 40098 9104
rect 41233 9095 41291 9101
rect 41233 9061 41245 9095
rect 41279 9092 41291 9095
rect 41279 9064 46888 9092
rect 41279 9061 41291 9064
rect 41233 9055 41291 9061
rect 37553 9027 37611 9033
rect 37553 9024 37565 9027
rect 32824 8996 37565 9024
rect 32824 8984 32830 8996
rect 37553 8993 37565 8996
rect 37599 8993 37611 9027
rect 37553 8987 37611 8993
rect 37645 9027 37703 9033
rect 37645 8993 37657 9027
rect 37691 8993 37703 9027
rect 38841 9027 38899 9033
rect 38841 9024 38853 9027
rect 37645 8987 37703 8993
rect 37752 8996 38853 9024
rect 22281 8959 22339 8965
rect 22281 8956 22293 8959
rect 22066 8928 22293 8956
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 22066 8820 22094 8928
rect 22281 8925 22293 8928
rect 22327 8956 22339 8959
rect 23201 8959 23259 8965
rect 23201 8956 23213 8959
rect 22327 8928 23213 8956
rect 22327 8925 22339 8928
rect 22281 8919 22339 8925
rect 23201 8925 23213 8928
rect 23247 8925 23259 8959
rect 23201 8919 23259 8925
rect 24762 8916 24768 8968
rect 24820 8956 24826 8968
rect 25317 8959 25375 8965
rect 25317 8956 25329 8959
rect 24820 8928 25329 8956
rect 24820 8916 24826 8928
rect 25317 8925 25329 8928
rect 25363 8925 25375 8959
rect 25317 8919 25375 8925
rect 28810 8916 28816 8968
rect 28868 8916 28874 8968
rect 31386 8956 31392 8968
rect 31142 8928 31392 8956
rect 31386 8916 31392 8928
rect 31444 8916 31450 8968
rect 33229 8959 33287 8965
rect 33229 8925 33241 8959
rect 33275 8956 33287 8959
rect 34422 8956 34428 8968
rect 33275 8928 34428 8956
rect 33275 8925 33287 8928
rect 33229 8919 33287 8925
rect 34422 8916 34428 8928
rect 34480 8916 34486 8968
rect 34882 8916 34888 8968
rect 34940 8916 34946 8968
rect 36170 8916 36176 8968
rect 36228 8956 36234 8968
rect 36998 8956 37004 8968
rect 36228 8928 37004 8956
rect 36228 8916 36234 8928
rect 36998 8916 37004 8928
rect 37056 8916 37062 8968
rect 37752 8956 37780 8996
rect 38841 8993 38853 8996
rect 38887 8993 38899 9027
rect 38841 8987 38899 8993
rect 37108 8928 37780 8956
rect 23109 8891 23167 8897
rect 23109 8857 23121 8891
rect 23155 8888 23167 8891
rect 23290 8888 23296 8900
rect 23155 8860 23296 8888
rect 23155 8857 23167 8860
rect 23109 8851 23167 8857
rect 23290 8848 23296 8860
rect 23348 8848 23354 8900
rect 26602 8848 26608 8900
rect 26660 8848 26666 8900
rect 28905 8891 28963 8897
rect 28905 8888 28917 8891
rect 26896 8860 28917 8888
rect 2648 8792 22094 8820
rect 2648 8780 2654 8792
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 26896 8820 26924 8860
rect 28905 8857 28917 8860
rect 28951 8857 28963 8891
rect 28905 8851 28963 8857
rect 35158 8848 35164 8900
rect 35216 8848 35222 8900
rect 23532 8792 26924 8820
rect 23532 8780 23538 8792
rect 31478 8780 31484 8832
rect 31536 8780 31542 8832
rect 32309 8823 32367 8829
rect 32309 8789 32321 8823
rect 32355 8820 32367 8823
rect 32582 8820 32588 8832
rect 32355 8792 32588 8820
rect 32355 8789 32367 8792
rect 32309 8783 32367 8789
rect 32582 8780 32588 8792
rect 32640 8780 32646 8832
rect 33134 8780 33140 8832
rect 33192 8820 33198 8832
rect 33321 8823 33379 8829
rect 33321 8820 33333 8823
rect 33192 8792 33333 8820
rect 33192 8780 33198 8792
rect 33321 8789 33333 8792
rect 33367 8789 33379 8823
rect 33321 8783 33379 8789
rect 33410 8780 33416 8832
rect 33468 8820 33474 8832
rect 36633 8823 36691 8829
rect 36633 8820 36645 8823
rect 33468 8792 36645 8820
rect 33468 8780 33474 8792
rect 36633 8789 36645 8792
rect 36679 8820 36691 8823
rect 37108 8820 37136 8928
rect 38654 8916 38660 8968
rect 38712 8916 38718 8968
rect 38749 8959 38807 8965
rect 38749 8925 38761 8959
rect 38795 8956 38807 8959
rect 38930 8956 38936 8968
rect 38795 8928 38936 8956
rect 38795 8925 38807 8928
rect 38749 8919 38807 8925
rect 38930 8916 38936 8928
rect 38988 8916 38994 8968
rect 40221 8959 40279 8965
rect 40221 8925 40233 8959
rect 40267 8956 40279 8959
rect 40310 8956 40316 8968
rect 40267 8928 40316 8956
rect 40267 8925 40279 8928
rect 40221 8919 40279 8925
rect 40310 8916 40316 8928
rect 40368 8916 40374 8968
rect 41417 8959 41475 8965
rect 41417 8925 41429 8959
rect 41463 8925 41475 8959
rect 41417 8919 41475 8925
rect 37458 8848 37464 8900
rect 37516 8848 37522 8900
rect 38470 8848 38476 8900
rect 38528 8888 38534 8900
rect 39022 8888 39028 8900
rect 38528 8860 39028 8888
rect 38528 8848 38534 8860
rect 39022 8848 39028 8860
rect 39080 8848 39086 8900
rect 36679 8792 37136 8820
rect 36679 8789 36691 8792
rect 36633 8783 36691 8789
rect 37274 8780 37280 8832
rect 37332 8820 37338 8832
rect 41432 8820 41460 8919
rect 44174 8916 44180 8968
rect 44232 8956 44238 8968
rect 46860 8965 46888 9064
rect 46109 8959 46167 8965
rect 46109 8956 46121 8959
rect 44232 8928 46121 8956
rect 44232 8916 44238 8928
rect 46109 8925 46121 8928
rect 46155 8925 46167 8959
rect 46109 8919 46167 8925
rect 46845 8959 46903 8965
rect 46845 8925 46857 8959
rect 46891 8925 46903 8959
rect 46845 8919 46903 8925
rect 47949 8959 48007 8965
rect 47949 8925 47961 8959
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 45278 8848 45284 8900
rect 45336 8848 45342 8900
rect 37332 8792 41460 8820
rect 46661 8823 46719 8829
rect 37332 8780 37338 8792
rect 46661 8789 46673 8823
rect 46707 8820 46719 8823
rect 47964 8820 47992 8919
rect 49142 8848 49148 8900
rect 49200 8848 49206 8900
rect 46707 8792 47992 8820
rect 46707 8789 46719 8792
rect 46661 8783 46719 8789
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 23474 8576 23480 8628
rect 23532 8576 23538 8628
rect 23934 8576 23940 8628
rect 23992 8576 23998 8628
rect 24673 8619 24731 8625
rect 24673 8585 24685 8619
rect 24719 8616 24731 8619
rect 30929 8619 30987 8625
rect 24719 8588 29224 8616
rect 24719 8585 24731 8588
rect 24673 8579 24731 8585
rect 18506 8508 18512 8560
rect 18564 8548 18570 8560
rect 25041 8551 25099 8557
rect 25041 8548 25053 8551
rect 18564 8520 25053 8548
rect 18564 8508 18570 8520
rect 25041 8517 25053 8520
rect 25087 8517 25099 8551
rect 25041 8511 25099 8517
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 22066 8452 23029 8480
rect 22066 8356 22094 8452
rect 23017 8449 23029 8452
rect 23063 8480 23075 8483
rect 23845 8483 23903 8489
rect 23845 8480 23857 8483
rect 23063 8452 23857 8480
rect 23063 8449 23075 8452
rect 23017 8443 23075 8449
rect 23845 8449 23857 8452
rect 23891 8449 23903 8483
rect 25056 8480 25084 8511
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 25774 8508 25780 8560
rect 25832 8548 25838 8560
rect 27522 8548 27528 8560
rect 25832 8520 27528 8548
rect 25832 8508 25838 8520
rect 27522 8508 27528 8520
rect 27580 8508 27586 8560
rect 29196 8548 29224 8588
rect 30929 8585 30941 8619
rect 30975 8616 30987 8619
rect 30975 8588 31754 8616
rect 30975 8585 30987 8588
rect 30929 8579 30987 8585
rect 31389 8551 31447 8557
rect 31389 8548 31401 8551
rect 27632 8520 28382 8548
rect 29196 8520 31401 8548
rect 25869 8483 25927 8489
rect 25869 8480 25881 8483
rect 25056 8452 25881 8480
rect 23845 8443 23903 8449
rect 25869 8449 25881 8452
rect 25915 8449 25927 8483
rect 25869 8443 25927 8449
rect 26418 8440 26424 8492
rect 26476 8440 26482 8492
rect 26602 8440 26608 8492
rect 26660 8480 26666 8492
rect 27632 8480 27660 8520
rect 31389 8517 31401 8520
rect 31435 8517 31447 8551
rect 31726 8548 31754 8588
rect 32306 8576 32312 8628
rect 32364 8576 32370 8628
rect 32677 8619 32735 8625
rect 32677 8585 32689 8619
rect 32723 8616 32735 8619
rect 34422 8616 34428 8628
rect 32723 8588 34428 8616
rect 32723 8585 32735 8588
rect 32677 8579 32735 8585
rect 34422 8576 34428 8588
rect 34480 8576 34486 8628
rect 34514 8576 34520 8628
rect 34572 8576 34578 8628
rect 35250 8576 35256 8628
rect 35308 8616 35314 8628
rect 35308 8588 35664 8616
rect 35308 8576 35314 8588
rect 34333 8551 34391 8557
rect 31726 8520 34008 8548
rect 31389 8511 31447 8517
rect 26660 8452 27660 8480
rect 31297 8483 31355 8489
rect 26660 8440 26666 8452
rect 31297 8449 31309 8483
rect 31343 8480 31355 8483
rect 32306 8480 32312 8492
rect 31343 8452 32312 8480
rect 31343 8449 31355 8452
rect 31297 8443 31355 8449
rect 32306 8440 32312 8452
rect 32364 8440 32370 8492
rect 32674 8440 32680 8492
rect 32732 8480 32738 8492
rect 32732 8452 32904 8480
rect 32732 8440 32738 8452
rect 24118 8372 24124 8424
rect 24176 8372 24182 8424
rect 25317 8415 25375 8421
rect 25317 8381 25329 8415
rect 25363 8381 25375 8415
rect 25317 8375 25375 8381
rect 22002 8304 22008 8356
rect 22060 8316 22094 8356
rect 25332 8344 25360 8375
rect 26234 8372 26240 8424
rect 26292 8412 26298 8424
rect 26513 8415 26571 8421
rect 26513 8412 26525 8415
rect 26292 8384 26525 8412
rect 26292 8372 26298 8384
rect 26513 8381 26525 8384
rect 26559 8381 26571 8415
rect 26513 8375 26571 8381
rect 26694 8372 26700 8424
rect 26752 8372 26758 8424
rect 27614 8372 27620 8424
rect 27672 8421 27678 8424
rect 27672 8412 27682 8421
rect 29365 8415 29423 8421
rect 27672 8384 27717 8412
rect 27672 8375 27682 8384
rect 29365 8381 29377 8415
rect 29411 8412 29423 8415
rect 30926 8412 30932 8424
rect 29411 8384 30932 8412
rect 29411 8381 29423 8384
rect 29365 8375 29423 8381
rect 27672 8372 27678 8375
rect 30926 8372 30932 8384
rect 30984 8412 30990 8424
rect 31481 8415 31539 8421
rect 31481 8412 31493 8415
rect 30984 8384 31493 8412
rect 30984 8372 30990 8384
rect 31481 8381 31493 8384
rect 31527 8381 31539 8415
rect 31481 8375 31539 8381
rect 31662 8372 31668 8424
rect 31720 8412 31726 8424
rect 32876 8421 32904 8452
rect 32769 8415 32827 8421
rect 32769 8412 32781 8415
rect 31720 8384 32781 8412
rect 31720 8372 31754 8384
rect 32769 8381 32781 8384
rect 32815 8381 32827 8415
rect 32769 8375 32827 8381
rect 32861 8415 32919 8421
rect 32861 8381 32873 8415
rect 32907 8381 32919 8415
rect 33980 8412 34008 8520
rect 34333 8517 34345 8551
rect 34379 8548 34391 8551
rect 34532 8548 34560 8576
rect 35636 8548 35664 8588
rect 35710 8576 35716 8628
rect 35768 8616 35774 8628
rect 35805 8619 35863 8625
rect 35805 8616 35817 8619
rect 35768 8588 35817 8616
rect 35768 8576 35774 8588
rect 35805 8585 35817 8588
rect 35851 8585 35863 8619
rect 35805 8579 35863 8585
rect 36446 8576 36452 8628
rect 36504 8616 36510 8628
rect 39485 8619 39543 8625
rect 39485 8616 39497 8619
rect 36504 8588 39497 8616
rect 36504 8576 36510 8588
rect 39485 8585 39497 8588
rect 39531 8585 39543 8619
rect 39485 8579 39543 8585
rect 40310 8576 40316 8628
rect 40368 8576 40374 8628
rect 36170 8548 36176 8560
rect 34379 8520 34560 8548
rect 35558 8520 36176 8548
rect 34379 8517 34391 8520
rect 34333 8511 34391 8517
rect 36170 8508 36176 8520
rect 36228 8508 36234 8560
rect 36722 8508 36728 8560
rect 36780 8508 36786 8560
rect 37182 8508 37188 8560
rect 37240 8548 37246 8560
rect 38470 8548 38476 8560
rect 37240 8520 38476 8548
rect 37240 8508 37246 8520
rect 38470 8508 38476 8520
rect 38528 8508 38534 8560
rect 40126 8508 40132 8560
rect 40184 8548 40190 8560
rect 40405 8551 40463 8557
rect 40405 8548 40417 8551
rect 40184 8520 40417 8548
rect 40184 8508 40190 8520
rect 40405 8517 40417 8520
rect 40451 8517 40463 8551
rect 40405 8511 40463 8517
rect 45186 8508 45192 8560
rect 45244 8548 45250 8560
rect 46661 8551 46719 8557
rect 46661 8548 46673 8551
rect 45244 8520 46673 8548
rect 45244 8508 45250 8520
rect 46661 8517 46673 8520
rect 46707 8517 46719 8551
rect 46661 8511 46719 8517
rect 34054 8440 34060 8492
rect 34112 8440 34118 8492
rect 36354 8480 36360 8492
rect 35544 8452 36360 8480
rect 35544 8412 35572 8452
rect 36354 8440 36360 8452
rect 36412 8440 36418 8492
rect 40218 8440 40224 8492
rect 40276 8480 40282 8492
rect 40276 8452 40540 8480
rect 40276 8440 40282 8452
rect 33980 8384 35572 8412
rect 32861 8375 32919 8381
rect 35802 8372 35808 8424
rect 35860 8412 35866 8424
rect 37737 8415 37795 8421
rect 37737 8412 37749 8415
rect 35860 8384 37749 8412
rect 35860 8372 35866 8384
rect 37737 8381 37749 8384
rect 37783 8381 37795 8415
rect 37737 8375 37795 8381
rect 38013 8415 38071 8421
rect 38013 8381 38025 8415
rect 38059 8412 38071 8415
rect 40328 8412 40356 8452
rect 40512 8421 40540 8452
rect 47854 8440 47860 8492
rect 47912 8480 47918 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 47912 8452 47961 8480
rect 47912 8440 47918 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 38059 8384 40356 8412
rect 40497 8415 40555 8421
rect 38059 8381 38071 8384
rect 38013 8375 38071 8381
rect 40497 8381 40509 8415
rect 40543 8381 40555 8415
rect 40497 8375 40555 8381
rect 49142 8372 49148 8424
rect 49200 8372 49206 8424
rect 25332 8316 27660 8344
rect 22060 8304 22066 8316
rect 26053 8279 26111 8285
rect 26053 8245 26065 8279
rect 26099 8276 26111 8279
rect 26142 8276 26148 8288
rect 26099 8248 26148 8276
rect 26099 8245 26111 8248
rect 26053 8239 26111 8245
rect 26142 8236 26148 8248
rect 26200 8236 26206 8288
rect 27632 8276 27660 8316
rect 30650 8304 30656 8356
rect 30708 8344 30714 8356
rect 31726 8344 31754 8372
rect 30708 8316 31754 8344
rect 30708 8304 30714 8316
rect 35342 8304 35348 8356
rect 35400 8344 35406 8356
rect 36909 8347 36967 8353
rect 36909 8344 36921 8347
rect 35400 8316 36921 8344
rect 35400 8304 35406 8316
rect 36909 8313 36921 8316
rect 36955 8313 36967 8347
rect 36909 8307 36967 8313
rect 39945 8347 40003 8353
rect 39945 8313 39957 8347
rect 39991 8344 40003 8347
rect 41230 8344 41236 8356
rect 39991 8316 41236 8344
rect 39991 8313 40003 8316
rect 39945 8307 40003 8313
rect 41230 8304 41236 8316
rect 41288 8304 41294 8356
rect 46842 8304 46848 8356
rect 46900 8304 46906 8356
rect 27890 8285 27896 8288
rect 27874 8279 27896 8285
rect 27874 8276 27886 8279
rect 27632 8248 27886 8276
rect 27874 8245 27886 8248
rect 27874 8239 27896 8245
rect 27890 8236 27896 8239
rect 27948 8236 27954 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 27801 8075 27859 8081
rect 27801 8041 27813 8075
rect 27847 8072 27859 8075
rect 27890 8072 27896 8084
rect 27847 8044 27896 8072
rect 27847 8041 27859 8044
rect 27801 8035 27859 8041
rect 27890 8032 27896 8044
rect 27948 8032 27954 8084
rect 28994 8032 29000 8084
rect 29052 8072 29058 8084
rect 29052 8044 31708 8072
rect 29052 8032 29058 8044
rect 31680 8016 31708 8044
rect 32306 8032 32312 8084
rect 32364 8032 32370 8084
rect 35158 8032 35164 8084
rect 35216 8072 35222 8084
rect 37553 8075 37611 8081
rect 37553 8072 37565 8075
rect 35216 8044 37565 8072
rect 35216 8032 35222 8044
rect 37553 8041 37565 8044
rect 37599 8041 37611 8075
rect 37553 8035 37611 8041
rect 40037 8075 40095 8081
rect 40037 8041 40049 8075
rect 40083 8072 40095 8075
rect 44174 8072 44180 8084
rect 40083 8044 44180 8072
rect 40083 8041 40095 8044
rect 40037 8035 40095 8041
rect 44174 8032 44180 8044
rect 44232 8032 44238 8084
rect 28261 8007 28319 8013
rect 28261 7973 28273 8007
rect 28307 8004 28319 8007
rect 30006 8004 30012 8016
rect 28307 7976 30012 8004
rect 28307 7973 28319 7976
rect 28261 7967 28319 7973
rect 30006 7964 30012 7976
rect 30064 7964 30070 8016
rect 31662 7964 31668 8016
rect 31720 8004 31726 8016
rect 34606 8004 34612 8016
rect 31720 7976 34612 8004
rect 31720 7964 31726 7976
rect 34606 7964 34612 7976
rect 34664 7964 34670 8016
rect 38381 8007 38439 8013
rect 38381 7973 38393 8007
rect 38427 8004 38439 8007
rect 45278 8004 45284 8016
rect 38427 7976 45284 8004
rect 38427 7973 38439 7976
rect 38381 7967 38439 7973
rect 45278 7964 45284 7976
rect 45336 7964 45342 8016
rect 25774 7896 25780 7948
rect 25832 7936 25838 7948
rect 26053 7939 26111 7945
rect 26053 7936 26065 7939
rect 25832 7908 26065 7936
rect 25832 7896 25838 7908
rect 26053 7905 26065 7908
rect 26099 7905 26111 7939
rect 26053 7899 26111 7905
rect 26329 7939 26387 7945
rect 26329 7905 26341 7939
rect 26375 7936 26387 7939
rect 27062 7936 27068 7948
rect 26375 7908 27068 7936
rect 26375 7905 26387 7908
rect 26329 7899 26387 7905
rect 27062 7896 27068 7908
rect 27120 7896 27126 7948
rect 28626 7896 28632 7948
rect 28684 7936 28690 7948
rect 28721 7939 28779 7945
rect 28721 7936 28733 7939
rect 28684 7908 28733 7936
rect 28684 7896 28690 7908
rect 28721 7905 28733 7908
rect 28767 7905 28779 7939
rect 28721 7899 28779 7905
rect 28905 7939 28963 7945
rect 28905 7905 28917 7939
rect 28951 7936 28963 7939
rect 31478 7936 31484 7948
rect 28951 7908 31484 7936
rect 28951 7905 28963 7908
rect 28905 7899 28963 7905
rect 31478 7896 31484 7908
rect 31536 7896 31542 7948
rect 31573 7939 31631 7945
rect 31573 7905 31585 7939
rect 31619 7936 31631 7939
rect 32582 7936 32588 7948
rect 31619 7908 32588 7936
rect 31619 7905 31631 7908
rect 31573 7899 31631 7905
rect 32582 7896 32588 7908
rect 32640 7896 32646 7948
rect 36081 7939 36139 7945
rect 36081 7905 36093 7939
rect 36127 7936 36139 7939
rect 37734 7936 37740 7948
rect 36127 7908 37740 7936
rect 36127 7905 36139 7908
rect 36081 7899 36139 7905
rect 37734 7896 37740 7908
rect 37792 7896 37798 7948
rect 28810 7828 28816 7880
rect 28868 7868 28874 7880
rect 31297 7871 31355 7877
rect 31297 7868 31309 7871
rect 28868 7840 31309 7868
rect 28868 7828 28874 7840
rect 31297 7837 31309 7840
rect 31343 7837 31355 7871
rect 31297 7831 31355 7837
rect 31389 7871 31447 7877
rect 31389 7837 31401 7871
rect 31435 7868 31447 7871
rect 31662 7868 31668 7880
rect 31435 7840 31668 7868
rect 31435 7837 31447 7840
rect 31389 7831 31447 7837
rect 31662 7828 31668 7840
rect 31720 7828 31726 7880
rect 32398 7828 32404 7880
rect 32456 7868 32462 7880
rect 32953 7871 33011 7877
rect 32953 7868 32965 7871
rect 32456 7840 32965 7868
rect 32456 7828 32462 7840
rect 32953 7837 32965 7840
rect 32999 7837 33011 7871
rect 32953 7831 33011 7837
rect 35253 7871 35311 7877
rect 35253 7837 35265 7871
rect 35299 7868 35311 7871
rect 35710 7868 35716 7880
rect 35299 7840 35716 7868
rect 35299 7837 35311 7840
rect 35253 7831 35311 7837
rect 35710 7828 35716 7840
rect 35768 7828 35774 7880
rect 35802 7828 35808 7880
rect 35860 7828 35866 7880
rect 37182 7828 37188 7880
rect 37240 7828 37246 7880
rect 38565 7871 38623 7877
rect 38565 7837 38577 7871
rect 38611 7837 38623 7871
rect 38565 7831 38623 7837
rect 26786 7760 26792 7812
rect 26844 7760 26850 7812
rect 35526 7800 35532 7812
rect 30944 7772 35532 7800
rect 23842 7692 23848 7744
rect 23900 7732 23906 7744
rect 30944 7741 30972 7772
rect 35526 7760 35532 7772
rect 35584 7760 35590 7812
rect 28629 7735 28687 7741
rect 28629 7732 28641 7735
rect 23900 7704 28641 7732
rect 23900 7692 23906 7704
rect 28629 7701 28641 7704
rect 28675 7701 28687 7735
rect 28629 7695 28687 7701
rect 30929 7735 30987 7741
rect 30929 7701 30941 7735
rect 30975 7701 30987 7735
rect 30929 7695 30987 7701
rect 33410 7692 33416 7744
rect 33468 7732 33474 7744
rect 38580 7732 38608 7831
rect 40218 7828 40224 7880
rect 40276 7828 40282 7880
rect 33468 7704 38608 7732
rect 33468 7692 33474 7704
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 34882 7528 34888 7540
rect 33152 7500 34888 7528
rect 28534 7420 28540 7472
rect 28592 7460 28598 7472
rect 28629 7463 28687 7469
rect 28629 7460 28641 7463
rect 28592 7432 28641 7460
rect 28592 7420 28598 7432
rect 28629 7429 28641 7432
rect 28675 7429 28687 7463
rect 28629 7423 28687 7429
rect 32490 7420 32496 7472
rect 32548 7420 32554 7472
rect 33152 7401 33180 7500
rect 34882 7488 34888 7500
rect 34940 7528 34946 7540
rect 35802 7528 35808 7540
rect 34940 7500 35808 7528
rect 34940 7488 34946 7500
rect 35802 7488 35808 7500
rect 35860 7488 35866 7540
rect 34698 7460 34704 7472
rect 34638 7432 34704 7460
rect 34698 7420 34704 7432
rect 34756 7460 34762 7472
rect 35250 7460 35256 7472
rect 34756 7432 35256 7460
rect 34756 7420 34762 7432
rect 35250 7420 35256 7432
rect 35308 7420 35314 7472
rect 35710 7420 35716 7472
rect 35768 7420 35774 7472
rect 46290 7420 46296 7472
rect 46348 7460 46354 7472
rect 46348 7432 47992 7460
rect 46348 7420 46354 7432
rect 33137 7395 33195 7401
rect 33137 7361 33149 7395
rect 33183 7361 33195 7395
rect 33137 7355 33195 7361
rect 35526 7352 35532 7404
rect 35584 7392 35590 7404
rect 35805 7395 35863 7401
rect 35805 7392 35817 7395
rect 35584 7364 35817 7392
rect 35584 7352 35590 7364
rect 35805 7361 35817 7364
rect 35851 7361 35863 7395
rect 35805 7355 35863 7361
rect 41230 7352 41236 7404
rect 41288 7392 41294 7404
rect 43257 7395 43315 7401
rect 43257 7392 43269 7395
rect 41288 7364 43269 7392
rect 41288 7352 41294 7364
rect 43257 7361 43269 7364
rect 43303 7361 43315 7395
rect 43257 7355 43315 7361
rect 45462 7352 45468 7404
rect 45520 7392 45526 7404
rect 47964 7401 47992 7432
rect 47121 7395 47179 7401
rect 47121 7392 47133 7395
rect 45520 7364 47133 7392
rect 45520 7352 45526 7364
rect 47121 7361 47133 7364
rect 47167 7361 47179 7395
rect 47121 7355 47179 7361
rect 47949 7395 48007 7401
rect 47949 7361 47961 7395
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 33413 7327 33471 7333
rect 33413 7293 33425 7327
rect 33459 7324 33471 7327
rect 34146 7324 34152 7336
rect 33459 7296 34152 7324
rect 33459 7293 33471 7296
rect 33413 7287 33471 7293
rect 34146 7284 34152 7296
rect 34204 7324 34210 7336
rect 34204 7296 34468 7324
rect 34204 7284 34210 7296
rect 28813 7259 28871 7265
rect 28813 7225 28825 7259
rect 28859 7256 28871 7259
rect 29270 7256 29276 7268
rect 28859 7228 29276 7256
rect 28859 7225 28871 7228
rect 28813 7219 28871 7225
rect 29270 7216 29276 7228
rect 29328 7216 29334 7268
rect 34440 7256 34468 7296
rect 34606 7284 34612 7336
rect 34664 7324 34670 7336
rect 34885 7327 34943 7333
rect 34885 7324 34897 7327
rect 34664 7296 34897 7324
rect 34664 7284 34670 7296
rect 34885 7293 34897 7296
rect 34931 7293 34943 7327
rect 35897 7327 35955 7333
rect 35897 7324 35909 7327
rect 34885 7287 34943 7293
rect 34992 7296 35909 7324
rect 34992 7256 35020 7296
rect 35897 7293 35909 7296
rect 35943 7293 35955 7327
rect 35897 7287 35955 7293
rect 49142 7284 49148 7336
rect 49200 7284 49206 7336
rect 34440 7228 35020 7256
rect 35345 7259 35403 7265
rect 35345 7225 35357 7259
rect 35391 7256 35403 7259
rect 40218 7256 40224 7268
rect 35391 7228 40224 7256
rect 35391 7225 35403 7228
rect 35345 7219 35403 7225
rect 40218 7216 40224 7228
rect 40276 7216 40282 7268
rect 32585 7191 32643 7197
rect 32585 7157 32597 7191
rect 32631 7188 32643 7191
rect 34422 7188 34428 7200
rect 32631 7160 34428 7188
rect 32631 7157 32643 7160
rect 32585 7151 32643 7157
rect 34422 7148 34428 7160
rect 34480 7148 34486 7200
rect 38473 7191 38531 7197
rect 38473 7157 38485 7191
rect 38519 7188 38531 7191
rect 39022 7188 39028 7200
rect 38519 7160 39028 7188
rect 38519 7157 38531 7160
rect 38473 7151 38531 7157
rect 39022 7148 39028 7160
rect 39080 7148 39086 7200
rect 43073 7191 43131 7197
rect 43073 7157 43085 7191
rect 43119 7188 43131 7191
rect 45462 7188 45468 7200
rect 43119 7160 45468 7188
rect 43119 7157 43131 7160
rect 43073 7151 43131 7157
rect 45462 7148 45468 7160
rect 45520 7148 45526 7200
rect 46934 7148 46940 7200
rect 46992 7148 46998 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 29996 6987 30054 6993
rect 29996 6953 30008 6987
rect 30042 6984 30054 6987
rect 31478 6984 31484 6996
rect 30042 6956 31484 6984
rect 30042 6953 30054 6956
rect 29996 6947 30054 6953
rect 31478 6944 31484 6956
rect 31536 6944 31542 6996
rect 36446 6944 36452 6996
rect 36504 6984 36510 6996
rect 36706 6987 36764 6993
rect 36706 6984 36718 6987
rect 36504 6956 36718 6984
rect 36504 6944 36510 6956
rect 36706 6953 36718 6956
rect 36752 6953 36764 6987
rect 36706 6947 36764 6953
rect 29730 6808 29736 6860
rect 29788 6848 29794 6860
rect 31941 6851 31999 6857
rect 31941 6848 31953 6851
rect 29788 6820 31953 6848
rect 29788 6808 29794 6820
rect 31941 6817 31953 6820
rect 31987 6848 31999 6851
rect 32306 6848 32312 6860
rect 31987 6820 32312 6848
rect 31987 6817 31999 6820
rect 31941 6811 31999 6817
rect 32306 6808 32312 6820
rect 32364 6848 32370 6860
rect 34054 6848 34060 6860
rect 32364 6820 34060 6848
rect 32364 6808 32370 6820
rect 34054 6808 34060 6820
rect 34112 6808 34118 6860
rect 35802 6808 35808 6860
rect 35860 6848 35866 6860
rect 36449 6851 36507 6857
rect 36449 6848 36461 6851
rect 35860 6820 36461 6848
rect 35860 6808 35866 6820
rect 36449 6817 36461 6820
rect 36495 6817 36507 6851
rect 36449 6811 36507 6817
rect 37734 6808 37740 6860
rect 37792 6848 37798 6860
rect 38197 6851 38255 6857
rect 38197 6848 38209 6851
rect 37792 6820 38209 6848
rect 37792 6808 37798 6820
rect 38197 6817 38209 6820
rect 38243 6848 38255 6851
rect 39209 6851 39267 6857
rect 39209 6848 39221 6851
rect 38243 6820 39221 6848
rect 38243 6817 38255 6820
rect 38197 6811 38255 6817
rect 39209 6817 39221 6820
rect 39255 6817 39267 6851
rect 39209 6811 39267 6817
rect 34238 6740 34244 6792
rect 34296 6780 34302 6792
rect 34977 6783 35035 6789
rect 34977 6780 34989 6783
rect 34296 6752 34989 6780
rect 34296 6740 34302 6752
rect 34977 6749 34989 6752
rect 35023 6749 35035 6783
rect 34977 6743 35035 6749
rect 35161 6783 35219 6789
rect 35161 6749 35173 6783
rect 35207 6780 35219 6783
rect 36354 6780 36360 6792
rect 35207 6752 36360 6780
rect 35207 6749 35219 6752
rect 35161 6743 35219 6749
rect 36354 6740 36360 6752
rect 36412 6740 36418 6792
rect 39022 6740 39028 6792
rect 39080 6740 39086 6792
rect 39114 6740 39120 6792
rect 39172 6740 39178 6792
rect 40034 6740 40040 6792
rect 40092 6780 40098 6792
rect 41693 6783 41751 6789
rect 41693 6780 41705 6783
rect 40092 6752 41705 6780
rect 40092 6740 40098 6752
rect 41693 6749 41705 6752
rect 41739 6749 41751 6783
rect 41693 6743 41751 6749
rect 47026 6740 47032 6792
rect 47084 6780 47090 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47084 6752 47961 6780
rect 47084 6740 47090 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 31386 6712 31392 6724
rect 31234 6684 31392 6712
rect 31386 6672 31392 6684
rect 31444 6672 31450 6724
rect 32214 6712 32220 6724
rect 31726 6684 32220 6712
rect 31481 6647 31539 6653
rect 31481 6613 31493 6647
rect 31527 6644 31539 6647
rect 31726 6644 31754 6684
rect 32214 6672 32220 6684
rect 32272 6672 32278 6724
rect 34698 6712 34704 6724
rect 33442 6684 34704 6712
rect 34698 6672 34704 6684
rect 34756 6672 34762 6724
rect 35618 6672 35624 6724
rect 35676 6712 35682 6724
rect 35805 6715 35863 6721
rect 35805 6712 35817 6715
rect 35676 6684 35817 6712
rect 35676 6672 35682 6684
rect 35805 6681 35817 6684
rect 35851 6681 35863 6715
rect 35805 6675 35863 6681
rect 37182 6672 37188 6724
rect 37240 6672 37246 6724
rect 38930 6712 38936 6724
rect 38580 6684 38936 6712
rect 31527 6616 31754 6644
rect 31527 6613 31539 6616
rect 31481 6607 31539 6613
rect 32582 6604 32588 6656
rect 32640 6644 32646 6656
rect 33689 6647 33747 6653
rect 33689 6644 33701 6647
rect 32640 6616 33701 6644
rect 32640 6604 32646 6616
rect 33689 6613 33701 6616
rect 33735 6613 33747 6647
rect 33689 6607 33747 6613
rect 35897 6647 35955 6653
rect 35897 6613 35909 6647
rect 35943 6644 35955 6647
rect 38580 6644 38608 6684
rect 38930 6672 38936 6684
rect 38988 6672 38994 6724
rect 49142 6672 49148 6724
rect 49200 6672 49206 6724
rect 35943 6616 38608 6644
rect 38657 6647 38715 6653
rect 35943 6613 35955 6616
rect 35897 6607 35955 6613
rect 38657 6613 38669 6647
rect 38703 6644 38715 6647
rect 40586 6644 40592 6656
rect 38703 6616 40592 6644
rect 38703 6613 38715 6616
rect 38657 6607 38715 6613
rect 40586 6604 40592 6616
rect 40644 6604 40650 6656
rect 41509 6647 41567 6653
rect 41509 6613 41521 6647
rect 41555 6644 41567 6647
rect 44082 6644 44088 6656
rect 41555 6616 44088 6644
rect 41555 6613 41567 6616
rect 41509 6607 41567 6613
rect 44082 6604 44088 6616
rect 44140 6604 44146 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 31386 6400 31392 6452
rect 31444 6440 31450 6452
rect 34057 6443 34115 6449
rect 31444 6412 33916 6440
rect 31444 6400 31450 6412
rect 32582 6332 32588 6384
rect 32640 6332 32646 6384
rect 33888 6372 33916 6412
rect 34057 6409 34069 6443
rect 34103 6440 34115 6443
rect 34146 6440 34152 6452
rect 34103 6412 34152 6440
rect 34103 6409 34115 6412
rect 34057 6403 34115 6409
rect 34146 6400 34152 6412
rect 34204 6400 34210 6452
rect 34698 6372 34704 6384
rect 33810 6344 34704 6372
rect 34698 6332 34704 6344
rect 34756 6332 34762 6384
rect 37550 6332 37556 6384
rect 37608 6332 37614 6384
rect 38286 6332 38292 6384
rect 38344 6332 38350 6384
rect 39482 6332 39488 6384
rect 39540 6332 39546 6384
rect 32306 6264 32312 6316
rect 32364 6264 32370 6316
rect 37182 6264 37188 6316
rect 37240 6304 37246 6316
rect 37240 6276 41414 6304
rect 37240 6264 37246 6276
rect 37737 6239 37795 6245
rect 37737 6205 37749 6239
rect 37783 6236 37795 6239
rect 40034 6236 40040 6248
rect 37783 6208 40040 6236
rect 37783 6205 37795 6208
rect 37737 6199 37795 6205
rect 40034 6196 40040 6208
rect 40092 6196 40098 6248
rect 41386 6236 41414 6276
rect 45186 6264 45192 6316
rect 45244 6304 45250 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 45244 6276 47961 6304
rect 45244 6264 45250 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 48498 6236 48504 6248
rect 41386 6208 48504 6236
rect 48498 6196 48504 6208
rect 48556 6196 48562 6248
rect 49145 6239 49203 6245
rect 49145 6205 49157 6239
rect 49191 6236 49203 6239
rect 49234 6236 49240 6248
rect 49191 6208 49240 6236
rect 49191 6205 49203 6208
rect 49145 6199 49203 6205
rect 49234 6196 49240 6208
rect 49292 6196 49298 6248
rect 38473 6171 38531 6177
rect 38473 6137 38485 6171
rect 38519 6168 38531 6171
rect 39482 6168 39488 6180
rect 38519 6140 39488 6168
rect 38519 6137 38531 6140
rect 38473 6131 38531 6137
rect 39482 6128 39488 6140
rect 39540 6128 39546 6180
rect 39577 6103 39635 6109
rect 39577 6069 39589 6103
rect 39623 6100 39635 6103
rect 42610 6100 42616 6112
rect 39623 6072 42616 6100
rect 39623 6069 39635 6072
rect 39577 6063 39635 6069
rect 42610 6060 42616 6072
rect 42668 6060 42674 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 32033 5899 32091 5905
rect 32033 5865 32045 5899
rect 32079 5896 32091 5899
rect 33410 5896 33416 5908
rect 32079 5868 33416 5896
rect 32079 5865 32091 5868
rect 32033 5859 32091 5865
rect 33410 5856 33416 5868
rect 33468 5856 33474 5908
rect 39025 5899 39083 5905
rect 39025 5865 39037 5899
rect 39071 5896 39083 5899
rect 40218 5896 40224 5908
rect 39071 5868 40224 5896
rect 39071 5865 39083 5868
rect 39025 5859 39083 5865
rect 40218 5856 40224 5868
rect 40276 5856 40282 5908
rect 45186 5856 45192 5908
rect 45244 5856 45250 5908
rect 40313 5831 40371 5837
rect 40313 5797 40325 5831
rect 40359 5828 40371 5831
rect 43346 5828 43352 5840
rect 40359 5800 43352 5828
rect 40359 5797 40371 5800
rect 40313 5791 40371 5797
rect 43346 5788 43352 5800
rect 43404 5788 43410 5840
rect 46842 5788 46848 5840
rect 46900 5788 46906 5840
rect 32214 5720 32220 5772
rect 32272 5760 32278 5772
rect 32585 5763 32643 5769
rect 32585 5760 32597 5763
rect 32272 5732 32597 5760
rect 32272 5720 32278 5732
rect 32585 5729 32597 5732
rect 32631 5729 32643 5763
rect 32585 5723 32643 5729
rect 38381 5763 38439 5769
rect 38381 5729 38393 5763
rect 38427 5760 38439 5763
rect 40126 5760 40132 5772
rect 38427 5732 40132 5760
rect 38427 5729 38439 5732
rect 38381 5723 38439 5729
rect 40126 5720 40132 5732
rect 40184 5720 40190 5772
rect 40402 5720 40408 5772
rect 40460 5760 40466 5772
rect 46860 5760 46888 5788
rect 40460 5732 45416 5760
rect 46860 5732 47992 5760
rect 40460 5720 40466 5732
rect 29178 5652 29184 5704
rect 29236 5692 29242 5704
rect 29825 5695 29883 5701
rect 29825 5692 29837 5695
rect 29236 5664 29837 5692
rect 29236 5652 29242 5664
rect 29825 5661 29837 5664
rect 29871 5661 29883 5695
rect 29825 5655 29883 5661
rect 32398 5652 32404 5704
rect 32456 5652 32462 5704
rect 37366 5652 37372 5704
rect 37424 5692 37430 5704
rect 38197 5695 38255 5701
rect 38197 5692 38209 5695
rect 37424 5664 38209 5692
rect 37424 5652 37430 5664
rect 38197 5661 38209 5664
rect 38243 5661 38255 5695
rect 38197 5655 38255 5661
rect 39206 5652 39212 5704
rect 39264 5692 39270 5704
rect 39264 5664 40264 5692
rect 39264 5652 39270 5664
rect 30006 5584 30012 5636
rect 30064 5624 30070 5636
rect 32493 5627 32551 5633
rect 32493 5624 32505 5627
rect 30064 5596 32505 5624
rect 30064 5584 30070 5596
rect 32493 5593 32505 5596
rect 32539 5593 32551 5627
rect 32493 5587 32551 5593
rect 36814 5584 36820 5636
rect 36872 5624 36878 5636
rect 38933 5627 38991 5633
rect 38933 5624 38945 5627
rect 36872 5596 38945 5624
rect 36872 5584 36878 5596
rect 38933 5593 38945 5596
rect 38979 5593 38991 5627
rect 38933 5587 38991 5593
rect 40129 5627 40187 5633
rect 40129 5593 40141 5627
rect 40175 5593 40187 5627
rect 40236 5624 40264 5664
rect 40586 5652 40592 5704
rect 40644 5692 40650 5704
rect 45388 5701 45416 5732
rect 42245 5695 42303 5701
rect 42245 5692 42257 5695
rect 40644 5664 42257 5692
rect 40644 5652 40650 5664
rect 42245 5661 42257 5664
rect 42291 5661 42303 5695
rect 42245 5655 42303 5661
rect 45373 5695 45431 5701
rect 45373 5661 45385 5695
rect 45419 5661 45431 5695
rect 45373 5655 45431 5661
rect 45462 5652 45468 5704
rect 45520 5692 45526 5704
rect 47964 5701 47992 5732
rect 46845 5695 46903 5701
rect 46845 5692 46857 5695
rect 45520 5664 46857 5692
rect 45520 5652 45526 5664
rect 46845 5661 46857 5664
rect 46891 5661 46903 5695
rect 46845 5655 46903 5661
rect 47949 5695 48007 5701
rect 47949 5661 47961 5695
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 40865 5627 40923 5633
rect 40865 5624 40877 5627
rect 40236 5596 40877 5624
rect 40129 5587 40187 5593
rect 40865 5593 40877 5596
rect 40911 5593 40923 5627
rect 40865 5587 40923 5593
rect 41049 5627 41107 5633
rect 41049 5593 41061 5627
rect 41095 5624 41107 5627
rect 42794 5624 42800 5636
rect 41095 5596 42800 5624
rect 41095 5593 41107 5596
rect 41049 5587 41107 5593
rect 27522 5516 27528 5568
rect 27580 5556 27586 5568
rect 29917 5559 29975 5565
rect 29917 5556 29929 5559
rect 27580 5528 29929 5556
rect 27580 5516 27586 5528
rect 29917 5525 29929 5528
rect 29963 5525 29975 5559
rect 40144 5556 40172 5587
rect 42794 5584 42800 5596
rect 42852 5584 42858 5636
rect 47026 5584 47032 5636
rect 47084 5584 47090 5636
rect 49142 5584 49148 5636
rect 49200 5584 49206 5636
rect 40494 5556 40500 5568
rect 40144 5528 40500 5556
rect 29917 5519 29975 5525
rect 40494 5516 40500 5528
rect 40552 5516 40558 5568
rect 42061 5559 42119 5565
rect 42061 5525 42073 5559
rect 42107 5556 42119 5559
rect 45462 5556 45468 5568
rect 42107 5528 45468 5556
rect 42107 5525 42119 5528
rect 42061 5519 42119 5525
rect 45462 5516 45468 5528
rect 45520 5516 45526 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 36630 5244 36636 5296
rect 36688 5284 36694 5296
rect 39945 5287 40003 5293
rect 39945 5284 39957 5287
rect 36688 5256 39957 5284
rect 36688 5244 36694 5256
rect 39945 5253 39957 5256
rect 39991 5253 40003 5287
rect 39945 5247 40003 5253
rect 40862 5244 40868 5296
rect 40920 5244 40926 5296
rect 44082 5176 44088 5228
rect 44140 5216 44146 5228
rect 46201 5219 46259 5225
rect 46201 5216 46213 5219
rect 44140 5188 46213 5216
rect 44140 5176 44146 5188
rect 46201 5185 46213 5188
rect 46247 5185 46259 5219
rect 46201 5179 46259 5185
rect 46934 5176 46940 5228
rect 46992 5216 46998 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 46992 5188 47961 5216
rect 46992 5176 46998 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 40129 5151 40187 5157
rect 40129 5117 40141 5151
rect 40175 5148 40187 5151
rect 47762 5148 47768 5160
rect 40175 5120 47768 5148
rect 40175 5117 40187 5120
rect 40129 5111 40187 5117
rect 47762 5108 47768 5120
rect 47820 5108 47826 5160
rect 49142 5108 49148 5160
rect 49200 5108 49206 5160
rect 41049 5083 41107 5089
rect 41049 5049 41061 5083
rect 41095 5080 41107 5083
rect 42702 5080 42708 5092
rect 41095 5052 42708 5080
rect 41095 5049 41107 5052
rect 41049 5043 41107 5049
rect 42702 5040 42708 5052
rect 42760 5040 42766 5092
rect 24670 4972 24676 5024
rect 24728 5012 24734 5024
rect 37642 5012 37648 5024
rect 24728 4984 37648 5012
rect 24728 4972 24734 4984
rect 37642 4972 37648 4984
rect 37700 4972 37706 5024
rect 46017 5015 46075 5021
rect 46017 4981 46029 5015
rect 46063 5012 46075 5015
rect 47946 5012 47952 5024
rect 46063 4984 47952 5012
rect 46063 4981 46075 4984
rect 46017 4975 46075 4981
rect 47946 4972 47952 4984
rect 48004 4972 48010 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 26878 4808 26884 4820
rect 10652 4780 26884 4808
rect 10652 4768 10658 4780
rect 26878 4768 26884 4780
rect 26936 4768 26942 4820
rect 31294 4768 31300 4820
rect 31352 4808 31358 4820
rect 46382 4808 46388 4820
rect 31352 4780 46388 4808
rect 31352 4768 31358 4780
rect 46382 4768 46388 4780
rect 46440 4768 46446 4820
rect 13446 4700 13452 4752
rect 13504 4740 13510 4752
rect 24026 4740 24032 4752
rect 13504 4712 24032 4740
rect 13504 4700 13510 4712
rect 24026 4700 24032 4712
rect 24084 4700 24090 4752
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11471 4644 16574 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 16546 4604 16574 4644
rect 47854 4632 47860 4684
rect 47912 4672 47918 4684
rect 48409 4675 48467 4681
rect 48409 4672 48421 4675
rect 47912 4644 48421 4672
rect 47912 4632 47918 4644
rect 48409 4641 48421 4644
rect 48455 4641 48467 4675
rect 48409 4635 48467 4641
rect 24762 4604 24768 4616
rect 12834 4576 14412 4604
rect 16546 4576 24768 4604
rect 11698 4496 11704 4548
rect 11756 4496 11762 4548
rect 13446 4496 13452 4548
rect 13504 4496 13510 4548
rect 14384 4536 14412 4576
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 46106 4564 46112 4616
rect 46164 4564 46170 4616
rect 47946 4564 47952 4616
rect 48004 4564 48010 4616
rect 26786 4536 26792 4548
rect 14384 4508 26792 4536
rect 26786 4496 26792 4508
rect 26844 4496 26850 4548
rect 47305 4539 47363 4545
rect 47305 4505 47317 4539
rect 47351 4536 47363 4539
rect 48682 4536 48688 4548
rect 47351 4508 48688 4536
rect 47351 4505 47363 4508
rect 47305 4499 47363 4505
rect 48682 4496 48688 4508
rect 48740 4496 48746 4548
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 34149 4131 34207 4137
rect 34149 4097 34161 4131
rect 34195 4128 34207 4131
rect 35342 4128 35348 4140
rect 34195 4100 35348 4128
rect 34195 4097 34207 4100
rect 34149 4091 34207 4097
rect 35342 4088 35348 4100
rect 35400 4088 35406 4140
rect 38930 4088 38936 4140
rect 38988 4128 38994 4140
rect 39117 4131 39175 4137
rect 39117 4128 39129 4131
rect 38988 4100 39129 4128
rect 38988 4088 38994 4100
rect 39117 4097 39129 4100
rect 39163 4097 39175 4131
rect 39117 4091 39175 4097
rect 42794 4088 42800 4140
rect 42852 4128 42858 4140
rect 44269 4131 44327 4137
rect 44269 4128 44281 4131
rect 42852 4100 44281 4128
rect 42852 4088 42858 4100
rect 44269 4097 44281 4100
rect 44315 4097 44327 4131
rect 44269 4091 44327 4097
rect 45462 4088 45468 4140
rect 45520 4128 45526 4140
rect 46477 4131 46535 4137
rect 46477 4128 46489 4131
rect 45520 4100 46489 4128
rect 45520 4088 45526 4100
rect 46477 4097 46489 4100
rect 46523 4097 46535 4131
rect 46477 4091 46535 4097
rect 47026 4088 47032 4140
rect 47084 4128 47090 4140
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 47084 4100 47961 4128
rect 47084 4088 47090 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 33870 4020 33876 4072
rect 33928 4060 33934 4072
rect 34425 4063 34483 4069
rect 34425 4060 34437 4063
rect 33928 4032 34437 4060
rect 33928 4020 33934 4032
rect 34425 4029 34437 4032
rect 34471 4029 34483 4063
rect 34425 4023 34483 4029
rect 39022 4020 39028 4072
rect 39080 4060 39086 4072
rect 39577 4063 39635 4069
rect 39577 4060 39589 4063
rect 39080 4032 39589 4060
rect 39080 4020 39086 4032
rect 39577 4029 39589 4032
rect 39623 4029 39635 4063
rect 39577 4023 39635 4029
rect 44174 4020 44180 4072
rect 44232 4060 44238 4072
rect 44729 4063 44787 4069
rect 44729 4060 44741 4063
rect 44232 4032 44741 4060
rect 44232 4020 44238 4032
rect 44729 4029 44741 4032
rect 44775 4029 44787 4063
rect 44729 4023 44787 4029
rect 49142 4020 49148 4072
rect 49200 4020 49206 4072
rect 46290 3884 46296 3936
rect 46348 3884 46354 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 32122 3720 32128 3732
rect 20956 3692 32128 3720
rect 20956 3680 20962 3692
rect 32122 3680 32128 3692
rect 32180 3680 32186 3732
rect 48498 3680 48504 3732
rect 48556 3680 48562 3732
rect 14366 3612 14372 3664
rect 14424 3652 14430 3664
rect 33318 3652 33324 3664
rect 14424 3624 28948 3652
rect 14424 3612 14430 3624
rect 20254 3544 20260 3596
rect 20312 3544 20318 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 25041 3587 25099 3593
rect 25041 3584 25053 3587
rect 24360 3556 25053 3584
rect 24360 3544 24366 3556
rect 25041 3553 25053 3556
rect 25087 3553 25099 3587
rect 25041 3547 25099 3553
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 17000 3488 17233 3516
rect 17000 3476 17006 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 19886 3476 19892 3528
rect 19944 3516 19950 3528
rect 19981 3519 20039 3525
rect 19981 3516 19993 3519
rect 19944 3488 19993 3516
rect 19944 3476 19950 3488
rect 19981 3485 19993 3488
rect 20027 3485 20039 3519
rect 19981 3479 20039 3485
rect 24670 3476 24676 3528
rect 24728 3476 24734 3528
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 23658 3448 23664 3460
rect 4028 3420 23664 3448
rect 4028 3408 4034 3420
rect 23658 3408 23664 3420
rect 23716 3408 23722 3460
rect 17037 3383 17095 3389
rect 17037 3349 17049 3383
rect 17083 3380 17095 3383
rect 28810 3380 28816 3392
rect 17083 3352 28816 3380
rect 17083 3349 17095 3352
rect 17037 3343 17095 3349
rect 28810 3340 28816 3352
rect 28868 3340 28874 3392
rect 28920 3380 28948 3624
rect 29932 3624 33324 3652
rect 29932 3525 29960 3624
rect 33318 3612 33324 3624
rect 33376 3612 33382 3664
rect 30193 3587 30251 3593
rect 30193 3553 30205 3587
rect 30239 3553 30251 3587
rect 30193 3547 30251 3553
rect 29917 3519 29975 3525
rect 29917 3485 29929 3519
rect 29963 3485 29975 3519
rect 29917 3479 29975 3485
rect 29454 3408 29460 3460
rect 29512 3448 29518 3460
rect 30208 3448 30236 3547
rect 30926 3544 30932 3596
rect 30984 3584 30990 3596
rect 32033 3587 32091 3593
rect 32033 3584 32045 3587
rect 30984 3556 32045 3584
rect 30984 3544 30990 3556
rect 32033 3553 32045 3556
rect 32079 3553 32091 3587
rect 32033 3547 32091 3553
rect 34606 3544 34612 3596
rect 34664 3584 34670 3596
rect 35345 3587 35403 3593
rect 35345 3584 35357 3587
rect 34664 3556 35357 3584
rect 34664 3544 34670 3556
rect 35345 3553 35357 3556
rect 35391 3553 35403 3587
rect 35345 3547 35403 3553
rect 36078 3544 36084 3596
rect 36136 3584 36142 3596
rect 37185 3587 37243 3593
rect 37185 3584 37197 3587
rect 36136 3556 37197 3584
rect 36136 3544 36142 3556
rect 37185 3553 37197 3556
rect 37231 3553 37243 3587
rect 37185 3547 37243 3553
rect 39758 3544 39764 3596
rect 39816 3584 39822 3596
rect 40497 3587 40555 3593
rect 40497 3584 40509 3587
rect 39816 3556 40509 3584
rect 39816 3544 39822 3556
rect 40497 3553 40509 3556
rect 40543 3553 40555 3587
rect 40497 3547 40555 3553
rect 41230 3544 41236 3596
rect 41288 3584 41294 3596
rect 42337 3587 42395 3593
rect 42337 3584 42349 3587
rect 41288 3556 42349 3584
rect 41288 3544 41294 3556
rect 42337 3553 42349 3556
rect 42383 3553 42395 3587
rect 42337 3547 42395 3553
rect 44910 3544 44916 3596
rect 44968 3584 44974 3596
rect 45649 3587 45707 3593
rect 45649 3584 45661 3587
rect 44968 3556 45661 3584
rect 44968 3544 44974 3556
rect 45649 3553 45661 3556
rect 45695 3553 45707 3587
rect 45649 3547 45707 3553
rect 31665 3519 31723 3525
rect 31665 3485 31677 3519
rect 31711 3485 31723 3519
rect 31665 3479 31723 3485
rect 29512 3420 30236 3448
rect 29512 3408 29518 3420
rect 30742 3380 30748 3392
rect 28920 3352 30748 3380
rect 30742 3340 30748 3352
rect 30800 3340 30806 3392
rect 31680 3380 31708 3479
rect 34422 3476 34428 3528
rect 34480 3516 34486 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34480 3488 34897 3516
rect 34480 3476 34486 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 36909 3519 36967 3525
rect 36909 3485 36921 3519
rect 36955 3516 36967 3519
rect 38562 3516 38568 3528
rect 36955 3488 38568 3516
rect 36955 3485 36967 3488
rect 36909 3479 36967 3485
rect 38562 3476 38568 3488
rect 38620 3476 38626 3528
rect 40034 3476 40040 3528
rect 40092 3476 40098 3528
rect 40126 3476 40132 3528
rect 40184 3516 40190 3528
rect 41877 3519 41935 3525
rect 41877 3516 41889 3519
rect 40184 3488 41889 3516
rect 40184 3476 40190 3488
rect 41877 3485 41889 3488
rect 41923 3485 41935 3519
rect 41877 3479 41935 3485
rect 42702 3476 42708 3528
rect 42760 3516 42766 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 42760 3488 45201 3516
rect 42760 3476 42766 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 47118 3408 47124 3460
rect 47176 3448 47182 3460
rect 47213 3451 47271 3457
rect 47213 3448 47225 3451
rect 47176 3420 47225 3448
rect 47176 3408 47182 3420
rect 47213 3417 47225 3420
rect 47259 3417 47271 3451
rect 47213 3411 47271 3417
rect 35986 3380 35992 3392
rect 31680 3352 35992 3380
rect 35986 3340 35992 3352
rect 36044 3340 36050 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 3970 3136 3976 3188
rect 4028 3136 4034 3188
rect 6733 3179 6791 3185
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 11701 3179 11759 3185
rect 6779 3148 6914 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 6886 3108 6914 3148
rect 11701 3145 11713 3179
rect 11747 3176 11759 3179
rect 22002 3176 22008 3188
rect 11747 3148 22008 3176
rect 11747 3145 11759 3148
rect 11701 3139 11759 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 33502 3176 33508 3188
rect 22480 3148 33508 3176
rect 18598 3108 18604 3120
rect 6886 3080 18604 3108
rect 18598 3068 18604 3080
rect 18656 3068 18662 3120
rect 2590 3000 2596 3052
rect 2648 3000 2654 3052
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3752 3012 3893 3040
rect 3752 3000 3758 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6696 3012 6929 3040
rect 6696 3000 6702 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8904 3012 9045 3040
rect 8904 3000 8910 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11885 3043 11943 3049
rect 11885 3040 11897 3043
rect 11112 3012 11897 3040
rect 11112 3000 11118 3012
rect 11885 3009 11897 3012
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3040 12955 3043
rect 13354 3040 13360 3052
rect 12943 3012 13360 3040
rect 12943 3009 12955 3012
rect 12897 3003 12955 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 22370 3040 22376 3052
rect 18095 3012 22376 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 22370 3000 22376 3012
rect 22428 3000 22434 3052
rect 22480 3049 22508 3148
rect 33502 3136 33508 3148
rect 33560 3136 33566 3188
rect 30558 3108 30564 3120
rect 24964 3080 30564 3108
rect 22465 3043 22523 3049
rect 22465 3009 22477 3043
rect 22511 3009 22523 3043
rect 22465 3003 22523 3009
rect 2222 2932 2228 2984
rect 2280 2972 2286 2984
rect 2317 2975 2375 2981
rect 2317 2972 2329 2975
rect 2280 2944 2329 2972
rect 2280 2932 2286 2944
rect 2317 2941 2329 2944
rect 2363 2941 2375 2975
rect 2317 2935 2375 2941
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 12621 2975 12679 2981
rect 12621 2972 12633 2975
rect 12584 2944 12633 2972
rect 12584 2932 12590 2944
rect 12621 2941 12633 2944
rect 12667 2941 12679 2975
rect 12621 2935 12679 2941
rect 13998 2932 14004 2984
rect 14056 2972 14062 2984
rect 14093 2975 14151 2981
rect 14093 2972 14105 2975
rect 14056 2944 14105 2972
rect 14056 2932 14062 2944
rect 14093 2941 14105 2944
rect 14139 2941 14151 2975
rect 14093 2935 14151 2941
rect 17678 2932 17684 2984
rect 17736 2972 17742 2984
rect 17773 2975 17831 2981
rect 17773 2972 17785 2975
rect 17736 2944 17785 2972
rect 17736 2932 17742 2944
rect 17773 2941 17785 2944
rect 17819 2941 17831 2975
rect 17773 2935 17831 2941
rect 19150 2932 19156 2984
rect 19208 2972 19214 2984
rect 19245 2975 19303 2981
rect 19245 2972 19257 2975
rect 19208 2944 19257 2972
rect 19208 2932 19214 2944
rect 19245 2941 19257 2944
rect 19291 2941 19303 2975
rect 19245 2935 19303 2941
rect 19521 2975 19579 2981
rect 19521 2941 19533 2975
rect 19567 2941 19579 2975
rect 19521 2935 19579 2941
rect 9217 2907 9275 2913
rect 9217 2873 9229 2907
rect 9263 2904 9275 2907
rect 19536 2904 19564 2935
rect 20622 2932 20628 2984
rect 20680 2932 20686 2984
rect 20898 2932 20904 2984
rect 20956 2932 20962 2984
rect 22094 2932 22100 2984
rect 22152 2972 22158 2984
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 22152 2944 22201 2972
rect 22152 2932 22158 2944
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 24964 2972 24992 3080
rect 30558 3068 30564 3080
rect 30616 3068 30622 3120
rect 44542 3108 44548 3120
rect 39500 3080 44548 3108
rect 25314 3000 25320 3052
rect 25372 3000 25378 3052
rect 27522 3000 27528 3052
rect 27580 3000 27586 3052
rect 29365 3043 29423 3049
rect 29365 3009 29377 3043
rect 29411 3040 29423 3043
rect 29546 3040 29552 3052
rect 29411 3012 29552 3040
rect 29411 3009 29423 3012
rect 29365 3003 29423 3009
rect 29546 3000 29552 3012
rect 29604 3000 29610 3052
rect 32493 3043 32551 3049
rect 32493 3009 32505 3043
rect 32539 3040 32551 3043
rect 33962 3040 33968 3052
rect 32539 3012 33968 3040
rect 32539 3009 32551 3012
rect 32493 3003 32551 3009
rect 33962 3000 33968 3012
rect 34020 3000 34026 3052
rect 34333 3043 34391 3049
rect 34333 3009 34345 3043
rect 34379 3040 34391 3043
rect 34974 3040 34980 3052
rect 34379 3012 34980 3040
rect 34379 3009 34391 3012
rect 34333 3003 34391 3009
rect 34974 3000 34980 3012
rect 35032 3000 35038 3052
rect 37645 3043 37703 3049
rect 37645 3009 37657 3043
rect 37691 3040 37703 3043
rect 38838 3040 38844 3052
rect 37691 3012 38844 3040
rect 37691 3009 37703 3012
rect 37645 3003 37703 3009
rect 38838 3000 38844 3012
rect 38896 3000 38902 3052
rect 39500 3049 39528 3080
rect 44542 3068 44548 3080
rect 44600 3068 44606 3120
rect 49142 3068 49148 3120
rect 49200 3068 49206 3120
rect 39485 3043 39543 3049
rect 39485 3009 39497 3043
rect 39531 3009 39543 3043
rect 39485 3003 39543 3009
rect 42610 3000 42616 3052
rect 42668 3000 42674 3052
rect 43346 3000 43352 3052
rect 43404 3040 43410 3052
rect 44453 3043 44511 3049
rect 44453 3040 44465 3043
rect 43404 3012 44465 3040
rect 43404 3000 43410 3012
rect 44453 3009 44465 3012
rect 44499 3009 44511 3043
rect 44453 3003 44511 3009
rect 46290 3000 46296 3052
rect 46348 3040 46354 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 46348 3012 47961 3040
rect 46348 3000 46354 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 22189 2935 22247 2941
rect 22296 2944 24992 2972
rect 22296 2904 22324 2944
rect 25038 2932 25044 2984
rect 25096 2972 25102 2984
rect 25593 2975 25651 2981
rect 25593 2972 25605 2975
rect 25096 2944 25605 2972
rect 25096 2932 25102 2944
rect 25593 2941 25605 2944
rect 25639 2941 25651 2975
rect 25593 2935 25651 2941
rect 27246 2932 27252 2984
rect 27304 2972 27310 2984
rect 27801 2975 27859 2981
rect 27801 2972 27813 2975
rect 27304 2944 27813 2972
rect 27304 2932 27310 2944
rect 27801 2941 27813 2944
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 29641 2975 29699 2981
rect 29641 2972 29653 2975
rect 28776 2944 29653 2972
rect 28776 2932 28782 2944
rect 29641 2941 29653 2944
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 31662 2932 31668 2984
rect 31720 2972 31726 2984
rect 32769 2975 32827 2981
rect 32769 2972 32781 2975
rect 31720 2944 32781 2972
rect 31720 2932 31726 2944
rect 32769 2941 32781 2944
rect 32815 2941 32827 2975
rect 32769 2935 32827 2941
rect 34609 2975 34667 2981
rect 34609 2941 34621 2975
rect 34655 2941 34667 2975
rect 34609 2935 34667 2941
rect 9263 2876 16574 2904
rect 19536 2876 22324 2904
rect 9263 2873 9275 2876
rect 9217 2867 9275 2873
rect 16546 2836 16574 2876
rect 22370 2864 22376 2916
rect 22428 2904 22434 2916
rect 31110 2904 31116 2916
rect 22428 2876 31116 2904
rect 22428 2864 22434 2876
rect 31110 2864 31116 2876
rect 31168 2864 31174 2916
rect 32398 2864 32404 2916
rect 32456 2904 32462 2916
rect 34624 2904 34652 2935
rect 36814 2932 36820 2984
rect 36872 2972 36878 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 36872 2944 37933 2972
rect 36872 2932 36878 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 39761 2975 39819 2981
rect 39761 2941 39773 2975
rect 39807 2941 39819 2975
rect 39761 2935 39819 2941
rect 32456 2876 34652 2904
rect 32456 2864 32462 2876
rect 37550 2864 37556 2916
rect 37608 2904 37614 2916
rect 39776 2904 39804 2935
rect 41966 2932 41972 2984
rect 42024 2972 42030 2984
rect 43073 2975 43131 2981
rect 43073 2972 43085 2975
rect 42024 2944 43085 2972
rect 42024 2932 42030 2944
rect 43073 2941 43085 2944
rect 43119 2941 43131 2975
rect 43073 2935 43131 2941
rect 44913 2975 44971 2981
rect 44913 2941 44925 2975
rect 44959 2941 44971 2975
rect 44913 2935 44971 2941
rect 37608 2876 39804 2904
rect 37608 2864 37614 2876
rect 42702 2864 42708 2916
rect 42760 2904 42766 2916
rect 44928 2904 44956 2935
rect 42760 2876 44956 2904
rect 42760 2864 42766 2876
rect 27798 2836 27804 2848
rect 16546 2808 27804 2836
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 28350 2796 28356 2848
rect 28408 2836 28414 2848
rect 30374 2836 30380 2848
rect 28408 2808 30380 2836
rect 28408 2796 28414 2808
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 45646 2796 45652 2848
rect 45704 2836 45710 2848
rect 48314 2836 48320 2848
rect 45704 2808 48320 2836
rect 45704 2796 45710 2808
rect 48314 2796 48320 2808
rect 48372 2796 48378 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 11698 2632 11704 2644
rect 1627 2604 11704 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 15059 2635 15117 2641
rect 15059 2601 15071 2635
rect 15105 2632 15117 2635
rect 30834 2632 30840 2644
rect 15105 2604 30840 2632
rect 15105 2601 15117 2604
rect 15059 2595 15117 2601
rect 30834 2592 30840 2604
rect 30892 2592 30898 2644
rect 45370 2632 45376 2644
rect 40144 2604 45376 2632
rect 19794 2564 19800 2576
rect 6886 2536 19800 2564
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 6886 2496 6914 2536
rect 19794 2524 19800 2536
rect 19852 2524 19858 2576
rect 22557 2567 22615 2573
rect 22557 2533 22569 2567
rect 22603 2533 22615 2567
rect 22557 2527 22615 2533
rect 2915 2468 6914 2496
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 10594 2456 10600 2508
rect 10652 2456 10658 2508
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2496 12955 2499
rect 13262 2496 13268 2508
rect 12943 2468 13268 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 18049 2499 18107 2505
rect 14660 2468 18000 2496
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1544 2400 1777 2428
rect 1544 2388 1550 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2958 2428 2964 2440
rect 2639 2400 2964 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 7374 2388 7380 2440
rect 7432 2428 7438 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7432 2400 7665 2428
rect 7432 2388 7438 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8527 2400 10272 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 4430 2320 4436 2372
rect 4488 2360 4494 2372
rect 4617 2363 4675 2369
rect 4617 2360 4629 2363
rect 4488 2332 4629 2360
rect 4488 2320 4494 2332
rect 4617 2329 4629 2332
rect 4663 2329 4675 2363
rect 4617 2323 4675 2329
rect 5166 2320 5172 2372
rect 5224 2360 5230 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5224 2332 5365 2360
rect 5224 2320 5230 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5353 2323 5411 2329
rect 5534 2320 5540 2372
rect 5592 2320 5598 2372
rect 5902 2320 5908 2372
rect 5960 2360 5966 2372
rect 6641 2363 6699 2369
rect 6641 2360 6653 2363
rect 5960 2332 6653 2360
rect 5960 2320 5966 2332
rect 6641 2329 6653 2332
rect 6687 2329 6699 2363
rect 6641 2323 6699 2329
rect 8294 2320 8300 2372
rect 8352 2320 8358 2372
rect 9582 2320 9588 2372
rect 9640 2360 9646 2372
rect 9677 2363 9735 2369
rect 9677 2360 9689 2363
rect 9640 2332 9689 2360
rect 9640 2320 9646 2332
rect 9677 2329 9689 2332
rect 9723 2329 9735 2363
rect 9677 2323 9735 2329
rect 9858 2320 9864 2372
rect 9916 2320 9922 2372
rect 10244 2360 10272 2400
rect 10318 2388 10324 2440
rect 10376 2388 10382 2440
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 11848 2400 12081 2428
rect 11848 2388 11854 2400
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 14660 2428 14688 2468
rect 13219 2400 14688 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14792 2400 14841 2428
rect 14792 2388 14798 2400
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 16301 2431 16359 2437
rect 16301 2428 16313 2431
rect 15528 2400 16313 2428
rect 15528 2388 15534 2400
rect 16301 2397 16313 2400
rect 16347 2397 16359 2431
rect 16301 2391 16359 2397
rect 16482 2388 16488 2440
rect 16540 2428 16546 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16540 2400 17049 2428
rect 16540 2388 16546 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17972 2428 18000 2468
rect 18049 2465 18061 2499
rect 18095 2496 18107 2499
rect 18414 2496 18420 2508
rect 18095 2468 18420 2496
rect 18095 2465 18107 2468
rect 18049 2459 18107 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 22572 2496 22600 2527
rect 24578 2524 24584 2576
rect 24636 2564 24642 2576
rect 28994 2564 29000 2576
rect 24636 2536 29000 2564
rect 24636 2524 24642 2536
rect 28994 2524 29000 2536
rect 29052 2524 29058 2576
rect 33594 2564 33600 2576
rect 29196 2536 33600 2564
rect 22572 2468 24992 2496
rect 19978 2428 19984 2440
rect 17972 2400 19984 2428
rect 17037 2391 17095 2397
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 22741 2431 22799 2437
rect 22741 2397 22753 2431
rect 22787 2428 22799 2431
rect 22830 2428 22836 2440
rect 22787 2400 22836 2428
rect 22787 2397 22799 2400
rect 22741 2391 22799 2397
rect 22830 2388 22836 2400
rect 22888 2388 22894 2440
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2428 23259 2431
rect 23566 2428 23572 2440
rect 23247 2400 23572 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 23566 2388 23572 2400
rect 23624 2388 23630 2440
rect 24412 2400 24900 2428
rect 21174 2360 21180 2372
rect 10244 2332 21180 2360
rect 21174 2320 21180 2332
rect 21232 2320 21238 2372
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 21358 2360 21364 2372
rect 21315 2332 21364 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 21453 2363 21511 2369
rect 21453 2329 21465 2363
rect 21499 2360 21511 2363
rect 24412 2360 24440 2400
rect 21499 2332 24440 2360
rect 21499 2329 21511 2332
rect 21453 2323 21511 2329
rect 4706 2252 4712 2304
rect 4764 2252 4770 2304
rect 6730 2252 6736 2304
rect 6788 2252 6794 2304
rect 7466 2252 7472 2304
rect 7524 2252 7530 2304
rect 11882 2252 11888 2304
rect 11940 2252 11946 2304
rect 16114 2252 16120 2304
rect 16172 2252 16178 2304
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 17310 2292 17316 2304
rect 16899 2264 17316 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 18279 2295 18337 2301
rect 18279 2261 18291 2295
rect 18325 2292 18337 2295
rect 22278 2292 22284 2304
rect 18325 2264 22284 2292
rect 18325 2261 18337 2264
rect 18279 2255 18337 2261
rect 22278 2252 22284 2264
rect 22336 2252 22342 2304
rect 23431 2295 23489 2301
rect 23431 2261 23443 2295
rect 23477 2292 23489 2295
rect 24578 2292 24584 2304
rect 23477 2264 24584 2292
rect 23477 2261 23489 2264
rect 23431 2255 23489 2261
rect 24578 2252 24584 2264
rect 24636 2252 24642 2304
rect 24872 2292 24900 2400
rect 24964 2360 24992 2468
rect 25774 2456 25780 2508
rect 25832 2456 25838 2508
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26568 2468 27629 2496
rect 26568 2456 26574 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 27341 2431 27399 2437
rect 27341 2397 27353 2431
rect 27387 2428 27399 2431
rect 29196 2428 29224 2536
rect 33594 2524 33600 2536
rect 33652 2524 33658 2576
rect 30374 2456 30380 2508
rect 30432 2456 30438 2508
rect 32769 2499 32827 2505
rect 32769 2496 32781 2499
rect 30484 2468 32781 2496
rect 27387 2400 29224 2428
rect 27387 2397 27399 2400
rect 27341 2391 27399 2397
rect 29270 2388 29276 2440
rect 29328 2428 29334 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29328 2400 29745 2428
rect 29328 2388 29334 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30190 2388 30196 2440
rect 30248 2428 30254 2440
rect 30484 2428 30512 2468
rect 32769 2465 32781 2468
rect 32815 2465 32827 2499
rect 32769 2459 32827 2465
rect 35342 2456 35348 2508
rect 35400 2496 35406 2508
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 35400 2468 37933 2496
rect 35400 2456 35406 2468
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 30248 2400 30512 2428
rect 32493 2431 32551 2437
rect 30248 2388 30254 2400
rect 32493 2397 32505 2431
rect 32539 2428 32551 2431
rect 33778 2428 33784 2440
rect 32539 2400 33784 2428
rect 32539 2397 32551 2400
rect 32493 2391 32551 2397
rect 33778 2388 33784 2400
rect 33836 2388 33842 2440
rect 35069 2431 35127 2437
rect 35069 2397 35081 2431
rect 35115 2428 35127 2431
rect 36262 2428 36268 2440
rect 35115 2400 36268 2428
rect 35115 2397 35127 2400
rect 35069 2391 35127 2397
rect 36262 2388 36268 2400
rect 36320 2388 36326 2440
rect 36354 2388 36360 2440
rect 36412 2428 36418 2440
rect 40144 2437 40172 2604
rect 45370 2592 45376 2604
rect 45428 2592 45434 2644
rect 40218 2524 40224 2576
rect 40276 2564 40282 2576
rect 40276 2536 43208 2564
rect 40276 2524 40282 2536
rect 40586 2456 40592 2508
rect 40644 2496 40650 2508
rect 43073 2499 43131 2505
rect 43073 2496 43085 2499
rect 40644 2468 43085 2496
rect 40644 2456 40650 2468
rect 43073 2465 43085 2468
rect 43119 2465 43131 2499
rect 43073 2459 43131 2465
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 36412 2400 37473 2428
rect 36412 2388 36418 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 40129 2431 40187 2437
rect 40129 2397 40141 2431
rect 40175 2397 40187 2431
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 40129 2391 40187 2397
rect 40420 2400 42625 2428
rect 30650 2360 30656 2372
rect 24964 2332 30656 2360
rect 30650 2320 30656 2332
rect 30708 2320 30714 2372
rect 35805 2363 35863 2369
rect 35805 2329 35817 2363
rect 35851 2329 35863 2363
rect 35805 2323 35863 2329
rect 29362 2292 29368 2304
rect 24872 2264 29368 2292
rect 29362 2252 29368 2264
rect 29420 2252 29426 2304
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 35820 2292 35848 2323
rect 39482 2320 39488 2372
rect 39540 2360 39546 2372
rect 40420 2360 40448 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 43180 2428 43208 2536
rect 43438 2456 43444 2508
rect 43496 2496 43502 2508
rect 45649 2499 45707 2505
rect 45649 2496 45661 2499
rect 43496 2468 45661 2496
rect 43496 2456 43502 2468
rect 45649 2465 45661 2468
rect 45695 2465 45707 2499
rect 45649 2459 45707 2465
rect 48314 2456 48320 2508
rect 48372 2456 48378 2508
rect 45189 2431 45247 2437
rect 45189 2428 45201 2431
rect 43180 2400 45201 2428
rect 42613 2391 42671 2397
rect 45189 2397 45201 2400
rect 45235 2397 45247 2431
rect 45189 2391 45247 2397
rect 47762 2388 47768 2440
rect 47820 2388 47826 2440
rect 39540 2332 40448 2360
rect 40957 2363 41015 2369
rect 39540 2320 39546 2332
rect 40957 2329 40969 2363
rect 41003 2329 41015 2363
rect 40957 2323 41015 2329
rect 33192 2264 35848 2292
rect 33192 2252 33198 2264
rect 38286 2252 38292 2304
rect 38344 2292 38350 2304
rect 40972 2292 41000 2323
rect 38344 2264 41000 2292
rect 38344 2252 38350 2264
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
rect 7466 2048 7472 2100
rect 7524 2088 7530 2100
rect 17218 2088 17224 2100
rect 7524 2060 17224 2088
rect 7524 2048 7530 2060
rect 17218 2048 17224 2060
rect 17276 2048 17282 2100
rect 17310 2048 17316 2100
rect 17368 2088 17374 2100
rect 23842 2088 23848 2100
rect 17368 2060 23848 2088
rect 17368 2048 17374 2060
rect 23842 2048 23848 2060
rect 23900 2048 23906 2100
rect 3418 1980 3424 2032
rect 3476 2020 3482 2032
rect 41598 2020 41604 2032
rect 3476 1992 41604 2020
rect 3476 1980 3482 1992
rect 41598 1980 41604 1992
rect 41656 1980 41662 2032
rect 4706 1912 4712 1964
rect 4764 1952 4770 1964
rect 17218 1952 17224 1964
rect 4764 1924 17224 1952
rect 4764 1912 4770 1924
rect 17218 1912 17224 1924
rect 17276 1912 17282 1964
rect 17328 1924 18644 1952
rect 5534 1844 5540 1896
rect 5592 1884 5598 1896
rect 17328 1884 17356 1924
rect 18506 1884 18512 1896
rect 5592 1856 17356 1884
rect 17420 1856 18512 1884
rect 5592 1844 5598 1856
rect 11882 1776 11888 1828
rect 11940 1816 11946 1828
rect 17420 1816 17448 1856
rect 18506 1844 18512 1856
rect 18564 1844 18570 1896
rect 18616 1884 18644 1924
rect 21174 1912 21180 1964
rect 21232 1952 21238 1964
rect 27706 1952 27712 1964
rect 21232 1924 27712 1952
rect 21232 1912 21238 1924
rect 27706 1912 27712 1924
rect 27764 1912 27770 1964
rect 24946 1884 24952 1896
rect 18616 1856 24952 1884
rect 24946 1844 24952 1856
rect 25004 1844 25010 1896
rect 11940 1788 17448 1816
rect 11940 1776 11946 1788
rect 22278 1776 22284 1828
rect 22336 1816 22342 1828
rect 31570 1816 31576 1828
rect 22336 1788 31576 1816
rect 22336 1776 22342 1788
rect 31570 1776 31576 1788
rect 31628 1776 31634 1828
rect 16114 1708 16120 1760
rect 16172 1748 16178 1760
rect 26234 1748 26240 1760
rect 16172 1720 26240 1748
rect 16172 1708 16178 1720
rect 26234 1708 26240 1720
rect 26292 1708 26298 1760
rect 17218 1640 17224 1692
rect 17276 1680 17282 1692
rect 25682 1680 25688 1692
rect 17276 1652 25688 1680
rect 17276 1640 17282 1652
rect 25682 1640 25688 1652
rect 25740 1640 25746 1692
rect 6730 1504 6736 1556
rect 6788 1544 6794 1556
rect 23382 1544 23388 1556
rect 6788 1516 23388 1544
rect 6788 1504 6794 1516
rect 23382 1504 23388 1516
rect 23440 1504 23446 1556
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 27950 54374 28002 54426
rect 28014 54374 28066 54426
rect 28078 54374 28130 54426
rect 28142 54374 28194 54426
rect 28206 54374 28258 54426
rect 37950 54374 38002 54426
rect 38014 54374 38066 54426
rect 38078 54374 38130 54426
rect 38142 54374 38194 54426
rect 38206 54374 38258 54426
rect 47950 54374 48002 54426
rect 48014 54374 48066 54426
rect 48078 54374 48130 54426
rect 48142 54374 48194 54426
rect 48206 54374 48258 54426
rect 29552 54272 29604 54324
rect 8392 54204 8444 54256
rect 36084 54204 36136 54256
rect 46756 54204 46808 54256
rect 1400 54068 1452 54120
rect 7104 54136 7156 54188
rect 9588 54179 9640 54188
rect 9588 54145 9597 54179
rect 9597 54145 9631 54179
rect 9631 54145 9640 54179
rect 9588 54136 9640 54145
rect 12256 54179 12308 54188
rect 12256 54145 12265 54179
rect 12265 54145 12299 54179
rect 12299 54145 12308 54179
rect 12256 54136 12308 54145
rect 15016 54179 15068 54188
rect 15016 54145 15025 54179
rect 15025 54145 15059 54179
rect 15059 54145 15068 54179
rect 15016 54136 15068 54145
rect 17684 54179 17736 54188
rect 17684 54145 17693 54179
rect 17693 54145 17727 54179
rect 17727 54145 17736 54179
rect 17684 54136 17736 54145
rect 20260 54179 20312 54188
rect 20260 54145 20269 54179
rect 20269 54145 20303 54179
rect 20303 54145 20312 54179
rect 20260 54136 20312 54145
rect 22836 54179 22888 54188
rect 22836 54145 22845 54179
rect 22845 54145 22879 54179
rect 22879 54145 22888 54179
rect 22836 54136 22888 54145
rect 25412 54136 25464 54188
rect 28356 54179 28408 54188
rect 28356 54145 28365 54179
rect 28365 54145 28399 54179
rect 28399 54145 28408 54179
rect 28356 54136 28408 54145
rect 30748 54136 30800 54188
rect 33416 54136 33468 54188
rect 38752 54136 38804 54188
rect 41420 54136 41472 54188
rect 44088 54136 44140 54188
rect 48320 54179 48372 54188
rect 48320 54145 48329 54179
rect 48329 54145 48363 54179
rect 48363 54145 48372 54179
rect 48320 54136 48372 54145
rect 49056 54179 49108 54188
rect 49056 54145 49065 54179
rect 49065 54145 49099 54179
rect 49099 54145 49108 54179
rect 49056 54136 49108 54145
rect 4068 54068 4120 54120
rect 7012 54068 7064 54120
rect 9404 54068 9456 54120
rect 12348 54068 12400 54120
rect 14740 54068 14792 54120
rect 17868 54068 17920 54120
rect 20168 54068 20220 54120
rect 22744 54068 22796 54120
rect 15200 54000 15252 54052
rect 20536 53932 20588 53984
rect 24400 53932 24452 53984
rect 25688 53932 25740 53984
rect 30840 53975 30892 53984
rect 30840 53941 30849 53975
rect 30849 53941 30883 53975
rect 30883 53941 30892 53975
rect 30840 53932 30892 53941
rect 39028 53975 39080 53984
rect 39028 53941 39037 53975
rect 39037 53941 39071 53975
rect 39071 53941 39080 53975
rect 39028 53932 39080 53941
rect 41696 53975 41748 53984
rect 41696 53941 41705 53975
rect 41705 53941 41739 53975
rect 41739 53941 41748 53975
rect 41696 53932 41748 53941
rect 44364 53975 44416 53984
rect 44364 53941 44373 53975
rect 44373 53941 44407 53975
rect 44407 53941 44416 53975
rect 44364 53932 44416 53941
rect 46940 53975 46992 53984
rect 46940 53941 46949 53975
rect 46949 53941 46983 53975
rect 46983 53941 46992 53975
rect 46940 53932 46992 53941
rect 48504 53975 48556 53984
rect 48504 53941 48513 53975
rect 48513 53941 48547 53975
rect 48547 53941 48556 53975
rect 48504 53932 48556 53941
rect 48872 53932 48924 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 32950 53830 33002 53882
rect 33014 53830 33066 53882
rect 33078 53830 33130 53882
rect 33142 53830 33194 53882
rect 33206 53830 33258 53882
rect 42950 53830 43002 53882
rect 43014 53830 43066 53882
rect 43078 53830 43130 53882
rect 43142 53830 43194 53882
rect 43206 53830 43258 53882
rect 49424 53592 49476 53644
rect 48412 53524 48464 53576
rect 49148 53524 49200 53576
rect 43444 53388 43496 53440
rect 48412 53388 48464 53440
rect 50160 53388 50212 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 27950 53286 28002 53338
rect 28014 53286 28066 53338
rect 28078 53286 28130 53338
rect 28142 53286 28194 53338
rect 28206 53286 28258 53338
rect 37950 53286 38002 53338
rect 38014 53286 38066 53338
rect 38078 53286 38130 53338
rect 38142 53286 38194 53338
rect 38206 53286 38258 53338
rect 47950 53286 48002 53338
rect 48014 53286 48066 53338
rect 48078 53286 48130 53338
rect 48142 53286 48194 53338
rect 48206 53286 48258 53338
rect 8392 53184 8444 53236
rect 13728 53048 13780 53100
rect 49056 53091 49108 53100
rect 49056 53057 49065 53091
rect 49065 53057 49099 53091
rect 49099 53057 49108 53091
rect 49056 53048 49108 53057
rect 34704 52844 34756 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 32950 52742 33002 52794
rect 33014 52742 33066 52794
rect 33078 52742 33130 52794
rect 33142 52742 33194 52794
rect 33206 52742 33258 52794
rect 42950 52742 43002 52794
rect 43014 52742 43066 52794
rect 43078 52742 43130 52794
rect 43142 52742 43194 52794
rect 43206 52742 43258 52794
rect 49976 52436 50028 52488
rect 48964 52411 49016 52420
rect 48964 52377 48973 52411
rect 48973 52377 49007 52411
rect 49007 52377 49016 52411
rect 48964 52368 49016 52377
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 27950 52198 28002 52250
rect 28014 52198 28066 52250
rect 28078 52198 28130 52250
rect 28142 52198 28194 52250
rect 28206 52198 28258 52250
rect 37950 52198 38002 52250
rect 38014 52198 38066 52250
rect 38078 52198 38130 52250
rect 38142 52198 38194 52250
rect 38206 52198 38258 52250
rect 47950 52198 48002 52250
rect 48014 52198 48066 52250
rect 48078 52198 48130 52250
rect 48142 52198 48194 52250
rect 48206 52198 48258 52250
rect 7104 52096 7156 52148
rect 19800 51960 19852 52012
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 32950 51654 33002 51706
rect 33014 51654 33066 51706
rect 33078 51654 33130 51706
rect 33142 51654 33194 51706
rect 33206 51654 33258 51706
rect 42950 51654 43002 51706
rect 43014 51654 43066 51706
rect 43078 51654 43130 51706
rect 43142 51654 43194 51706
rect 43206 51654 43258 51706
rect 15016 51552 15068 51604
rect 12256 51484 12308 51536
rect 21640 51416 21692 51468
rect 17500 51348 17552 51400
rect 22744 51280 22796 51332
rect 48964 51323 49016 51332
rect 48964 51289 48973 51323
rect 48973 51289 49007 51323
rect 49007 51289 49016 51323
rect 48964 51280 49016 51289
rect 49608 51280 49660 51332
rect 9588 51212 9640 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 27950 51110 28002 51162
rect 28014 51110 28066 51162
rect 28078 51110 28130 51162
rect 28142 51110 28194 51162
rect 28206 51110 28258 51162
rect 37950 51110 38002 51162
rect 38014 51110 38066 51162
rect 38078 51110 38130 51162
rect 38142 51110 38194 51162
rect 38206 51110 38258 51162
rect 47950 51110 48002 51162
rect 48014 51110 48066 51162
rect 48078 51110 48130 51162
rect 48142 51110 48194 51162
rect 48206 51110 48258 51162
rect 48964 50915 49016 50924
rect 48964 50881 48973 50915
rect 48973 50881 49007 50915
rect 49007 50881 49016 50915
rect 48964 50872 49016 50881
rect 35716 50668 35768 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 32950 50566 33002 50618
rect 33014 50566 33066 50618
rect 33078 50566 33130 50618
rect 33142 50566 33194 50618
rect 33206 50566 33258 50618
rect 42950 50566 43002 50618
rect 43014 50566 43066 50618
rect 43078 50566 43130 50618
rect 43142 50566 43194 50618
rect 43206 50566 43258 50618
rect 15200 50464 15252 50516
rect 16120 50464 16172 50516
rect 17684 50464 17736 50516
rect 13728 50396 13780 50448
rect 17316 50396 17368 50448
rect 20536 50260 20588 50312
rect 20628 50192 20680 50244
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 27950 50022 28002 50074
rect 28014 50022 28066 50074
rect 28078 50022 28130 50074
rect 28142 50022 28194 50074
rect 28206 50022 28258 50074
rect 37950 50022 38002 50074
rect 38014 50022 38066 50074
rect 38078 50022 38130 50074
rect 38142 50022 38194 50074
rect 38206 50022 38258 50074
rect 47950 50022 48002 50074
rect 48014 50022 48066 50074
rect 48078 50022 48130 50074
rect 48142 50022 48194 50074
rect 48206 50022 48258 50074
rect 49148 49827 49200 49836
rect 49148 49793 49157 49827
rect 49157 49793 49191 49827
rect 49191 49793 49200 49827
rect 49148 49784 49200 49793
rect 49516 49716 49568 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 32950 49478 33002 49530
rect 33014 49478 33066 49530
rect 33078 49478 33130 49530
rect 33142 49478 33194 49530
rect 33206 49478 33258 49530
rect 42950 49478 43002 49530
rect 43014 49478 43066 49530
rect 43078 49478 43130 49530
rect 43142 49478 43194 49530
rect 43206 49478 43258 49530
rect 20260 49376 20312 49428
rect 22836 49376 22888 49428
rect 21456 49104 21508 49156
rect 23296 49104 23348 49156
rect 49148 49147 49200 49156
rect 49148 49113 49157 49147
rect 49157 49113 49191 49147
rect 49191 49113 49200 49147
rect 49148 49104 49200 49113
rect 50436 49104 50488 49156
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 27950 48934 28002 48986
rect 28014 48934 28066 48986
rect 28078 48934 28130 48986
rect 28142 48934 28194 48986
rect 28206 48934 28258 48986
rect 37950 48934 38002 48986
rect 38014 48934 38066 48986
rect 38078 48934 38130 48986
rect 38142 48934 38194 48986
rect 38206 48934 38258 48986
rect 47950 48934 48002 48986
rect 48014 48934 48066 48986
rect 48078 48934 48130 48986
rect 48142 48934 48194 48986
rect 48206 48934 48258 48986
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 32950 48390 33002 48442
rect 33014 48390 33066 48442
rect 33078 48390 33130 48442
rect 33142 48390 33194 48442
rect 33206 48390 33258 48442
rect 42950 48390 43002 48442
rect 43014 48390 43066 48442
rect 43078 48390 43130 48442
rect 43142 48390 43194 48442
rect 43206 48390 43258 48442
rect 16120 48263 16172 48272
rect 16120 48229 16129 48263
rect 16129 48229 16163 48263
rect 16163 48229 16172 48263
rect 16120 48220 16172 48229
rect 19432 48152 19484 48204
rect 18328 48016 18380 48068
rect 49148 48059 49200 48068
rect 49148 48025 49157 48059
rect 49157 48025 49191 48059
rect 49191 48025 49200 48059
rect 49148 48016 49200 48025
rect 19524 47948 19576 48000
rect 33692 47948 33744 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 27950 47846 28002 47898
rect 28014 47846 28066 47898
rect 28078 47846 28130 47898
rect 28142 47846 28194 47898
rect 28206 47846 28258 47898
rect 37950 47846 38002 47898
rect 38014 47846 38066 47898
rect 38078 47846 38130 47898
rect 38142 47846 38194 47898
rect 38206 47846 38258 47898
rect 47950 47846 48002 47898
rect 48014 47846 48066 47898
rect 48078 47846 48130 47898
rect 48142 47846 48194 47898
rect 48206 47846 48258 47898
rect 19800 47787 19852 47796
rect 19800 47753 19809 47787
rect 19809 47753 19843 47787
rect 19843 47753 19852 47787
rect 19800 47744 19852 47753
rect 20536 47676 20588 47728
rect 17316 47540 17368 47592
rect 49332 47651 49384 47660
rect 49332 47617 49341 47651
rect 49341 47617 49375 47651
rect 49375 47617 49384 47651
rect 49332 47608 49384 47617
rect 19524 47540 19576 47592
rect 21180 47540 21232 47592
rect 22008 47404 22060 47456
rect 46204 47404 46256 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 32950 47302 33002 47354
rect 33014 47302 33066 47354
rect 33078 47302 33130 47354
rect 33142 47302 33194 47354
rect 33206 47302 33258 47354
rect 42950 47302 43002 47354
rect 43014 47302 43066 47354
rect 43078 47302 43130 47354
rect 43142 47302 43194 47354
rect 43206 47302 43258 47354
rect 25688 47107 25740 47116
rect 25688 47073 25697 47107
rect 25697 47073 25731 47107
rect 25731 47073 25740 47107
rect 25688 47064 25740 47073
rect 19800 46996 19852 47048
rect 27528 46971 27580 46980
rect 27528 46937 27537 46971
rect 27537 46937 27571 46971
rect 27571 46937 27580 46971
rect 27528 46928 27580 46937
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 27950 46758 28002 46810
rect 28014 46758 28066 46810
rect 28078 46758 28130 46810
rect 28142 46758 28194 46810
rect 28206 46758 28258 46810
rect 37950 46758 38002 46810
rect 38014 46758 38066 46810
rect 38078 46758 38130 46810
rect 38142 46758 38194 46810
rect 38206 46758 38258 46810
rect 47950 46758 48002 46810
rect 48014 46758 48066 46810
rect 48078 46758 48130 46810
rect 48142 46758 48194 46810
rect 48206 46758 48258 46810
rect 20536 46656 20588 46708
rect 22468 46656 22520 46708
rect 24400 46588 24452 46640
rect 49332 46563 49384 46572
rect 49332 46529 49341 46563
rect 49341 46529 49375 46563
rect 49375 46529 49384 46563
rect 49332 46520 49384 46529
rect 22008 46452 22060 46504
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 41236 46316 41288 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 32950 46214 33002 46266
rect 33014 46214 33066 46266
rect 33078 46214 33130 46266
rect 33142 46214 33194 46266
rect 33206 46214 33258 46266
rect 42950 46214 43002 46266
rect 43014 46214 43066 46266
rect 43078 46214 43130 46266
rect 43142 46214 43194 46266
rect 43206 46214 43258 46266
rect 17500 46155 17552 46164
rect 17500 46121 17509 46155
rect 17509 46121 17543 46155
rect 17543 46121 17552 46155
rect 17500 46112 17552 46121
rect 21548 46112 21600 46164
rect 21640 46155 21692 46164
rect 21640 46121 21649 46155
rect 21649 46121 21683 46155
rect 21683 46121 21692 46155
rect 21640 46112 21692 46121
rect 20996 46044 21048 46096
rect 17316 46019 17368 46028
rect 17316 45985 17325 46019
rect 17325 45985 17359 46019
rect 17359 45985 17368 46019
rect 17316 45976 17368 45985
rect 17132 45951 17184 45960
rect 17132 45917 17141 45951
rect 17141 45917 17175 45951
rect 17175 45917 17184 45951
rect 17132 45908 17184 45917
rect 20536 45908 20588 45960
rect 30840 46044 30892 46096
rect 28908 46019 28960 46028
rect 28908 45985 28917 46019
rect 28917 45985 28951 46019
rect 28951 45985 28960 46019
rect 28908 45976 28960 45985
rect 49332 45951 49384 45960
rect 49332 45917 49341 45951
rect 49341 45917 49375 45951
rect 49375 45917 49384 45951
rect 49332 45908 49384 45917
rect 49884 45772 49936 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 27950 45670 28002 45722
rect 28014 45670 28066 45722
rect 28078 45670 28130 45722
rect 28142 45670 28194 45722
rect 28206 45670 28258 45722
rect 37950 45670 38002 45722
rect 38014 45670 38066 45722
rect 38078 45670 38130 45722
rect 38142 45670 38194 45722
rect 38206 45670 38258 45722
rect 47950 45670 48002 45722
rect 48014 45670 48066 45722
rect 48078 45670 48130 45722
rect 48142 45670 48194 45722
rect 48206 45670 48258 45722
rect 22836 45432 22888 45484
rect 29552 45475 29604 45484
rect 29552 45441 29561 45475
rect 29561 45441 29595 45475
rect 29595 45441 29604 45475
rect 29552 45432 29604 45441
rect 31392 45407 31444 45416
rect 31392 45373 31401 45407
rect 31401 45373 31435 45407
rect 31435 45373 31444 45407
rect 31392 45364 31444 45373
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 32950 45126 33002 45178
rect 33014 45126 33066 45178
rect 33078 45126 33130 45178
rect 33142 45126 33194 45178
rect 33206 45126 33258 45178
rect 42950 45126 43002 45178
rect 43014 45126 43066 45178
rect 43078 45126 43130 45178
rect 43142 45126 43194 45178
rect 43206 45126 43258 45178
rect 21180 45067 21232 45076
rect 21180 45033 21189 45067
rect 21189 45033 21223 45067
rect 21223 45033 21232 45067
rect 21180 45024 21232 45033
rect 21548 44888 21600 44940
rect 19432 44863 19484 44872
rect 19432 44829 19441 44863
rect 19441 44829 19475 44863
rect 19475 44829 19484 44863
rect 19432 44820 19484 44829
rect 49332 44863 49384 44872
rect 49332 44829 49341 44863
rect 49341 44829 49375 44863
rect 49375 44829 49384 44863
rect 49332 44820 49384 44829
rect 18328 44684 18380 44736
rect 23388 44752 23440 44804
rect 48688 44684 48740 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 27950 44582 28002 44634
rect 28014 44582 28066 44634
rect 28078 44582 28130 44634
rect 28142 44582 28194 44634
rect 28206 44582 28258 44634
rect 37950 44582 38002 44634
rect 38014 44582 38066 44634
rect 38078 44582 38130 44634
rect 38142 44582 38194 44634
rect 38206 44582 38258 44634
rect 47950 44582 48002 44634
rect 48014 44582 48066 44634
rect 48078 44582 48130 44634
rect 48142 44582 48194 44634
rect 48206 44582 48258 44634
rect 20628 44523 20680 44532
rect 20628 44489 20637 44523
rect 20637 44489 20671 44523
rect 20671 44489 20680 44523
rect 20628 44480 20680 44489
rect 22836 44480 22888 44532
rect 19800 44344 19852 44396
rect 22468 44387 22520 44396
rect 22468 44353 22477 44387
rect 22477 44353 22511 44387
rect 22511 44353 22520 44387
rect 22468 44344 22520 44353
rect 49148 44387 49200 44396
rect 49148 44353 49157 44387
rect 49157 44353 49191 44387
rect 49191 44353 49200 44387
rect 49148 44344 49200 44353
rect 19984 44319 20036 44328
rect 19984 44285 19993 44319
rect 19993 44285 20027 44319
rect 20027 44285 20036 44319
rect 19984 44276 20036 44285
rect 49700 44208 49752 44260
rect 22560 44183 22612 44192
rect 22560 44149 22569 44183
rect 22569 44149 22603 44183
rect 22603 44149 22612 44183
rect 22560 44140 22612 44149
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 32950 44038 33002 44090
rect 33014 44038 33066 44090
rect 33078 44038 33130 44090
rect 33142 44038 33194 44090
rect 33206 44038 33258 44090
rect 42950 44038 43002 44090
rect 43014 44038 43066 44090
rect 43078 44038 43130 44090
rect 43142 44038 43194 44090
rect 43206 44038 43258 44090
rect 43444 43800 43496 43852
rect 41420 43732 41472 43784
rect 42800 43664 42852 43716
rect 34980 43596 35032 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 27950 43494 28002 43546
rect 28014 43494 28066 43546
rect 28078 43494 28130 43546
rect 28142 43494 28194 43546
rect 28206 43494 28258 43546
rect 37950 43494 38002 43546
rect 38014 43494 38066 43546
rect 38078 43494 38130 43546
rect 38142 43494 38194 43546
rect 38206 43494 38258 43546
rect 47950 43494 48002 43546
rect 48014 43494 48066 43546
rect 48078 43494 48130 43546
rect 48142 43494 48194 43546
rect 48206 43494 48258 43546
rect 49148 43299 49200 43308
rect 49148 43265 49157 43299
rect 49157 43265 49191 43299
rect 49191 43265 49200 43299
rect 49148 43256 49200 43265
rect 49792 43120 49844 43172
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 32950 42950 33002 43002
rect 33014 42950 33066 43002
rect 33078 42950 33130 43002
rect 33142 42950 33194 43002
rect 33206 42950 33258 43002
rect 42950 42950 43002 43002
rect 43014 42950 43066 43002
rect 43078 42950 43130 43002
rect 43142 42950 43194 43002
rect 43206 42950 43258 43002
rect 49148 42619 49200 42628
rect 49148 42585 49157 42619
rect 49157 42585 49191 42619
rect 49191 42585 49200 42619
rect 49148 42576 49200 42585
rect 49240 42551 49292 42560
rect 49240 42517 49249 42551
rect 49249 42517 49283 42551
rect 49283 42517 49292 42551
rect 49240 42508 49292 42517
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 27950 42406 28002 42458
rect 28014 42406 28066 42458
rect 28078 42406 28130 42458
rect 28142 42406 28194 42458
rect 28206 42406 28258 42458
rect 37950 42406 38002 42458
rect 38014 42406 38066 42458
rect 38078 42406 38130 42458
rect 38142 42406 38194 42458
rect 38206 42406 38258 42458
rect 47950 42406 48002 42458
rect 48014 42406 48066 42458
rect 48078 42406 48130 42458
rect 48142 42406 48194 42458
rect 48206 42406 48258 42458
rect 21456 42347 21508 42356
rect 21456 42313 21465 42347
rect 21465 42313 21499 42347
rect 21499 42313 21508 42347
rect 21456 42304 21508 42313
rect 23296 42304 23348 42356
rect 20996 42211 21048 42220
rect 20996 42177 21005 42211
rect 21005 42177 21039 42211
rect 21039 42177 21048 42211
rect 20996 42168 21048 42177
rect 22652 42168 22704 42220
rect 20812 42143 20864 42152
rect 20812 42109 20821 42143
rect 20821 42109 20855 42143
rect 20855 42109 20864 42143
rect 20812 42100 20864 42109
rect 22836 42100 22888 42152
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 32950 41862 33002 41914
rect 33014 41862 33066 41914
rect 33078 41862 33130 41914
rect 33142 41862 33194 41914
rect 33206 41862 33258 41914
rect 42950 41862 43002 41914
rect 43014 41862 43066 41914
rect 43078 41862 43130 41914
rect 43142 41862 43194 41914
rect 43206 41862 43258 41914
rect 21548 41760 21600 41812
rect 19432 41624 19484 41676
rect 22836 41624 22888 41676
rect 23388 41624 23440 41676
rect 24308 41556 24360 41608
rect 22560 41420 22612 41472
rect 23388 41488 23440 41540
rect 49148 41531 49200 41540
rect 49148 41497 49157 41531
rect 49157 41497 49191 41531
rect 49191 41497 49200 41531
rect 49148 41488 49200 41497
rect 36820 41420 36872 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 27950 41318 28002 41370
rect 28014 41318 28066 41370
rect 28078 41318 28130 41370
rect 28142 41318 28194 41370
rect 28206 41318 28258 41370
rect 37950 41318 38002 41370
rect 38014 41318 38066 41370
rect 38078 41318 38130 41370
rect 38142 41318 38194 41370
rect 38206 41318 38258 41370
rect 47950 41318 48002 41370
rect 48014 41318 48066 41370
rect 48078 41318 48130 41370
rect 48142 41318 48194 41370
rect 48206 41318 48258 41370
rect 49332 41123 49384 41132
rect 49332 41089 49341 41123
rect 49341 41089 49375 41123
rect 49375 41089 49384 41123
rect 49332 41080 49384 41089
rect 48320 40876 48372 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 32950 40774 33002 40826
rect 33014 40774 33066 40826
rect 33078 40774 33130 40826
rect 33142 40774 33194 40826
rect 33206 40774 33258 40826
rect 42950 40774 43002 40826
rect 43014 40774 43066 40826
rect 43078 40774 43130 40826
rect 43142 40774 43194 40826
rect 43206 40774 43258 40826
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 27950 40230 28002 40282
rect 28014 40230 28066 40282
rect 28078 40230 28130 40282
rect 28142 40230 28194 40282
rect 28206 40230 28258 40282
rect 37950 40230 38002 40282
rect 38014 40230 38066 40282
rect 38078 40230 38130 40282
rect 38142 40230 38194 40282
rect 38206 40230 38258 40282
rect 47950 40230 48002 40282
rect 48014 40230 48066 40282
rect 48078 40230 48130 40282
rect 48142 40230 48194 40282
rect 48206 40230 48258 40282
rect 49056 40128 49108 40180
rect 49332 40035 49384 40044
rect 49332 40001 49341 40035
rect 49341 40001 49375 40035
rect 49375 40001 49384 40035
rect 49332 39992 49384 40001
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 32950 39686 33002 39738
rect 33014 39686 33066 39738
rect 33078 39686 33130 39738
rect 33142 39686 33194 39738
rect 33206 39686 33258 39738
rect 42950 39686 43002 39738
rect 43014 39686 43066 39738
rect 43078 39686 43130 39738
rect 43142 39686 43194 39738
rect 43206 39686 43258 39738
rect 49332 39423 49384 39432
rect 49332 39389 49341 39423
rect 49341 39389 49375 39423
rect 49375 39389 49384 39423
rect 49332 39380 49384 39389
rect 48596 39244 48648 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 27950 39142 28002 39194
rect 28014 39142 28066 39194
rect 28078 39142 28130 39194
rect 28142 39142 28194 39194
rect 28206 39142 28258 39194
rect 37950 39142 38002 39194
rect 38014 39142 38066 39194
rect 38078 39142 38130 39194
rect 38142 39142 38194 39194
rect 38206 39142 38258 39194
rect 47950 39142 48002 39194
rect 48014 39142 48066 39194
rect 48078 39142 48130 39194
rect 48142 39142 48194 39194
rect 48206 39142 48258 39194
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 32950 38598 33002 38650
rect 33014 38598 33066 38650
rect 33078 38598 33130 38650
rect 33142 38598 33194 38650
rect 33206 38598 33258 38650
rect 42950 38598 43002 38650
rect 43014 38598 43066 38650
rect 43078 38598 43130 38650
rect 43142 38598 43194 38650
rect 43206 38598 43258 38650
rect 49332 38335 49384 38344
rect 49332 38301 49341 38335
rect 49341 38301 49375 38335
rect 49375 38301 49384 38335
rect 49332 38292 49384 38301
rect 48964 38156 49016 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 27950 38054 28002 38106
rect 28014 38054 28066 38106
rect 28078 38054 28130 38106
rect 28142 38054 28194 38106
rect 28206 38054 28258 38106
rect 37950 38054 38002 38106
rect 38014 38054 38066 38106
rect 38078 38054 38130 38106
rect 38142 38054 38194 38106
rect 38206 38054 38258 38106
rect 47950 38054 48002 38106
rect 48014 38054 48066 38106
rect 48078 38054 48130 38106
rect 48142 38054 48194 38106
rect 48206 38054 48258 38106
rect 49148 37859 49200 37868
rect 49148 37825 49157 37859
rect 49157 37825 49191 37859
rect 49191 37825 49200 37859
rect 49148 37816 49200 37825
rect 50528 37680 50580 37732
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 32950 37510 33002 37562
rect 33014 37510 33066 37562
rect 33078 37510 33130 37562
rect 33142 37510 33194 37562
rect 33206 37510 33258 37562
rect 42950 37510 43002 37562
rect 43014 37510 43066 37562
rect 43078 37510 43130 37562
rect 43142 37510 43194 37562
rect 43206 37510 43258 37562
rect 22560 37204 22612 37256
rect 17132 37068 17184 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 27950 36966 28002 37018
rect 28014 36966 28066 37018
rect 28078 36966 28130 37018
rect 28142 36966 28194 37018
rect 28206 36966 28258 37018
rect 37950 36966 38002 37018
rect 38014 36966 38066 37018
rect 38078 36966 38130 37018
rect 38142 36966 38194 37018
rect 38206 36966 38258 37018
rect 47950 36966 48002 37018
rect 48014 36966 48066 37018
rect 48078 36966 48130 37018
rect 48142 36966 48194 37018
rect 48206 36966 48258 37018
rect 49148 36771 49200 36780
rect 49148 36737 49157 36771
rect 49157 36737 49191 36771
rect 49191 36737 49200 36771
rect 49148 36728 49200 36737
rect 48780 36524 48832 36576
rect 49424 36524 49476 36576
rect 49700 36524 49752 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 32950 36422 33002 36474
rect 33014 36422 33066 36474
rect 33078 36422 33130 36474
rect 33142 36422 33194 36474
rect 33206 36422 33258 36474
rect 42950 36422 43002 36474
rect 43014 36422 43066 36474
rect 43078 36422 43130 36474
rect 43142 36422 43194 36474
rect 43206 36422 43258 36474
rect 49332 36159 49384 36168
rect 49332 36125 49341 36159
rect 49341 36125 49375 36159
rect 49375 36125 49384 36159
rect 49332 36116 49384 36125
rect 49700 35980 49752 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 27950 35878 28002 35930
rect 28014 35878 28066 35930
rect 28078 35878 28130 35930
rect 28142 35878 28194 35930
rect 28206 35878 28258 35930
rect 37950 35878 38002 35930
rect 38014 35878 38066 35930
rect 38078 35878 38130 35930
rect 38142 35878 38194 35930
rect 38206 35878 38258 35930
rect 47950 35878 48002 35930
rect 48014 35878 48066 35930
rect 48078 35878 48130 35930
rect 48142 35878 48194 35930
rect 48206 35878 48258 35930
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 32950 35334 33002 35386
rect 33014 35334 33066 35386
rect 33078 35334 33130 35386
rect 33142 35334 33194 35386
rect 33206 35334 33258 35386
rect 42950 35334 43002 35386
rect 43014 35334 43066 35386
rect 43078 35334 43130 35386
rect 43142 35334 43194 35386
rect 43206 35334 43258 35386
rect 49332 35071 49384 35080
rect 49332 35037 49341 35071
rect 49341 35037 49375 35071
rect 49375 35037 49384 35071
rect 49332 35028 49384 35037
rect 50068 34892 50120 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 27950 34790 28002 34842
rect 28014 34790 28066 34842
rect 28078 34790 28130 34842
rect 28142 34790 28194 34842
rect 28206 34790 28258 34842
rect 37950 34790 38002 34842
rect 38014 34790 38066 34842
rect 38078 34790 38130 34842
rect 38142 34790 38194 34842
rect 38206 34790 38258 34842
rect 47950 34790 48002 34842
rect 48014 34790 48066 34842
rect 48078 34790 48130 34842
rect 48142 34790 48194 34842
rect 48206 34790 48258 34842
rect 23388 34688 23440 34740
rect 44180 34688 44232 34740
rect 24308 34552 24360 34604
rect 49332 34595 49384 34604
rect 49332 34561 49341 34595
rect 49341 34561 49375 34595
rect 49375 34561 49384 34595
rect 49332 34552 49384 34561
rect 22836 34484 22888 34536
rect 24216 34348 24268 34400
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 32950 34246 33002 34298
rect 33014 34246 33066 34298
rect 33078 34246 33130 34298
rect 33142 34246 33194 34298
rect 33206 34246 33258 34298
rect 42950 34246 43002 34298
rect 43014 34246 43066 34298
rect 43078 34246 43130 34298
rect 43142 34246 43194 34298
rect 43206 34246 43258 34298
rect 19984 34144 20036 34196
rect 38384 34076 38436 34128
rect 41236 34008 41288 34060
rect 22744 33940 22796 33992
rect 39672 33940 39724 33992
rect 27528 33804 27580 33856
rect 43720 34076 43772 34128
rect 42708 34051 42760 34060
rect 42708 34017 42717 34051
rect 42717 34017 42751 34051
rect 42751 34017 42760 34051
rect 42708 34008 42760 34017
rect 42892 34008 42944 34060
rect 49884 34008 49936 34060
rect 40960 33847 41012 33856
rect 40960 33813 40969 33847
rect 40969 33813 41003 33847
rect 41003 33813 41012 33847
rect 40960 33804 41012 33813
rect 41236 33804 41288 33856
rect 42892 33804 42944 33856
rect 43812 33804 43864 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 27950 33702 28002 33754
rect 28014 33702 28066 33754
rect 28078 33702 28130 33754
rect 28142 33702 28194 33754
rect 28206 33702 28258 33754
rect 37950 33702 38002 33754
rect 38014 33702 38066 33754
rect 38078 33702 38130 33754
rect 38142 33702 38194 33754
rect 38206 33702 38258 33754
rect 47950 33702 48002 33754
rect 48014 33702 48066 33754
rect 48078 33702 48130 33754
rect 48142 33702 48194 33754
rect 48206 33702 48258 33754
rect 48688 33600 48740 33652
rect 31392 33328 31444 33380
rect 43628 33464 43680 33516
rect 49332 33507 49384 33516
rect 49332 33473 49341 33507
rect 49341 33473 49375 33507
rect 49375 33473 49384 33507
rect 49332 33464 49384 33473
rect 43536 33396 43588 33448
rect 40224 33260 40276 33312
rect 43628 33260 43680 33312
rect 46848 33260 46900 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 32950 33158 33002 33210
rect 33014 33158 33066 33210
rect 33078 33158 33130 33210
rect 33142 33158 33194 33210
rect 33206 33158 33258 33210
rect 42950 33158 43002 33210
rect 43014 33158 43066 33210
rect 43078 33158 43130 33210
rect 43142 33158 43194 33210
rect 43206 33158 43258 33210
rect 49332 32895 49384 32904
rect 49332 32861 49341 32895
rect 49341 32861 49375 32895
rect 49375 32861 49384 32895
rect 49332 32852 49384 32861
rect 47400 32716 47452 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 27950 32614 28002 32666
rect 28014 32614 28066 32666
rect 28078 32614 28130 32666
rect 28142 32614 28194 32666
rect 28206 32614 28258 32666
rect 37950 32614 38002 32666
rect 38014 32614 38066 32666
rect 38078 32614 38130 32666
rect 38142 32614 38194 32666
rect 38206 32614 38258 32666
rect 47950 32614 48002 32666
rect 48014 32614 48066 32666
rect 48078 32614 48130 32666
rect 48142 32614 48194 32666
rect 48206 32614 48258 32666
rect 40132 32444 40184 32496
rect 41512 32444 41564 32496
rect 38476 32351 38528 32360
rect 38476 32317 38485 32351
rect 38485 32317 38519 32351
rect 38519 32317 38528 32351
rect 38476 32308 38528 32317
rect 41788 32308 41840 32360
rect 38292 32172 38344 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 32950 32070 33002 32122
rect 33014 32070 33066 32122
rect 33078 32070 33130 32122
rect 33142 32070 33194 32122
rect 33206 32070 33258 32122
rect 42950 32070 43002 32122
rect 43014 32070 43066 32122
rect 43078 32070 43130 32122
rect 43142 32070 43194 32122
rect 43206 32070 43258 32122
rect 24400 31832 24452 31884
rect 24768 31832 24820 31884
rect 42892 31968 42944 32020
rect 41788 31943 41840 31952
rect 41788 31909 41797 31943
rect 41797 31909 41831 31943
rect 41831 31909 41840 31943
rect 41788 31900 41840 31909
rect 41880 31900 41932 31952
rect 45652 31900 45704 31952
rect 40316 31875 40368 31884
rect 40316 31841 40325 31875
rect 40325 31841 40359 31875
rect 40359 31841 40368 31875
rect 40316 31832 40368 31841
rect 40040 31807 40092 31816
rect 40040 31773 40049 31807
rect 40049 31773 40083 31807
rect 40083 31773 40092 31807
rect 40040 31764 40092 31773
rect 41512 31832 41564 31884
rect 42708 31832 42760 31884
rect 43352 31832 43404 31884
rect 42892 31764 42944 31816
rect 48320 31764 48372 31816
rect 49332 31807 49384 31816
rect 49332 31773 49341 31807
rect 49341 31773 49375 31807
rect 49375 31773 49384 31807
rect 49332 31764 49384 31773
rect 34336 31628 34388 31680
rect 46940 31628 46992 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 27950 31526 28002 31578
rect 28014 31526 28066 31578
rect 28078 31526 28130 31578
rect 28142 31526 28194 31578
rect 28206 31526 28258 31578
rect 37950 31526 38002 31578
rect 38014 31526 38066 31578
rect 38078 31526 38130 31578
rect 38142 31526 38194 31578
rect 38206 31526 38258 31578
rect 47950 31526 48002 31578
rect 48014 31526 48066 31578
rect 48078 31526 48130 31578
rect 48142 31526 48194 31578
rect 48206 31526 48258 31578
rect 34336 31288 34388 31340
rect 35164 31288 35216 31340
rect 38476 31356 38528 31408
rect 40132 31356 40184 31408
rect 40040 31288 40092 31340
rect 41420 31424 41472 31476
rect 41512 31424 41564 31476
rect 43720 31467 43772 31476
rect 43720 31433 43729 31467
rect 43729 31433 43763 31467
rect 43763 31433 43772 31467
rect 43720 31424 43772 31433
rect 49056 31424 49108 31476
rect 42800 31356 42852 31408
rect 42892 31356 42944 31408
rect 43904 31356 43956 31408
rect 49332 31331 49384 31340
rect 49332 31297 49341 31331
rect 49341 31297 49375 31331
rect 49375 31297 49384 31331
rect 49332 31288 49384 31297
rect 34980 31220 35032 31272
rect 35624 31220 35676 31272
rect 38292 31220 38344 31272
rect 38568 31220 38620 31272
rect 43536 31220 43588 31272
rect 31484 31152 31536 31204
rect 42524 31152 42576 31204
rect 39672 31127 39724 31136
rect 39672 31093 39681 31127
rect 39681 31093 39715 31127
rect 39715 31093 39724 31127
rect 39672 31084 39724 31093
rect 40316 31084 40368 31136
rect 43444 31084 43496 31136
rect 48320 31084 48372 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 32950 30982 33002 31034
rect 33014 30982 33066 31034
rect 33078 30982 33130 31034
rect 33142 30982 33194 31034
rect 33206 30982 33258 31034
rect 42950 30982 43002 31034
rect 43014 30982 43066 31034
rect 43078 30982 43130 31034
rect 43142 30982 43194 31034
rect 43206 30982 43258 31034
rect 20812 30880 20864 30932
rect 22652 30880 22704 30932
rect 43536 30880 43588 30932
rect 39948 30744 40000 30796
rect 41420 30787 41472 30796
rect 41420 30753 41429 30787
rect 41429 30753 41463 30787
rect 41463 30753 41472 30787
rect 41420 30744 41472 30753
rect 22468 30719 22520 30728
rect 22468 30685 22477 30719
rect 22477 30685 22511 30719
rect 22511 30685 22520 30719
rect 22468 30676 22520 30685
rect 23388 30676 23440 30728
rect 40592 30719 40644 30728
rect 40592 30685 40601 30719
rect 40601 30685 40635 30719
rect 40635 30685 40644 30719
rect 40592 30676 40644 30685
rect 42800 30676 42852 30728
rect 43628 30676 43680 30728
rect 32864 30608 32916 30660
rect 33508 30651 33560 30660
rect 33508 30617 33517 30651
rect 33517 30617 33551 30651
rect 33551 30617 33560 30651
rect 33508 30608 33560 30617
rect 35440 30651 35492 30660
rect 35440 30617 35449 30651
rect 35449 30617 35483 30651
rect 35483 30617 35492 30651
rect 35440 30608 35492 30617
rect 37464 30608 37516 30660
rect 41696 30651 41748 30660
rect 41696 30617 41705 30651
rect 41705 30617 41739 30651
rect 41739 30617 41748 30651
rect 41696 30608 41748 30617
rect 38292 30540 38344 30592
rect 48596 30540 48648 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 27950 30438 28002 30490
rect 28014 30438 28066 30490
rect 28078 30438 28130 30490
rect 28142 30438 28194 30490
rect 28206 30438 28258 30490
rect 37950 30438 38002 30490
rect 38014 30438 38066 30490
rect 38078 30438 38130 30490
rect 38142 30438 38194 30490
rect 38206 30438 38258 30490
rect 47950 30438 48002 30490
rect 48014 30438 48066 30490
rect 48078 30438 48130 30490
rect 48142 30438 48194 30490
rect 48206 30438 48258 30490
rect 39120 30336 39172 30388
rect 35900 30268 35952 30320
rect 35992 30200 36044 30252
rect 37464 30200 37516 30252
rect 38476 30268 38528 30320
rect 43260 30336 43312 30388
rect 43536 30336 43588 30388
rect 40132 30268 40184 30320
rect 43628 30268 43680 30320
rect 35624 30175 35676 30184
rect 35624 30141 35633 30175
rect 35633 30141 35667 30175
rect 35667 30141 35676 30175
rect 35624 30132 35676 30141
rect 39672 30132 39724 30184
rect 39488 30064 39540 30116
rect 41420 30200 41472 30252
rect 42616 30243 42668 30252
rect 42616 30209 42625 30243
rect 42625 30209 42659 30243
rect 42659 30209 42668 30243
rect 42616 30200 42668 30209
rect 49332 30243 49384 30252
rect 49332 30209 49341 30243
rect 49341 30209 49375 30243
rect 49375 30209 49384 30243
rect 49332 30200 49384 30209
rect 34704 29996 34756 30048
rect 35164 29996 35216 30048
rect 35808 29996 35860 30048
rect 39028 29996 39080 30048
rect 39764 29996 39816 30048
rect 40592 29996 40644 30048
rect 42984 30132 43036 30184
rect 43536 30132 43588 30184
rect 41512 29996 41564 30048
rect 41696 29996 41748 30048
rect 48688 29996 48740 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 32950 29894 33002 29946
rect 33014 29894 33066 29946
rect 33078 29894 33130 29946
rect 33142 29894 33194 29946
rect 33206 29894 33258 29946
rect 42950 29894 43002 29946
rect 43014 29894 43066 29946
rect 43078 29894 43130 29946
rect 43142 29894 43194 29946
rect 43206 29894 43258 29946
rect 35624 29792 35676 29844
rect 41512 29792 41564 29844
rect 48964 29792 49016 29844
rect 34520 29724 34572 29776
rect 35072 29724 35124 29776
rect 41604 29724 41656 29776
rect 22836 29588 22888 29640
rect 33508 29656 33560 29708
rect 35532 29699 35584 29708
rect 35532 29665 35541 29699
rect 35541 29665 35575 29699
rect 35575 29665 35584 29699
rect 35532 29656 35584 29665
rect 35900 29656 35952 29708
rect 41512 29656 41564 29708
rect 32680 29588 32732 29640
rect 34612 29588 34664 29640
rect 48872 29724 48924 29776
rect 42616 29656 42668 29708
rect 33324 29520 33376 29572
rect 48412 29588 48464 29640
rect 49332 29631 49384 29640
rect 49332 29597 49341 29631
rect 49341 29597 49375 29631
rect 49375 29597 49384 29631
rect 49332 29588 49384 29597
rect 41972 29520 42024 29572
rect 31668 29452 31720 29504
rect 33600 29452 33652 29504
rect 41512 29452 41564 29504
rect 50160 29520 50212 29572
rect 48412 29452 48464 29504
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 27950 29350 28002 29402
rect 28014 29350 28066 29402
rect 28078 29350 28130 29402
rect 28142 29350 28194 29402
rect 28206 29350 28258 29402
rect 37950 29350 38002 29402
rect 38014 29350 38066 29402
rect 38078 29350 38130 29402
rect 38142 29350 38194 29402
rect 38206 29350 38258 29402
rect 47950 29350 48002 29402
rect 48014 29350 48066 29402
rect 48078 29350 48130 29402
rect 48142 29350 48194 29402
rect 48206 29350 48258 29402
rect 31392 29248 31444 29300
rect 34520 29248 34572 29300
rect 35256 29248 35308 29300
rect 34796 29180 34848 29232
rect 34888 29180 34940 29232
rect 35808 29180 35860 29232
rect 39120 29180 39172 29232
rect 34520 29112 34572 29164
rect 30288 29044 30340 29096
rect 31576 28976 31628 29028
rect 35164 29112 35216 29164
rect 37464 29155 37516 29164
rect 37464 29121 37473 29155
rect 37473 29121 37507 29155
rect 37507 29121 37516 29155
rect 37464 29112 37516 29121
rect 40040 29180 40092 29232
rect 41420 29180 41472 29232
rect 34336 28908 34388 28960
rect 39948 29087 40000 29096
rect 35808 28976 35860 29028
rect 35716 28908 35768 28960
rect 39948 29053 39957 29087
rect 39957 29053 39991 29087
rect 39991 29053 40000 29087
rect 39948 29044 40000 29053
rect 43536 29248 43588 29300
rect 43628 29180 43680 29232
rect 42616 29155 42668 29164
rect 42616 29121 42625 29155
rect 42625 29121 42659 29155
rect 42659 29121 42668 29155
rect 42616 29112 42668 29121
rect 48504 29044 48556 29096
rect 38476 28908 38528 28960
rect 39948 28908 40000 28960
rect 42432 28908 42484 28960
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 32950 28806 33002 28858
rect 33014 28806 33066 28858
rect 33078 28806 33130 28858
rect 33142 28806 33194 28858
rect 33206 28806 33258 28858
rect 42950 28806 43002 28858
rect 43014 28806 43066 28858
rect 43078 28806 43130 28858
rect 43142 28806 43194 28858
rect 43206 28806 43258 28858
rect 30656 28568 30708 28620
rect 35532 28568 35584 28620
rect 42064 28704 42116 28756
rect 30472 28432 30524 28484
rect 31944 28432 31996 28484
rect 32864 28432 32916 28484
rect 33416 28432 33468 28484
rect 38476 28568 38528 28620
rect 36176 28500 36228 28552
rect 39028 28500 39080 28552
rect 39396 28543 39448 28552
rect 39396 28509 39405 28543
rect 39405 28509 39439 28543
rect 39439 28509 39448 28543
rect 39396 28500 39448 28509
rect 40040 28543 40092 28552
rect 40040 28509 40049 28543
rect 40049 28509 40083 28543
rect 40083 28509 40092 28543
rect 40040 28500 40092 28509
rect 41420 28500 41472 28552
rect 43628 28704 43680 28756
rect 42616 28568 42668 28620
rect 43628 28500 43680 28552
rect 49332 28543 49384 28552
rect 49332 28509 49341 28543
rect 49341 28509 49375 28543
rect 49375 28509 49384 28543
rect 49332 28500 49384 28509
rect 32036 28407 32088 28416
rect 32036 28373 32045 28407
rect 32045 28373 32079 28407
rect 32079 28373 32088 28407
rect 32036 28364 32088 28373
rect 34888 28407 34940 28416
rect 34888 28373 34897 28407
rect 34897 28373 34931 28407
rect 34931 28373 34940 28407
rect 34888 28364 34940 28373
rect 35348 28407 35400 28416
rect 35348 28373 35357 28407
rect 35357 28373 35391 28407
rect 35391 28373 35400 28407
rect 35348 28364 35400 28373
rect 38844 28432 38896 28484
rect 39948 28432 40000 28484
rect 42524 28475 42576 28484
rect 39488 28364 39540 28416
rect 42524 28441 42533 28475
rect 42533 28441 42567 28475
rect 42567 28441 42576 28475
rect 42524 28432 42576 28441
rect 42432 28364 42484 28416
rect 46940 28364 46992 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 27950 28262 28002 28314
rect 28014 28262 28066 28314
rect 28078 28262 28130 28314
rect 28142 28262 28194 28314
rect 28206 28262 28258 28314
rect 37950 28262 38002 28314
rect 38014 28262 38066 28314
rect 38078 28262 38130 28314
rect 38142 28262 38194 28314
rect 38206 28262 38258 28314
rect 47950 28262 48002 28314
rect 48014 28262 48066 28314
rect 48078 28262 48130 28314
rect 48142 28262 48194 28314
rect 48206 28262 48258 28314
rect 22560 28160 22612 28212
rect 25596 28092 25648 28144
rect 25504 28024 25556 28076
rect 28448 28024 28500 28076
rect 30656 28160 30708 28212
rect 31484 28203 31536 28212
rect 31484 28169 31493 28203
rect 31493 28169 31527 28203
rect 31527 28169 31536 28203
rect 31484 28160 31536 28169
rect 32864 28160 32916 28212
rect 28816 28135 28868 28144
rect 28816 28101 28825 28135
rect 28825 28101 28859 28135
rect 28859 28101 28868 28135
rect 28816 28092 28868 28101
rect 30104 28092 30156 28144
rect 31944 28092 31996 28144
rect 33508 28092 33560 28144
rect 39396 28160 39448 28212
rect 40224 28203 40276 28212
rect 40224 28169 40233 28203
rect 40233 28169 40267 28203
rect 40267 28169 40276 28203
rect 40224 28160 40276 28169
rect 43904 28203 43956 28212
rect 35440 28135 35492 28144
rect 35440 28101 35471 28135
rect 35471 28101 35492 28135
rect 35440 28092 35492 28101
rect 24216 27999 24268 28008
rect 24216 27965 24225 27999
rect 24225 27965 24259 27999
rect 24259 27965 24268 27999
rect 24216 27956 24268 27965
rect 27528 27956 27580 28008
rect 31668 27956 31720 28008
rect 28908 27820 28960 27872
rect 30288 27863 30340 27872
rect 30288 27829 30297 27863
rect 30297 27829 30331 27863
rect 30331 27829 30340 27863
rect 30288 27820 30340 27829
rect 34612 28024 34664 28076
rect 39028 28092 39080 28144
rect 38384 28024 38436 28076
rect 40408 28024 40460 28076
rect 41512 28024 41564 28076
rect 43904 28169 43913 28203
rect 43913 28169 43947 28203
rect 43947 28169 43956 28203
rect 43904 28160 43956 28169
rect 46204 28160 46256 28212
rect 44180 28092 44232 28144
rect 33508 27999 33560 28008
rect 33508 27965 33517 27999
rect 33517 27965 33551 27999
rect 33551 27965 33560 27999
rect 33508 27956 33560 27965
rect 36176 27999 36228 28008
rect 36176 27965 36185 27999
rect 36185 27965 36219 27999
rect 36219 27965 36228 27999
rect 36176 27956 36228 27965
rect 38568 27999 38620 28008
rect 38568 27965 38577 27999
rect 38577 27965 38611 27999
rect 38611 27965 38620 27999
rect 38568 27956 38620 27965
rect 40316 27999 40368 28008
rect 40316 27965 40325 27999
rect 40325 27965 40359 27999
rect 40359 27965 40368 27999
rect 40316 27956 40368 27965
rect 35348 27888 35400 27940
rect 35624 27888 35676 27940
rect 44364 28024 44416 28076
rect 49332 28067 49384 28076
rect 49332 28033 49341 28067
rect 49341 28033 49375 28067
rect 49375 28033 49384 28067
rect 49332 28024 49384 28033
rect 34704 27820 34756 27872
rect 34980 27863 35032 27872
rect 34980 27829 34989 27863
rect 34989 27829 35023 27863
rect 35023 27829 35032 27863
rect 34980 27820 35032 27829
rect 37648 27820 37700 27872
rect 38384 27820 38436 27872
rect 39856 27820 39908 27872
rect 41788 27820 41840 27872
rect 44088 27999 44140 28008
rect 44088 27965 44097 27999
rect 44097 27965 44131 27999
rect 44131 27965 44140 27999
rect 44088 27956 44140 27965
rect 42064 27888 42116 27940
rect 49608 27888 49660 27940
rect 42616 27820 42668 27872
rect 48872 27820 48924 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 32950 27718 33002 27770
rect 33014 27718 33066 27770
rect 33078 27718 33130 27770
rect 33142 27718 33194 27770
rect 33206 27718 33258 27770
rect 42950 27718 43002 27770
rect 43014 27718 43066 27770
rect 43078 27718 43130 27770
rect 43142 27718 43194 27770
rect 43206 27718 43258 27770
rect 26148 27616 26200 27668
rect 32036 27616 32088 27668
rect 28448 27480 28500 27532
rect 30656 27480 30708 27532
rect 32680 27616 32732 27668
rect 34612 27616 34664 27668
rect 40408 27659 40460 27668
rect 40408 27625 40417 27659
rect 40417 27625 40451 27659
rect 40451 27625 40460 27659
rect 40408 27616 40460 27625
rect 32220 27548 32272 27600
rect 32128 27412 32180 27464
rect 24308 27344 24360 27396
rect 24768 27344 24820 27396
rect 24216 27276 24268 27328
rect 30840 27276 30892 27328
rect 34980 27480 35032 27532
rect 35716 27480 35768 27532
rect 39764 27480 39816 27532
rect 43904 27523 43956 27532
rect 43904 27489 43913 27523
rect 43913 27489 43947 27523
rect 43947 27489 43956 27523
rect 43904 27480 43956 27489
rect 35900 27455 35952 27464
rect 35900 27421 35909 27455
rect 35909 27421 35943 27455
rect 35943 27421 35952 27455
rect 35900 27412 35952 27421
rect 41696 27412 41748 27464
rect 41972 27455 42024 27464
rect 41972 27421 41981 27455
rect 41981 27421 42015 27455
rect 42015 27421 42024 27455
rect 41972 27412 42024 27421
rect 43720 27455 43772 27464
rect 43720 27421 43729 27455
rect 43729 27421 43763 27455
rect 43763 27421 43772 27455
rect 43720 27412 43772 27421
rect 46848 27412 46900 27464
rect 33600 27344 33652 27396
rect 40960 27344 41012 27396
rect 42708 27387 42760 27396
rect 42708 27353 42717 27387
rect 42717 27353 42751 27387
rect 42751 27353 42760 27387
rect 42708 27344 42760 27353
rect 33232 27276 33284 27328
rect 34888 27276 34940 27328
rect 35532 27319 35584 27328
rect 35532 27285 35541 27319
rect 35541 27285 35575 27319
rect 35575 27285 35584 27319
rect 35532 27276 35584 27285
rect 35992 27319 36044 27328
rect 35992 27285 36001 27319
rect 36001 27285 36035 27319
rect 36035 27285 36044 27319
rect 35992 27276 36044 27285
rect 40500 27276 40552 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 27950 27174 28002 27226
rect 28014 27174 28066 27226
rect 28078 27174 28130 27226
rect 28142 27174 28194 27226
rect 28206 27174 28258 27226
rect 37950 27174 38002 27226
rect 38014 27174 38066 27226
rect 38078 27174 38130 27226
rect 38142 27174 38194 27226
rect 38206 27174 38258 27226
rect 47950 27174 48002 27226
rect 48014 27174 48066 27226
rect 48078 27174 48130 27226
rect 48142 27174 48194 27226
rect 48206 27174 48258 27226
rect 30288 27072 30340 27124
rect 31392 27115 31444 27124
rect 31392 27081 31401 27115
rect 31401 27081 31435 27115
rect 31435 27081 31444 27115
rect 31392 27072 31444 27081
rect 31576 27072 31628 27124
rect 33324 27072 33376 27124
rect 33600 27072 33652 27124
rect 35256 27115 35308 27124
rect 35256 27081 35265 27115
rect 35265 27081 35299 27115
rect 35299 27081 35308 27115
rect 35256 27072 35308 27081
rect 39488 27115 39540 27124
rect 39488 27081 39497 27115
rect 39497 27081 39531 27115
rect 39531 27081 39540 27115
rect 39488 27072 39540 27081
rect 41696 27115 41748 27124
rect 41696 27081 41705 27115
rect 41705 27081 41739 27115
rect 41739 27081 41748 27115
rect 41696 27072 41748 27081
rect 41880 27072 41932 27124
rect 43812 27072 43864 27124
rect 47400 27072 47452 27124
rect 30104 27004 30156 27056
rect 39028 27004 39080 27056
rect 28448 26979 28500 26988
rect 28448 26945 28457 26979
rect 28457 26945 28491 26979
rect 28491 26945 28500 26979
rect 28448 26936 28500 26945
rect 34520 26936 34572 26988
rect 34704 26936 34756 26988
rect 49332 26979 49384 26988
rect 49332 26945 49341 26979
rect 49341 26945 49375 26979
rect 49375 26945 49384 26979
rect 49332 26936 49384 26945
rect 27712 26800 27764 26852
rect 24768 26732 24820 26784
rect 28172 26732 28224 26784
rect 32772 26868 32824 26920
rect 35164 26868 35216 26920
rect 35440 26911 35492 26920
rect 35440 26877 35449 26911
rect 35449 26877 35483 26911
rect 35483 26877 35492 26911
rect 35440 26868 35492 26877
rect 36176 26868 36228 26920
rect 39948 26868 40000 26920
rect 41604 26868 41656 26920
rect 45100 26868 45152 26920
rect 30104 26800 30156 26852
rect 30656 26732 30708 26784
rect 32680 26800 32732 26852
rect 41144 26732 41196 26784
rect 43628 26732 43680 26784
rect 47032 26732 47084 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 32950 26630 33002 26682
rect 33014 26630 33066 26682
rect 33078 26630 33130 26682
rect 33142 26630 33194 26682
rect 33206 26630 33258 26682
rect 42950 26630 43002 26682
rect 43014 26630 43066 26682
rect 43078 26630 43130 26682
rect 43142 26630 43194 26682
rect 43206 26630 43258 26682
rect 27344 26528 27396 26580
rect 30472 26528 30524 26580
rect 31484 26528 31536 26580
rect 27436 26435 27488 26444
rect 27436 26401 27445 26435
rect 27445 26401 27479 26435
rect 27479 26401 27488 26435
rect 27436 26392 27488 26401
rect 28448 26392 28500 26444
rect 30564 26435 30616 26444
rect 30564 26401 30573 26435
rect 30573 26401 30607 26435
rect 30607 26401 30616 26435
rect 30564 26392 30616 26401
rect 36268 26460 36320 26512
rect 44088 26460 44140 26512
rect 30840 26435 30892 26444
rect 30840 26401 30849 26435
rect 30849 26401 30883 26435
rect 30883 26401 30892 26435
rect 30840 26392 30892 26401
rect 33508 26392 33560 26444
rect 34152 26392 34204 26444
rect 35072 26392 35124 26444
rect 35440 26435 35492 26444
rect 35440 26401 35449 26435
rect 35449 26401 35483 26435
rect 35483 26401 35492 26435
rect 35440 26392 35492 26401
rect 38292 26392 38344 26444
rect 38844 26435 38896 26444
rect 38844 26401 38853 26435
rect 38853 26401 38887 26435
rect 38887 26401 38896 26435
rect 38844 26392 38896 26401
rect 42708 26392 42760 26444
rect 42892 26392 42944 26444
rect 43352 26392 43404 26444
rect 35256 26367 35308 26376
rect 35256 26333 35265 26367
rect 35265 26333 35299 26367
rect 35299 26333 35308 26367
rect 35256 26324 35308 26333
rect 40132 26367 40184 26376
rect 40132 26333 40141 26367
rect 40141 26333 40175 26367
rect 40175 26333 40184 26367
rect 40132 26324 40184 26333
rect 42524 26367 42576 26376
rect 42524 26333 42533 26367
rect 42533 26333 42567 26367
rect 42567 26333 42576 26367
rect 42524 26324 42576 26333
rect 48504 26367 48556 26376
rect 48504 26333 48513 26367
rect 48513 26333 48547 26367
rect 48547 26333 48556 26367
rect 48504 26324 48556 26333
rect 48596 26324 48648 26376
rect 25228 26256 25280 26308
rect 27712 26299 27764 26308
rect 27712 26265 27721 26299
rect 27721 26265 27755 26299
rect 27755 26265 27764 26299
rect 27712 26256 27764 26265
rect 28172 26256 28224 26308
rect 32128 26256 32180 26308
rect 39764 26256 39816 26308
rect 39028 26188 39080 26240
rect 43352 26256 43404 26308
rect 45468 26256 45520 26308
rect 41420 26188 41472 26240
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 27950 26086 28002 26138
rect 28014 26086 28066 26138
rect 28078 26086 28130 26138
rect 28142 26086 28194 26138
rect 28206 26086 28258 26138
rect 37950 26086 38002 26138
rect 38014 26086 38066 26138
rect 38078 26086 38130 26138
rect 38142 26086 38194 26138
rect 38206 26086 38258 26138
rect 47950 26086 48002 26138
rect 48014 26086 48066 26138
rect 48078 26086 48130 26138
rect 48142 26086 48194 26138
rect 48206 26086 48258 26138
rect 32036 25984 32088 26036
rect 27436 25916 27488 25968
rect 31852 25916 31904 25968
rect 33048 25916 33100 25968
rect 34428 25916 34480 25968
rect 28540 25848 28592 25900
rect 35532 25984 35584 26036
rect 35808 26027 35860 26036
rect 35808 25993 35817 26027
rect 35817 25993 35851 26027
rect 35851 25993 35860 26027
rect 35808 25984 35860 25993
rect 40132 25984 40184 26036
rect 42524 25984 42576 26036
rect 41420 25916 41472 25968
rect 41880 25916 41932 25968
rect 42708 25984 42760 26036
rect 26424 25780 26476 25832
rect 27528 25780 27580 25832
rect 28724 25712 28776 25764
rect 28816 25644 28868 25696
rect 29000 25644 29052 25696
rect 34980 25780 35032 25832
rect 44364 25848 44416 25900
rect 45100 25959 45152 25968
rect 45100 25925 45109 25959
rect 45109 25925 45143 25959
rect 45143 25925 45152 25959
rect 45100 25916 45152 25925
rect 46112 25916 46164 25968
rect 41696 25780 41748 25832
rect 33600 25644 33652 25696
rect 36176 25712 36228 25764
rect 39948 25712 40000 25764
rect 35348 25687 35400 25696
rect 35348 25653 35357 25687
rect 35357 25653 35391 25687
rect 35391 25653 35400 25687
rect 35348 25644 35400 25653
rect 37740 25644 37792 25696
rect 40408 25644 40460 25696
rect 42432 25780 42484 25832
rect 43536 25780 43588 25832
rect 43444 25644 43496 25696
rect 43996 25644 44048 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 32950 25542 33002 25594
rect 33014 25542 33066 25594
rect 33078 25542 33130 25594
rect 33142 25542 33194 25594
rect 33206 25542 33258 25594
rect 42950 25542 43002 25594
rect 43014 25542 43066 25594
rect 43078 25542 43130 25594
rect 43142 25542 43194 25594
rect 43206 25542 43258 25594
rect 24860 25440 24912 25492
rect 28724 25440 28776 25492
rect 32496 25440 32548 25492
rect 30472 25372 30524 25424
rect 30656 25347 30708 25356
rect 30656 25313 30665 25347
rect 30665 25313 30699 25347
rect 30699 25313 30708 25347
rect 30656 25304 30708 25313
rect 38568 25372 38620 25424
rect 32772 25304 32824 25356
rect 32956 25304 33008 25356
rect 33324 25304 33376 25356
rect 34152 25347 34204 25356
rect 34152 25313 34161 25347
rect 34161 25313 34195 25347
rect 34195 25313 34204 25347
rect 34152 25304 34204 25313
rect 34520 25304 34572 25356
rect 38476 25304 38528 25356
rect 40684 25304 40736 25356
rect 41788 25415 41840 25424
rect 41788 25381 41797 25415
rect 41797 25381 41831 25415
rect 41831 25381 41840 25415
rect 41788 25372 41840 25381
rect 43904 25372 43956 25424
rect 44088 25304 44140 25356
rect 45652 25347 45704 25356
rect 45652 25313 45661 25347
rect 45661 25313 45695 25347
rect 45695 25313 45704 25347
rect 45652 25304 45704 25313
rect 45928 25304 45980 25356
rect 37740 25279 37792 25288
rect 37740 25245 37749 25279
rect 37749 25245 37783 25279
rect 37783 25245 37792 25279
rect 37740 25236 37792 25245
rect 40040 25279 40092 25288
rect 40040 25245 40049 25279
rect 40049 25245 40083 25279
rect 40083 25245 40092 25279
rect 40040 25236 40092 25245
rect 44364 25236 44416 25288
rect 45468 25236 45520 25288
rect 49148 25279 49200 25288
rect 49148 25245 49157 25279
rect 49157 25245 49191 25279
rect 49191 25245 49200 25279
rect 49148 25236 49200 25245
rect 30380 25168 30432 25220
rect 30564 25143 30616 25152
rect 30564 25109 30573 25143
rect 30573 25109 30607 25143
rect 30607 25109 30616 25143
rect 30564 25100 30616 25109
rect 31300 25168 31352 25220
rect 35900 25168 35952 25220
rect 40592 25168 40644 25220
rect 41880 25168 41932 25220
rect 32864 25143 32916 25152
rect 32864 25109 32873 25143
rect 32873 25109 32907 25143
rect 32907 25109 32916 25143
rect 32864 25100 32916 25109
rect 35072 25100 35124 25152
rect 36636 25100 36688 25152
rect 36728 25143 36780 25152
rect 36728 25109 36737 25143
rect 36737 25109 36771 25143
rect 36771 25109 36780 25143
rect 36728 25100 36780 25109
rect 37372 25143 37424 25152
rect 37372 25109 37381 25143
rect 37381 25109 37415 25143
rect 37415 25109 37424 25143
rect 37372 25100 37424 25109
rect 43996 25100 44048 25152
rect 45560 25143 45612 25152
rect 45560 25109 45569 25143
rect 45569 25109 45603 25143
rect 45603 25109 45612 25143
rect 45560 25100 45612 25109
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 27950 24998 28002 25050
rect 28014 24998 28066 25050
rect 28078 24998 28130 25050
rect 28142 24998 28194 25050
rect 28206 24998 28258 25050
rect 37950 24998 38002 25050
rect 38014 24998 38066 25050
rect 38078 24998 38130 25050
rect 38142 24998 38194 25050
rect 38206 24998 38258 25050
rect 47950 24998 48002 25050
rect 48014 24998 48066 25050
rect 48078 24998 48130 25050
rect 48142 24998 48194 25050
rect 48206 24998 48258 25050
rect 32680 24896 32732 24948
rect 33416 24896 33468 24948
rect 34612 24896 34664 24948
rect 35900 24896 35952 24948
rect 36544 24939 36596 24948
rect 36544 24905 36553 24939
rect 36553 24905 36587 24939
rect 36587 24905 36596 24939
rect 36544 24896 36596 24905
rect 36728 24896 36780 24948
rect 43996 24896 44048 24948
rect 31484 24803 31536 24812
rect 31484 24769 31493 24803
rect 31493 24769 31527 24803
rect 31527 24769 31536 24803
rect 31484 24760 31536 24769
rect 34428 24828 34480 24880
rect 41880 24828 41932 24880
rect 44364 24828 44416 24880
rect 46020 24828 46072 24880
rect 36636 24803 36688 24812
rect 36636 24769 36645 24803
rect 36645 24769 36679 24803
rect 36679 24769 36688 24803
rect 36636 24760 36688 24769
rect 37740 24803 37792 24812
rect 37740 24769 37749 24803
rect 37749 24769 37783 24803
rect 37783 24769 37792 24803
rect 37740 24760 37792 24769
rect 38568 24803 38620 24812
rect 38568 24769 38577 24803
rect 38577 24769 38611 24803
rect 38611 24769 38620 24803
rect 38568 24760 38620 24769
rect 41696 24760 41748 24812
rect 42984 24803 43036 24812
rect 42984 24769 42993 24803
rect 42993 24769 43027 24803
rect 43027 24769 43036 24803
rect 42984 24760 43036 24769
rect 29460 24692 29512 24744
rect 32588 24692 32640 24744
rect 32956 24735 33008 24744
rect 32956 24701 32965 24735
rect 32965 24701 32999 24735
rect 32999 24701 33008 24735
rect 32956 24692 33008 24701
rect 33600 24735 33652 24744
rect 33600 24701 33609 24735
rect 33609 24701 33643 24735
rect 33643 24701 33652 24735
rect 33600 24692 33652 24701
rect 33876 24735 33928 24744
rect 33876 24701 33885 24735
rect 33885 24701 33919 24735
rect 33919 24701 33928 24735
rect 33876 24692 33928 24701
rect 33508 24624 33560 24676
rect 34888 24624 34940 24676
rect 42064 24624 42116 24676
rect 27068 24556 27120 24608
rect 29000 24556 29052 24608
rect 31024 24599 31076 24608
rect 31024 24565 31033 24599
rect 31033 24565 31067 24599
rect 31067 24565 31076 24599
rect 31024 24556 31076 24565
rect 31116 24556 31168 24608
rect 32404 24556 32456 24608
rect 35440 24556 35492 24608
rect 36636 24556 36688 24608
rect 37832 24599 37884 24608
rect 37832 24565 37841 24599
rect 37841 24565 37875 24599
rect 37875 24565 37884 24599
rect 37832 24556 37884 24565
rect 38384 24599 38436 24608
rect 38384 24565 38393 24599
rect 38393 24565 38427 24599
rect 38427 24565 38436 24599
rect 38384 24556 38436 24565
rect 39212 24556 39264 24608
rect 44088 24760 44140 24812
rect 45836 24760 45888 24812
rect 43444 24692 43496 24744
rect 45100 24692 45152 24744
rect 49148 24735 49200 24744
rect 49148 24701 49157 24735
rect 49157 24701 49191 24735
rect 49191 24701 49200 24735
rect 49148 24692 49200 24701
rect 48412 24556 48464 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 22836 24352 22888 24404
rect 27160 24284 27212 24336
rect 27528 24216 27580 24268
rect 28816 24284 28868 24336
rect 27804 24080 27856 24132
rect 28908 24259 28960 24268
rect 28908 24225 28917 24259
rect 28917 24225 28951 24259
rect 28951 24225 28960 24259
rect 28908 24216 28960 24225
rect 33508 24284 33560 24336
rect 31208 24216 31260 24268
rect 33600 24216 33652 24268
rect 35624 24284 35676 24336
rect 29736 24191 29788 24200
rect 29736 24157 29745 24191
rect 29745 24157 29779 24191
rect 29779 24157 29788 24191
rect 29736 24148 29788 24157
rect 34428 24148 34480 24200
rect 35256 24191 35308 24200
rect 35256 24157 35265 24191
rect 35265 24157 35299 24191
rect 35299 24157 35308 24191
rect 35256 24148 35308 24157
rect 31392 24080 31444 24132
rect 32128 24080 32180 24132
rect 32312 24080 32364 24132
rect 43168 24352 43220 24404
rect 49516 24352 49568 24404
rect 38384 24284 38436 24336
rect 46572 24284 46624 24336
rect 42800 24216 42852 24268
rect 45744 24259 45796 24268
rect 45744 24225 45753 24259
rect 45753 24225 45787 24259
rect 45787 24225 45796 24259
rect 45744 24216 45796 24225
rect 38660 24148 38712 24200
rect 40316 24148 40368 24200
rect 43260 24148 43312 24200
rect 43536 24148 43588 24200
rect 43812 24148 43864 24200
rect 48688 24216 48740 24268
rect 46572 24191 46624 24200
rect 46572 24157 46581 24191
rect 46581 24157 46615 24191
rect 46615 24157 46624 24191
rect 46572 24148 46624 24157
rect 28632 24012 28684 24064
rect 29368 24012 29420 24064
rect 32588 24012 32640 24064
rect 32956 24012 33008 24064
rect 37740 24080 37792 24132
rect 43168 24080 43220 24132
rect 43720 24080 43772 24132
rect 48320 24080 48372 24132
rect 33784 24012 33836 24064
rect 43352 24012 43404 24064
rect 43536 24055 43588 24064
rect 43536 24021 43545 24055
rect 43545 24021 43579 24055
rect 43579 24021 43588 24055
rect 43536 24012 43588 24021
rect 45192 24055 45244 24064
rect 45192 24021 45201 24055
rect 45201 24021 45235 24055
rect 45235 24021 45244 24055
rect 45192 24012 45244 24021
rect 46388 24055 46440 24064
rect 46388 24021 46397 24055
rect 46397 24021 46431 24055
rect 46431 24021 46440 24055
rect 46388 24012 46440 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 25596 23851 25648 23860
rect 25596 23817 25605 23851
rect 25605 23817 25639 23851
rect 25639 23817 25648 23851
rect 25596 23808 25648 23817
rect 27068 23808 27120 23860
rect 28540 23672 28592 23724
rect 29736 23808 29788 23860
rect 26056 23647 26108 23656
rect 26056 23613 26065 23647
rect 26065 23613 26099 23647
rect 26099 23613 26108 23647
rect 26056 23604 26108 23613
rect 26148 23647 26200 23656
rect 26148 23613 26157 23647
rect 26157 23613 26191 23647
rect 26191 23613 26200 23647
rect 26148 23604 26200 23613
rect 29368 23604 29420 23656
rect 28540 23536 28592 23588
rect 29000 23536 29052 23588
rect 28908 23511 28960 23520
rect 28908 23477 28917 23511
rect 28917 23477 28951 23511
rect 28951 23477 28960 23511
rect 28908 23468 28960 23477
rect 29460 23536 29512 23588
rect 31392 23740 31444 23792
rect 32404 23808 32456 23860
rect 32864 23808 32916 23860
rect 32036 23740 32088 23792
rect 34428 23740 34480 23792
rect 34704 23740 34756 23792
rect 34980 23740 35032 23792
rect 34796 23672 34848 23724
rect 35256 23740 35308 23792
rect 37740 23672 37792 23724
rect 38660 23783 38712 23792
rect 38660 23749 38669 23783
rect 38669 23749 38703 23783
rect 38703 23749 38712 23783
rect 38660 23740 38712 23749
rect 39856 23740 39908 23792
rect 40316 23783 40368 23792
rect 40316 23749 40325 23783
rect 40325 23749 40359 23783
rect 40359 23749 40368 23783
rect 40316 23740 40368 23749
rect 40500 23740 40552 23792
rect 41972 23740 42024 23792
rect 44088 23783 44140 23792
rect 44088 23749 44097 23783
rect 44097 23749 44131 23783
rect 44131 23749 44140 23783
rect 44088 23740 44140 23749
rect 39028 23672 39080 23724
rect 44640 23715 44692 23724
rect 44640 23681 44649 23715
rect 44649 23681 44683 23715
rect 44683 23681 44692 23715
rect 44640 23672 44692 23681
rect 46020 23672 46072 23724
rect 46388 23672 46440 23724
rect 31208 23647 31260 23656
rect 31208 23613 31217 23647
rect 31217 23613 31251 23647
rect 31251 23613 31260 23647
rect 31208 23604 31260 23613
rect 33876 23604 33928 23656
rect 35440 23647 35492 23656
rect 35440 23613 35449 23647
rect 35449 23613 35483 23647
rect 35483 23613 35492 23647
rect 35440 23604 35492 23613
rect 34796 23536 34848 23588
rect 35624 23604 35676 23656
rect 30932 23468 30984 23520
rect 32680 23468 32732 23520
rect 32956 23468 33008 23520
rect 35256 23468 35308 23520
rect 35532 23468 35584 23520
rect 37004 23604 37056 23656
rect 37556 23604 37608 23656
rect 36912 23536 36964 23588
rect 39948 23604 40000 23656
rect 40684 23604 40736 23656
rect 45928 23604 45980 23656
rect 46664 23604 46716 23656
rect 49148 23647 49200 23656
rect 49148 23613 49157 23647
rect 49157 23613 49191 23647
rect 49191 23613 49200 23647
rect 49148 23604 49200 23613
rect 38844 23468 38896 23520
rect 40040 23536 40092 23588
rect 41328 23536 41380 23588
rect 43444 23468 43496 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 24032 23264 24084 23316
rect 24860 23171 24912 23180
rect 24860 23137 24869 23171
rect 24869 23137 24903 23171
rect 24903 23137 24912 23171
rect 24860 23128 24912 23137
rect 25412 23128 25464 23180
rect 26148 23264 26200 23316
rect 28908 23128 28960 23180
rect 24584 23103 24636 23112
rect 24584 23069 24593 23103
rect 24593 23069 24627 23103
rect 24627 23069 24636 23103
rect 24584 23060 24636 23069
rect 30104 23103 30156 23112
rect 30104 23069 30113 23103
rect 30113 23069 30147 23103
rect 30147 23069 30156 23103
rect 30104 23060 30156 23069
rect 31116 23060 31168 23112
rect 26608 22992 26660 23044
rect 26700 22992 26752 23044
rect 34980 23264 35032 23316
rect 40868 23264 40920 23316
rect 35440 23196 35492 23248
rect 39120 23196 39172 23248
rect 42800 23196 42852 23248
rect 33416 23171 33468 23180
rect 33416 23137 33425 23171
rect 33425 23137 33459 23171
rect 33459 23137 33468 23171
rect 33416 23128 33468 23137
rect 38384 23128 38436 23180
rect 37740 23060 37792 23112
rect 39304 23128 39356 23180
rect 40040 23128 40092 23180
rect 41512 23128 41564 23180
rect 46940 23196 46992 23248
rect 44364 23128 44416 23180
rect 27252 22924 27304 22976
rect 30104 22924 30156 22976
rect 32220 22924 32272 22976
rect 32496 22924 32548 22976
rect 32864 22967 32916 22976
rect 32864 22933 32873 22967
rect 32873 22933 32907 22967
rect 32907 22933 32916 22967
rect 32864 22924 32916 22933
rect 33508 22992 33560 23044
rect 40132 23060 40184 23112
rect 41880 23060 41932 23112
rect 42984 23060 43036 23112
rect 40776 23035 40828 23044
rect 40776 23001 40785 23035
rect 40785 23001 40819 23035
rect 40819 23001 40828 23035
rect 40776 22992 40828 23001
rect 34060 22924 34112 22976
rect 43720 22992 43772 23044
rect 44180 22992 44232 23044
rect 46756 22992 46808 23044
rect 49148 23035 49200 23044
rect 49148 23001 49157 23035
rect 49157 23001 49191 23035
rect 49191 23001 49200 23035
rect 49148 22992 49200 23001
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 27620 22720 27672 22772
rect 33416 22720 33468 22772
rect 35348 22720 35400 22772
rect 36544 22720 36596 22772
rect 36728 22652 36780 22704
rect 33416 22584 33468 22636
rect 40040 22720 40092 22772
rect 40132 22720 40184 22772
rect 41420 22720 41472 22772
rect 41696 22720 41748 22772
rect 42984 22763 43036 22772
rect 42984 22729 42993 22763
rect 42993 22729 43027 22763
rect 43027 22729 43036 22763
rect 42984 22720 43036 22729
rect 43628 22720 43680 22772
rect 40592 22652 40644 22704
rect 41512 22584 41564 22636
rect 33968 22559 34020 22568
rect 33968 22525 33977 22559
rect 33977 22525 34011 22559
rect 34011 22525 34020 22559
rect 33968 22516 34020 22525
rect 33508 22448 33560 22500
rect 37740 22448 37792 22500
rect 39304 22559 39356 22568
rect 39304 22525 39313 22559
rect 39313 22525 39347 22559
rect 39347 22525 39356 22559
rect 39304 22516 39356 22525
rect 39396 22516 39448 22568
rect 40776 22559 40828 22568
rect 40776 22525 40785 22559
rect 40785 22525 40819 22559
rect 40819 22525 40828 22559
rect 40776 22516 40828 22525
rect 43996 22695 44048 22704
rect 43996 22661 44005 22695
rect 44005 22661 44039 22695
rect 44039 22661 44048 22695
rect 43996 22652 44048 22661
rect 45836 22720 45888 22772
rect 46664 22763 46716 22772
rect 46664 22729 46673 22763
rect 46673 22729 46707 22763
rect 46707 22729 46716 22763
rect 46664 22720 46716 22729
rect 45928 22652 45980 22704
rect 44640 22584 44692 22636
rect 44916 22627 44968 22636
rect 44916 22593 44925 22627
rect 44925 22593 44959 22627
rect 44959 22593 44968 22627
rect 44916 22584 44968 22593
rect 38476 22380 38528 22432
rect 39672 22380 39724 22432
rect 43352 22516 43404 22568
rect 44548 22516 44600 22568
rect 40408 22380 40460 22432
rect 47032 22380 47084 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 30196 22219 30248 22228
rect 24584 22108 24636 22160
rect 30196 22185 30226 22219
rect 30226 22185 30248 22219
rect 30196 22176 30248 22185
rect 34520 22176 34572 22228
rect 39488 22176 39540 22228
rect 40408 22176 40460 22228
rect 42800 22176 42852 22228
rect 26792 22040 26844 22092
rect 29184 22108 29236 22160
rect 25412 21972 25464 22024
rect 33324 22108 33376 22160
rect 33508 22108 33560 22160
rect 35900 22108 35952 22160
rect 32864 22040 32916 22092
rect 35440 22040 35492 22092
rect 39304 22108 39356 22160
rect 42064 22108 42116 22160
rect 29736 21972 29788 22024
rect 27068 21904 27120 21956
rect 30932 21904 30984 21956
rect 26424 21836 26476 21888
rect 27528 21879 27580 21888
rect 27528 21845 27537 21879
rect 27537 21845 27571 21879
rect 27571 21845 27580 21879
rect 27528 21836 27580 21845
rect 27804 21836 27856 21888
rect 30840 21836 30892 21888
rect 34980 21904 35032 21956
rect 31668 21879 31720 21888
rect 31668 21845 31677 21879
rect 31677 21845 31711 21879
rect 31711 21845 31720 21879
rect 31668 21836 31720 21845
rect 37280 21904 37332 21956
rect 39212 22083 39264 22092
rect 39212 22049 39221 22083
rect 39221 22049 39255 22083
rect 39255 22049 39264 22083
rect 39212 22040 39264 22049
rect 39396 22083 39448 22092
rect 39396 22049 39405 22083
rect 39405 22049 39439 22083
rect 39439 22049 39448 22083
rect 39396 22040 39448 22049
rect 39120 22015 39172 22024
rect 39120 21981 39129 22015
rect 39129 21981 39163 22015
rect 39163 21981 39172 22015
rect 39120 21972 39172 21981
rect 44180 22040 44232 22092
rect 45560 22040 45612 22092
rect 41328 21972 41380 22024
rect 44916 21972 44968 22024
rect 46756 21972 46808 22024
rect 49148 22015 49200 22024
rect 49148 21981 49157 22015
rect 49157 21981 49191 22015
rect 49191 21981 49200 22015
rect 49148 21972 49200 21981
rect 41604 21904 41656 21956
rect 45928 21904 45980 21956
rect 37188 21836 37240 21888
rect 43904 21836 43956 21888
rect 44548 21836 44600 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 25504 21675 25556 21684
rect 25504 21641 25513 21675
rect 25513 21641 25547 21675
rect 25547 21641 25556 21675
rect 25504 21632 25556 21641
rect 26608 21632 26660 21684
rect 26884 21632 26936 21684
rect 26976 21564 27028 21616
rect 30380 21632 30432 21684
rect 30840 21632 30892 21684
rect 31024 21632 31076 21684
rect 32772 21632 32824 21684
rect 38384 21632 38436 21684
rect 39028 21675 39080 21684
rect 39028 21641 39037 21675
rect 39037 21641 39071 21675
rect 39071 21641 39080 21675
rect 39028 21632 39080 21641
rect 43720 21632 43772 21684
rect 43996 21632 44048 21684
rect 44916 21632 44968 21684
rect 45744 21675 45796 21684
rect 45744 21641 45753 21675
rect 45753 21641 45787 21675
rect 45787 21641 45796 21675
rect 45744 21632 45796 21641
rect 29000 21564 29052 21616
rect 30472 21564 30524 21616
rect 34428 21564 34480 21616
rect 35348 21564 35400 21616
rect 38844 21564 38896 21616
rect 43812 21564 43864 21616
rect 45928 21564 45980 21616
rect 27528 21539 27580 21548
rect 27528 21505 27537 21539
rect 27537 21505 27571 21539
rect 27571 21505 27580 21539
rect 27528 21496 27580 21505
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 26516 21428 26568 21480
rect 26700 21360 26752 21412
rect 27344 21360 27396 21412
rect 27804 21428 27856 21480
rect 28724 21471 28776 21480
rect 28724 21437 28733 21471
rect 28733 21437 28767 21471
rect 28767 21437 28776 21471
rect 28724 21428 28776 21437
rect 37832 21539 37884 21548
rect 37832 21505 37841 21539
rect 37841 21505 37875 21539
rect 37875 21505 37884 21539
rect 37832 21496 37884 21505
rect 40592 21496 40644 21548
rect 24952 21335 25004 21344
rect 24952 21301 24961 21335
rect 24961 21301 24995 21335
rect 24995 21301 25004 21335
rect 24952 21292 25004 21301
rect 25136 21292 25188 21344
rect 31208 21471 31260 21480
rect 31208 21437 31217 21471
rect 31217 21437 31251 21471
rect 31251 21437 31260 21471
rect 31208 21428 31260 21437
rect 31024 21360 31076 21412
rect 31668 21360 31720 21412
rect 34520 21428 34572 21480
rect 35072 21471 35124 21480
rect 35072 21437 35081 21471
rect 35081 21437 35115 21471
rect 35115 21437 35124 21471
rect 35072 21428 35124 21437
rect 35440 21428 35492 21480
rect 38752 21428 38804 21480
rect 39028 21428 39080 21480
rect 38844 21360 38896 21412
rect 41788 21360 41840 21412
rect 47032 21496 47084 21548
rect 43996 21471 44048 21480
rect 43996 21437 44005 21471
rect 44005 21437 44039 21471
rect 44039 21437 44048 21471
rect 43996 21428 44048 21437
rect 48872 21428 48924 21480
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 30196 21335 30248 21344
rect 30196 21301 30205 21335
rect 30205 21301 30239 21335
rect 30239 21301 30248 21335
rect 30196 21292 30248 21301
rect 36452 21292 36504 21344
rect 36544 21335 36596 21344
rect 36544 21301 36553 21335
rect 36553 21301 36587 21335
rect 36587 21301 36596 21335
rect 36544 21292 36596 21301
rect 39212 21292 39264 21344
rect 42800 21335 42852 21344
rect 42800 21301 42809 21335
rect 42809 21301 42843 21335
rect 42843 21301 42852 21335
rect 42800 21292 42852 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 27528 21088 27580 21140
rect 30288 21088 30340 21140
rect 32680 21088 32732 21140
rect 37004 21088 37056 21140
rect 37832 21088 37884 21140
rect 42064 21088 42116 21140
rect 30564 21020 30616 21072
rect 36452 21020 36504 21072
rect 25228 20995 25280 21004
rect 25228 20961 25237 20995
rect 25237 20961 25271 20995
rect 25271 20961 25280 20995
rect 25228 20952 25280 20961
rect 26424 20995 26476 21004
rect 26424 20961 26433 20995
rect 26433 20961 26467 20995
rect 26467 20961 26476 20995
rect 26424 20952 26476 20961
rect 31024 20995 31076 21004
rect 31024 20961 31033 20995
rect 31033 20961 31067 20995
rect 31067 20961 31076 20995
rect 31024 20952 31076 20961
rect 31760 20952 31812 21004
rect 33600 20952 33652 21004
rect 36544 20952 36596 21004
rect 24952 20927 25004 20936
rect 24952 20893 24961 20927
rect 24961 20893 24995 20927
rect 24995 20893 25004 20927
rect 24952 20884 25004 20893
rect 25412 20884 25464 20936
rect 29736 20884 29788 20936
rect 33784 20884 33836 20936
rect 43628 21020 43680 21072
rect 43444 20995 43496 21004
rect 43444 20961 43453 20995
rect 43453 20961 43487 20995
rect 43487 20961 43496 20995
rect 43444 20952 43496 20961
rect 40040 20884 40092 20936
rect 41604 20884 41656 20936
rect 26884 20816 26936 20868
rect 27712 20816 27764 20868
rect 30932 20816 30984 20868
rect 25044 20791 25096 20800
rect 25044 20757 25053 20791
rect 25053 20757 25087 20791
rect 25087 20757 25096 20791
rect 25044 20748 25096 20757
rect 29276 20748 29328 20800
rect 35348 20816 35400 20868
rect 37096 20816 37148 20868
rect 38752 20816 38804 20868
rect 40500 20859 40552 20868
rect 40500 20825 40509 20859
rect 40509 20825 40543 20859
rect 40543 20825 40552 20859
rect 40500 20816 40552 20825
rect 34428 20748 34480 20800
rect 44088 20816 44140 20868
rect 43904 20748 43956 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 28724 20544 28776 20596
rect 31760 20587 31812 20596
rect 31760 20553 31769 20587
rect 31769 20553 31803 20587
rect 31803 20553 31812 20587
rect 31760 20544 31812 20553
rect 27528 20476 27580 20528
rect 29644 20476 29696 20528
rect 30288 20519 30340 20528
rect 30288 20485 30297 20519
rect 30297 20485 30331 20519
rect 30331 20485 30340 20519
rect 30288 20476 30340 20485
rect 30932 20476 30984 20528
rect 25320 20408 25372 20460
rect 26884 20408 26936 20460
rect 34520 20476 34572 20528
rect 36636 20587 36688 20596
rect 36636 20553 36645 20587
rect 36645 20553 36679 20587
rect 36679 20553 36688 20587
rect 36636 20544 36688 20553
rect 45192 20544 45244 20596
rect 38660 20476 38712 20528
rect 41604 20476 41656 20528
rect 47032 20476 47084 20528
rect 35348 20408 35400 20460
rect 35992 20408 36044 20460
rect 39948 20408 40000 20460
rect 46940 20408 46992 20460
rect 23756 20383 23808 20392
rect 23756 20349 23765 20383
rect 23765 20349 23799 20383
rect 23799 20349 23808 20383
rect 23756 20340 23808 20349
rect 24032 20383 24084 20392
rect 24032 20349 24041 20383
rect 24041 20349 24075 20383
rect 24075 20349 24084 20383
rect 24032 20340 24084 20349
rect 25412 20340 25464 20392
rect 26608 20272 26660 20324
rect 29736 20340 29788 20392
rect 34704 20340 34756 20392
rect 36636 20340 36688 20392
rect 26240 20204 26292 20256
rect 35440 20204 35492 20256
rect 38752 20340 38804 20392
rect 44548 20383 44600 20392
rect 44548 20349 44557 20383
rect 44557 20349 44591 20383
rect 44591 20349 44600 20383
rect 44548 20340 44600 20349
rect 49148 20383 49200 20392
rect 49148 20349 49157 20383
rect 49157 20349 49191 20383
rect 49191 20349 49200 20383
rect 49148 20340 49200 20349
rect 40040 20204 40092 20256
rect 40132 20247 40184 20256
rect 40132 20213 40141 20247
rect 40141 20213 40175 20247
rect 40175 20213 40184 20247
rect 40132 20204 40184 20213
rect 42156 20204 42208 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 29184 20043 29236 20052
rect 29184 20009 29193 20043
rect 29193 20009 29227 20043
rect 29227 20009 29236 20043
rect 29184 20000 29236 20009
rect 34796 20000 34848 20052
rect 39948 20000 40000 20052
rect 40132 20000 40184 20052
rect 41788 20043 41840 20052
rect 41788 20009 41797 20043
rect 41797 20009 41831 20043
rect 41831 20009 41840 20043
rect 41788 20000 41840 20009
rect 44364 20000 44416 20052
rect 23756 19864 23808 19916
rect 25412 19864 25464 19916
rect 27804 19864 27856 19916
rect 28908 19864 28960 19916
rect 32588 19839 32640 19848
rect 32588 19805 32597 19839
rect 32597 19805 32631 19839
rect 32631 19805 32640 19839
rect 32588 19796 32640 19805
rect 35072 19839 35124 19848
rect 35072 19805 35081 19839
rect 35081 19805 35115 19839
rect 35115 19805 35124 19839
rect 35072 19796 35124 19805
rect 40040 19907 40092 19916
rect 40040 19873 40049 19907
rect 40049 19873 40083 19907
rect 40083 19873 40092 19907
rect 40040 19864 40092 19873
rect 41328 19864 41380 19916
rect 43996 19864 44048 19916
rect 38844 19839 38896 19848
rect 38844 19805 38853 19839
rect 38853 19805 38887 19839
rect 38887 19805 38896 19839
rect 38844 19796 38896 19805
rect 39672 19796 39724 19848
rect 41604 19796 41656 19848
rect 25320 19728 25372 19780
rect 27620 19728 27672 19780
rect 26240 19660 26292 19712
rect 26608 19660 26660 19712
rect 27528 19660 27580 19712
rect 34152 19728 34204 19780
rect 35348 19728 35400 19780
rect 36176 19728 36228 19780
rect 34704 19660 34756 19712
rect 35624 19660 35676 19712
rect 40592 19728 40644 19780
rect 43904 19796 43956 19848
rect 36544 19660 36596 19712
rect 40500 19660 40552 19712
rect 41052 19660 41104 19712
rect 42984 19728 43036 19780
rect 49148 19771 49200 19780
rect 49148 19737 49157 19771
rect 49157 19737 49191 19771
rect 49191 19737 49200 19771
rect 49148 19728 49200 19737
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 23388 19456 23440 19508
rect 28908 19456 28960 19508
rect 30104 19456 30156 19508
rect 33508 19456 33560 19508
rect 35164 19499 35216 19508
rect 35164 19465 35173 19499
rect 35173 19465 35207 19499
rect 35207 19465 35216 19499
rect 35164 19456 35216 19465
rect 27804 19388 27856 19440
rect 30932 19388 30984 19440
rect 32496 19431 32548 19440
rect 32496 19397 32505 19431
rect 32505 19397 32539 19431
rect 32539 19397 32548 19431
rect 32496 19388 32548 19397
rect 33968 19431 34020 19440
rect 33968 19397 33977 19431
rect 33977 19397 34011 19431
rect 34011 19397 34020 19431
rect 33968 19388 34020 19397
rect 34336 19388 34388 19440
rect 23296 19320 23348 19372
rect 25320 19320 25372 19372
rect 27436 19320 27488 19372
rect 28816 19320 28868 19372
rect 32772 19320 32824 19372
rect 24124 19295 24176 19304
rect 24124 19261 24133 19295
rect 24133 19261 24167 19295
rect 24167 19261 24176 19295
rect 24124 19252 24176 19261
rect 28724 19184 28776 19236
rect 29736 19252 29788 19304
rect 31760 19252 31812 19304
rect 34428 19320 34480 19372
rect 32220 19184 32272 19236
rect 33876 19184 33928 19236
rect 35348 19295 35400 19304
rect 35348 19261 35357 19295
rect 35357 19261 35391 19295
rect 35391 19261 35400 19295
rect 35348 19252 35400 19261
rect 43352 19320 43404 19372
rect 47952 19456 48004 19508
rect 43904 19431 43956 19440
rect 43904 19397 43913 19431
rect 43913 19397 43947 19431
rect 43947 19397 43956 19431
rect 43904 19388 43956 19397
rect 43812 19252 43864 19304
rect 46940 19252 46992 19304
rect 42984 19184 43036 19236
rect 43996 19184 44048 19236
rect 30380 19116 30432 19168
rect 32128 19116 32180 19168
rect 32864 19116 32916 19168
rect 37004 19116 37056 19168
rect 42340 19116 42392 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 22468 18912 22520 18964
rect 35072 18912 35124 18964
rect 29368 18844 29420 18896
rect 32128 18844 32180 18896
rect 25504 18776 25556 18828
rect 26240 18776 26292 18828
rect 29736 18776 29788 18828
rect 32588 18819 32640 18828
rect 32588 18785 32597 18819
rect 32597 18785 32631 18819
rect 32631 18785 32640 18819
rect 32588 18776 32640 18785
rect 32864 18819 32916 18828
rect 32864 18785 32873 18819
rect 32873 18785 32907 18819
rect 32907 18785 32916 18819
rect 32864 18776 32916 18785
rect 35256 18776 35308 18828
rect 35624 18912 35676 18964
rect 41788 18912 41840 18964
rect 27252 18708 27304 18760
rect 28724 18751 28776 18760
rect 28724 18717 28733 18751
rect 28733 18717 28767 18751
rect 28767 18717 28776 18751
rect 28724 18708 28776 18717
rect 31668 18708 31720 18760
rect 27436 18640 27488 18692
rect 32404 18640 32456 18692
rect 34428 18708 34480 18760
rect 37648 18776 37700 18828
rect 40868 18776 40920 18828
rect 41052 18819 41104 18828
rect 41052 18785 41061 18819
rect 41061 18785 41095 18819
rect 41095 18785 41104 18819
rect 41052 18776 41104 18785
rect 41420 18776 41472 18828
rect 38292 18708 38344 18760
rect 47952 18751 48004 18760
rect 47952 18717 47961 18751
rect 47961 18717 47995 18751
rect 47995 18717 48004 18751
rect 47952 18708 48004 18717
rect 49148 18751 49200 18760
rect 49148 18717 49157 18751
rect 49157 18717 49191 18751
rect 49191 18717 49200 18751
rect 49148 18708 49200 18717
rect 32864 18640 32916 18692
rect 34152 18640 34204 18692
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 26332 18572 26384 18624
rect 26424 18572 26476 18624
rect 34336 18615 34388 18624
rect 34336 18581 34345 18615
rect 34345 18581 34379 18615
rect 34379 18581 34388 18615
rect 34336 18572 34388 18581
rect 40408 18640 40460 18692
rect 43996 18640 44048 18692
rect 35256 18615 35308 18624
rect 35256 18581 35265 18615
rect 35265 18581 35299 18615
rect 35299 18581 35308 18615
rect 35256 18572 35308 18581
rect 35716 18572 35768 18624
rect 39488 18572 39540 18624
rect 40868 18615 40920 18624
rect 40868 18581 40877 18615
rect 40877 18581 40911 18615
rect 40911 18581 40920 18615
rect 40868 18572 40920 18581
rect 42892 18572 42944 18624
rect 43352 18572 43404 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 26056 18368 26108 18420
rect 28632 18411 28684 18420
rect 28632 18377 28641 18411
rect 28641 18377 28675 18411
rect 28675 18377 28684 18411
rect 28632 18368 28684 18377
rect 32312 18368 32364 18420
rect 35256 18368 35308 18420
rect 35532 18411 35584 18420
rect 35532 18377 35541 18411
rect 35541 18377 35575 18411
rect 35575 18377 35584 18411
rect 35532 18368 35584 18377
rect 38384 18368 38436 18420
rect 44364 18411 44416 18420
rect 44364 18377 44373 18411
rect 44373 18377 44407 18411
rect 44407 18377 44416 18411
rect 44364 18368 44416 18377
rect 23664 18232 23716 18284
rect 25044 18300 25096 18352
rect 25964 18232 26016 18284
rect 25228 18164 25280 18216
rect 27804 18207 27856 18216
rect 27804 18173 27813 18207
rect 27813 18173 27847 18207
rect 27847 18173 27856 18207
rect 27804 18164 27856 18173
rect 30196 18300 30248 18352
rect 30380 18300 30432 18352
rect 31024 18300 31076 18352
rect 31576 18300 31628 18352
rect 37648 18300 37700 18352
rect 42892 18343 42944 18352
rect 42892 18309 42901 18343
rect 42901 18309 42935 18343
rect 42935 18309 42944 18343
rect 42892 18300 42944 18309
rect 28448 18232 28500 18284
rect 29920 18232 29972 18284
rect 36268 18232 36320 18284
rect 38844 18232 38896 18284
rect 41144 18232 41196 18284
rect 41420 18232 41472 18284
rect 43996 18232 44048 18284
rect 29184 18207 29236 18216
rect 29184 18173 29193 18207
rect 29193 18173 29227 18207
rect 29227 18173 29236 18207
rect 29184 18164 29236 18173
rect 29736 18164 29788 18216
rect 34336 18164 34388 18216
rect 37464 18207 37516 18216
rect 37464 18173 37473 18207
rect 37473 18173 37507 18207
rect 37507 18173 37516 18207
rect 37464 18164 37516 18173
rect 25596 18071 25648 18080
rect 25596 18037 25605 18071
rect 25605 18037 25639 18071
rect 25639 18037 25648 18071
rect 25596 18028 25648 18037
rect 30472 18028 30524 18080
rect 32128 18028 32180 18080
rect 32588 18028 32640 18080
rect 40776 18164 40828 18216
rect 40868 18164 40920 18216
rect 43444 18164 43496 18216
rect 39948 18096 40000 18148
rect 49148 18207 49200 18216
rect 49148 18173 49157 18207
rect 49157 18173 49191 18207
rect 49191 18173 49200 18207
rect 49148 18164 49200 18173
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 25688 17824 25740 17876
rect 27620 17824 27672 17876
rect 28908 17824 28960 17876
rect 37096 17824 37148 17876
rect 43444 17824 43496 17876
rect 25228 17756 25280 17808
rect 25412 17731 25464 17740
rect 25412 17697 25421 17731
rect 25421 17697 25455 17731
rect 25455 17697 25464 17731
rect 25412 17688 25464 17697
rect 34152 17799 34204 17808
rect 34152 17765 34161 17799
rect 34161 17765 34195 17799
rect 34195 17765 34204 17799
rect 34152 17756 34204 17765
rect 27620 17688 27672 17740
rect 32036 17688 32088 17740
rect 28724 17620 28776 17672
rect 29000 17620 29052 17672
rect 33416 17620 33468 17672
rect 34520 17688 34572 17740
rect 42524 17756 42576 17808
rect 37372 17688 37424 17740
rect 38660 17688 38712 17740
rect 37004 17620 37056 17672
rect 40408 17620 40460 17672
rect 41328 17688 41380 17740
rect 49792 17756 49844 17808
rect 42800 17620 42852 17672
rect 49700 17688 49752 17740
rect 50068 17620 50120 17672
rect 27344 17552 27396 17604
rect 27712 17484 27764 17536
rect 33324 17552 33376 17604
rect 34060 17552 34112 17604
rect 36176 17552 36228 17604
rect 28356 17527 28408 17536
rect 28356 17493 28365 17527
rect 28365 17493 28399 17527
rect 28399 17493 28408 17527
rect 28356 17484 28408 17493
rect 28540 17484 28592 17536
rect 34888 17484 34940 17536
rect 43536 17484 43588 17536
rect 44548 17552 44600 17604
rect 45468 17595 45520 17604
rect 45468 17561 45477 17595
rect 45477 17561 45511 17595
rect 45511 17561 45520 17595
rect 45468 17552 45520 17561
rect 49424 17484 49476 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 25136 17280 25188 17332
rect 25596 17280 25648 17332
rect 25964 17280 26016 17332
rect 27160 17212 27212 17264
rect 28540 17280 28592 17332
rect 31760 17280 31812 17332
rect 29184 17212 29236 17264
rect 32036 17212 32088 17264
rect 33416 17323 33468 17332
rect 33416 17289 33425 17323
rect 33425 17289 33459 17323
rect 33459 17289 33468 17323
rect 33416 17280 33468 17289
rect 37464 17280 37516 17332
rect 38568 17280 38620 17332
rect 39672 17280 39724 17332
rect 37004 17212 37056 17264
rect 20996 17144 21048 17196
rect 19800 17076 19852 17128
rect 26240 17144 26292 17196
rect 24860 17076 24912 17128
rect 29460 17144 29512 17196
rect 30748 17144 30800 17196
rect 30932 17187 30984 17196
rect 30932 17153 30941 17187
rect 30941 17153 30975 17187
rect 30975 17153 30984 17187
rect 30932 17144 30984 17153
rect 32128 17144 32180 17196
rect 27804 17076 27856 17128
rect 28540 17119 28592 17128
rect 28540 17085 28549 17119
rect 28549 17085 28583 17119
rect 28583 17085 28592 17119
rect 28540 17076 28592 17085
rect 28632 17076 28684 17128
rect 27712 17008 27764 17060
rect 28724 17008 28776 17060
rect 30380 17076 30432 17128
rect 38844 17144 38896 17196
rect 40408 17212 40460 17264
rect 42892 17212 42944 17264
rect 39672 17187 39724 17196
rect 39672 17153 39681 17187
rect 39681 17153 39715 17187
rect 39715 17153 39724 17187
rect 39672 17144 39724 17153
rect 44088 17280 44140 17332
rect 44272 17255 44324 17264
rect 44272 17221 44281 17255
rect 44281 17221 44315 17255
rect 44315 17221 44324 17255
rect 44272 17212 44324 17221
rect 45560 17144 45612 17196
rect 37740 17119 37792 17128
rect 37740 17085 37749 17119
rect 37749 17085 37783 17119
rect 37783 17085 37792 17119
rect 37740 17076 37792 17085
rect 37832 17076 37884 17128
rect 39948 17119 40000 17128
rect 39948 17085 39957 17119
rect 39957 17085 39991 17119
rect 39991 17085 40000 17119
rect 39948 17076 40000 17085
rect 40408 17076 40460 17128
rect 39028 17008 39080 17060
rect 29092 16983 29144 16992
rect 29092 16949 29101 16983
rect 29101 16949 29135 16983
rect 29135 16949 29144 16983
rect 29092 16940 29144 16949
rect 31760 16983 31812 16992
rect 31760 16949 31769 16983
rect 31769 16949 31803 16983
rect 31803 16949 31812 16983
rect 31760 16940 31812 16949
rect 41052 17008 41104 17060
rect 43352 17076 43404 17128
rect 49148 17119 49200 17128
rect 49148 17085 49157 17119
rect 49157 17085 49191 17119
rect 49191 17085 49200 17119
rect 49148 17076 49200 17085
rect 43996 17008 44048 17060
rect 46112 16940 46164 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 20996 16779 21048 16788
rect 20996 16745 21005 16779
rect 21005 16745 21039 16779
rect 21039 16745 21048 16779
rect 20996 16736 21048 16745
rect 23848 16736 23900 16788
rect 25228 16736 25280 16788
rect 29184 16736 29236 16788
rect 31944 16736 31996 16788
rect 35808 16736 35860 16788
rect 41328 16736 41380 16788
rect 23572 16600 23624 16652
rect 29092 16668 29144 16720
rect 33968 16668 34020 16720
rect 37832 16668 37884 16720
rect 25688 16643 25740 16652
rect 25688 16609 25697 16643
rect 25697 16609 25731 16643
rect 25731 16609 25740 16643
rect 25688 16600 25740 16609
rect 27160 16643 27212 16652
rect 27160 16609 27169 16643
rect 27169 16609 27203 16643
rect 27203 16609 27212 16643
rect 27160 16600 27212 16609
rect 27528 16600 27580 16652
rect 27620 16600 27672 16652
rect 28632 16643 28684 16652
rect 28632 16609 28641 16643
rect 28641 16609 28675 16643
rect 28675 16609 28684 16643
rect 28632 16600 28684 16609
rect 29644 16600 29696 16652
rect 29736 16643 29788 16652
rect 29736 16609 29745 16643
rect 29745 16609 29779 16643
rect 29779 16609 29788 16643
rect 29736 16600 29788 16609
rect 25780 16532 25832 16584
rect 26516 16532 26568 16584
rect 29000 16532 29052 16584
rect 31024 16532 31076 16584
rect 24768 16464 24820 16516
rect 24124 16396 24176 16448
rect 26792 16464 26844 16516
rect 27344 16464 27396 16516
rect 29644 16464 29696 16516
rect 26700 16439 26752 16448
rect 26700 16405 26709 16439
rect 26709 16405 26743 16439
rect 26743 16405 26752 16439
rect 26700 16396 26752 16405
rect 27068 16439 27120 16448
rect 27068 16405 27077 16439
rect 27077 16405 27111 16439
rect 27111 16405 27120 16439
rect 27068 16396 27120 16405
rect 29276 16396 29328 16448
rect 30380 16396 30432 16448
rect 31944 16643 31996 16652
rect 31944 16609 31953 16643
rect 31953 16609 31987 16643
rect 31987 16609 31996 16643
rect 31944 16600 31996 16609
rect 34336 16600 34388 16652
rect 36728 16600 36780 16652
rect 38476 16643 38528 16652
rect 38476 16609 38485 16643
rect 38485 16609 38519 16643
rect 38519 16609 38528 16643
rect 38476 16600 38528 16609
rect 39948 16600 40000 16652
rect 42616 16600 42668 16652
rect 46112 16600 46164 16652
rect 33324 16532 33376 16584
rect 35072 16532 35124 16584
rect 32128 16464 32180 16516
rect 32864 16396 32916 16448
rect 32956 16396 33008 16448
rect 35440 16464 35492 16516
rect 37188 16532 37240 16584
rect 40316 16532 40368 16584
rect 44456 16532 44508 16584
rect 36912 16464 36964 16516
rect 37372 16464 37424 16516
rect 33876 16396 33928 16448
rect 35532 16396 35584 16448
rect 40500 16464 40552 16516
rect 42800 16464 42852 16516
rect 49148 16507 49200 16516
rect 49148 16473 49157 16507
rect 49157 16473 49191 16507
rect 49191 16473 49200 16507
rect 49148 16464 49200 16473
rect 40040 16439 40092 16448
rect 40040 16405 40049 16439
rect 40049 16405 40083 16439
rect 40083 16405 40092 16439
rect 40040 16396 40092 16405
rect 40224 16396 40276 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 27712 16192 27764 16244
rect 28264 16192 28316 16244
rect 31760 16192 31812 16244
rect 24124 16124 24176 16176
rect 23572 15988 23624 16040
rect 24492 16031 24544 16040
rect 24492 15997 24501 16031
rect 24501 15997 24535 16031
rect 24535 15997 24544 16031
rect 24492 15988 24544 15997
rect 24768 15988 24820 16040
rect 27344 16124 27396 16176
rect 29644 16124 29696 16176
rect 31024 16124 31076 16176
rect 34520 16192 34572 16244
rect 34796 16192 34848 16244
rect 35072 16124 35124 16176
rect 36176 16124 36228 16176
rect 37556 16056 37608 16108
rect 39396 16056 39448 16108
rect 40776 16099 40828 16108
rect 40776 16065 40785 16099
rect 40785 16065 40819 16099
rect 40819 16065 40828 16099
rect 40776 16056 40828 16065
rect 27528 15988 27580 16040
rect 27712 15988 27764 16040
rect 28724 15988 28776 16040
rect 28908 15988 28960 16040
rect 30472 15988 30524 16040
rect 32036 15988 32088 16040
rect 32956 16031 33008 16040
rect 32956 15997 32965 16031
rect 32965 15997 32999 16031
rect 32999 15997 33008 16031
rect 32956 15988 33008 15997
rect 34796 15988 34848 16040
rect 35992 15920 36044 15972
rect 37556 15852 37608 15904
rect 38292 15852 38344 15904
rect 42708 15852 42760 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 23296 15691 23348 15700
rect 23296 15657 23305 15691
rect 23305 15657 23339 15691
rect 23339 15657 23348 15691
rect 23296 15648 23348 15657
rect 26976 15648 27028 15700
rect 31576 15648 31628 15700
rect 37740 15648 37792 15700
rect 23848 15555 23900 15564
rect 23848 15521 23857 15555
rect 23857 15521 23891 15555
rect 23891 15521 23900 15555
rect 23848 15512 23900 15521
rect 24492 15512 24544 15564
rect 26240 15512 26292 15564
rect 28264 15512 28316 15564
rect 31668 15555 31720 15564
rect 31668 15521 31677 15555
rect 31677 15521 31711 15555
rect 31711 15521 31720 15555
rect 31668 15512 31720 15521
rect 34520 15512 34572 15564
rect 35624 15555 35676 15564
rect 35624 15521 35633 15555
rect 35633 15521 35667 15555
rect 35667 15521 35676 15555
rect 35624 15512 35676 15521
rect 35900 15555 35952 15564
rect 35900 15521 35909 15555
rect 35909 15521 35943 15555
rect 35943 15521 35952 15555
rect 35900 15512 35952 15521
rect 40868 15580 40920 15632
rect 45560 15580 45612 15632
rect 28724 15444 28776 15496
rect 30656 15487 30708 15496
rect 30656 15453 30665 15487
rect 30665 15453 30699 15487
rect 30699 15453 30708 15487
rect 30656 15444 30708 15453
rect 34244 15444 34296 15496
rect 37280 15444 37332 15496
rect 43628 15444 43680 15496
rect 44732 15444 44784 15496
rect 49148 15487 49200 15496
rect 49148 15453 49157 15487
rect 49157 15453 49191 15487
rect 49191 15453 49200 15487
rect 49148 15444 49200 15453
rect 23388 15376 23440 15428
rect 25504 15419 25556 15428
rect 25504 15385 25513 15419
rect 25513 15385 25547 15419
rect 25547 15385 25556 15419
rect 25504 15376 25556 15385
rect 27344 15376 27396 15428
rect 29552 15376 29604 15428
rect 30840 15376 30892 15428
rect 33508 15376 33560 15428
rect 25872 15308 25924 15360
rect 29828 15308 29880 15360
rect 33692 15351 33744 15360
rect 33692 15317 33701 15351
rect 33701 15317 33735 15351
rect 33735 15317 33744 15351
rect 33692 15308 33744 15317
rect 36360 15376 36412 15428
rect 37464 15376 37516 15428
rect 38660 15376 38712 15428
rect 42524 15308 42576 15360
rect 47768 15376 47820 15428
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 25504 15104 25556 15156
rect 23572 15036 23624 15088
rect 26240 15036 26292 15088
rect 30656 15104 30708 15156
rect 24768 14968 24820 15020
rect 27436 14968 27488 15020
rect 27528 14968 27580 15020
rect 31944 15036 31996 15088
rect 32864 15104 32916 15156
rect 34520 15104 34572 15156
rect 38660 15104 38712 15156
rect 25504 14900 25556 14952
rect 32128 14968 32180 15020
rect 33324 15036 33376 15088
rect 25044 14832 25096 14884
rect 28264 14807 28316 14816
rect 28264 14773 28273 14807
rect 28273 14773 28307 14807
rect 28307 14773 28316 14807
rect 30288 14900 30340 14952
rect 30564 14943 30616 14952
rect 30564 14909 30573 14943
rect 30573 14909 30607 14943
rect 30607 14909 30616 14943
rect 30564 14900 30616 14909
rect 31852 14900 31904 14952
rect 34980 15036 35032 15088
rect 35348 15036 35400 15088
rect 35624 15079 35676 15088
rect 35624 15045 35633 15079
rect 35633 15045 35667 15079
rect 35667 15045 35676 15079
rect 35624 15036 35676 15045
rect 36544 15036 36596 15088
rect 39028 15079 39080 15088
rect 39028 15045 39037 15079
rect 39037 15045 39071 15079
rect 39071 15045 39080 15079
rect 39028 15036 39080 15045
rect 40408 15036 40460 15088
rect 32312 14832 32364 14884
rect 28264 14764 28316 14773
rect 30748 14764 30800 14816
rect 32404 14764 32456 14816
rect 36268 14968 36320 15020
rect 37280 14968 37332 15020
rect 38568 14968 38620 15020
rect 43536 14968 43588 15020
rect 47952 15011 48004 15020
rect 47952 14977 47961 15011
rect 47961 14977 47995 15011
rect 47995 14977 48004 15011
rect 47952 14968 48004 14977
rect 34060 14943 34112 14952
rect 34060 14909 34069 14943
rect 34069 14909 34103 14943
rect 34103 14909 34112 14943
rect 34060 14900 34112 14909
rect 49148 14943 49200 14952
rect 49148 14909 49157 14943
rect 49157 14909 49191 14943
rect 49191 14909 49200 14943
rect 49148 14900 49200 14909
rect 36452 14807 36504 14816
rect 36452 14773 36461 14807
rect 36461 14773 36495 14807
rect 36495 14773 36504 14807
rect 36452 14764 36504 14773
rect 39396 14764 39448 14816
rect 47860 14764 47912 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 25320 14560 25372 14612
rect 28448 14603 28500 14612
rect 28448 14569 28457 14603
rect 28457 14569 28491 14603
rect 28491 14569 28500 14603
rect 28448 14560 28500 14569
rect 30288 14560 30340 14612
rect 31484 14560 31536 14612
rect 32128 14560 32180 14612
rect 35348 14560 35400 14612
rect 30196 14492 30248 14544
rect 35072 14492 35124 14544
rect 41236 14492 41288 14544
rect 47952 14560 48004 14612
rect 49240 14492 49292 14544
rect 23848 14424 23900 14476
rect 26792 14424 26844 14476
rect 27712 14424 27764 14476
rect 28908 14424 28960 14476
rect 31484 14424 31536 14476
rect 34796 14424 34848 14476
rect 38568 14424 38620 14476
rect 39212 14467 39264 14476
rect 39212 14433 39221 14467
rect 39221 14433 39255 14467
rect 39255 14433 39264 14467
rect 39212 14424 39264 14433
rect 39396 14467 39448 14476
rect 39396 14433 39405 14467
rect 39405 14433 39439 14467
rect 39439 14433 39448 14467
rect 39396 14424 39448 14433
rect 26240 14356 26292 14408
rect 26976 14399 27028 14408
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 27436 14399 27488 14408
rect 27436 14365 27445 14399
rect 27445 14365 27479 14399
rect 27479 14365 27488 14399
rect 27436 14356 27488 14365
rect 28448 14356 28500 14408
rect 28816 14356 28868 14408
rect 30932 14356 30984 14408
rect 32036 14399 32088 14408
rect 32036 14365 32045 14399
rect 32045 14365 32079 14399
rect 32079 14365 32088 14399
rect 32036 14356 32088 14365
rect 39120 14356 39172 14408
rect 27344 14288 27396 14340
rect 26516 14220 26568 14272
rect 26608 14263 26660 14272
rect 26608 14229 26617 14263
rect 26617 14229 26651 14263
rect 26651 14229 26660 14263
rect 26608 14220 26660 14229
rect 26884 14220 26936 14272
rect 28816 14263 28868 14272
rect 28816 14229 28825 14263
rect 28825 14229 28859 14263
rect 28859 14229 28868 14263
rect 28816 14220 28868 14229
rect 28908 14263 28960 14272
rect 28908 14229 28917 14263
rect 28917 14229 28951 14263
rect 28951 14229 28960 14263
rect 28908 14220 28960 14229
rect 30932 14220 30984 14272
rect 31576 14263 31628 14272
rect 31576 14229 31585 14263
rect 31585 14229 31619 14263
rect 31619 14229 31628 14263
rect 31576 14220 31628 14229
rect 31852 14288 31904 14340
rect 34704 14288 34756 14340
rect 35624 14263 35676 14272
rect 35624 14229 35633 14263
rect 35633 14229 35667 14263
rect 35667 14229 35676 14263
rect 35624 14220 35676 14229
rect 35900 14288 35952 14340
rect 36268 14288 36320 14340
rect 41144 14424 41196 14476
rect 41328 14424 41380 14476
rect 50528 14424 50580 14476
rect 41236 14399 41288 14408
rect 41236 14365 41245 14399
rect 41245 14365 41279 14399
rect 41279 14365 41288 14399
rect 41236 14356 41288 14365
rect 42156 14288 42208 14340
rect 38752 14263 38804 14272
rect 38752 14229 38761 14263
rect 38761 14229 38795 14263
rect 38795 14229 38804 14263
rect 38752 14220 38804 14229
rect 38844 14220 38896 14272
rect 40960 14220 41012 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 23480 14016 23532 14068
rect 23756 14016 23808 14068
rect 23848 14016 23900 14068
rect 25872 14059 25924 14068
rect 25872 14025 25881 14059
rect 25881 14025 25915 14059
rect 25915 14025 25924 14059
rect 25872 14016 25924 14025
rect 26240 14059 26292 14068
rect 26240 14025 26249 14059
rect 26249 14025 26283 14059
rect 26283 14025 26292 14059
rect 26240 14016 26292 14025
rect 28172 14016 28224 14068
rect 29920 14016 29972 14068
rect 32128 14016 32180 14068
rect 33324 14016 33376 14068
rect 24768 13948 24820 14000
rect 25320 13948 25372 14000
rect 26240 13880 26292 13932
rect 27528 13880 27580 13932
rect 29644 13948 29696 14000
rect 27712 13923 27764 13932
rect 33416 13948 33468 14000
rect 34796 14016 34848 14068
rect 35072 14016 35124 14068
rect 37924 14059 37976 14068
rect 37924 14025 37933 14059
rect 37933 14025 37967 14059
rect 37967 14025 37976 14059
rect 37924 14016 37976 14025
rect 38752 14016 38804 14068
rect 42432 14016 42484 14068
rect 44456 14016 44508 14068
rect 34520 13948 34572 14000
rect 35256 13948 35308 14000
rect 27712 13889 27728 13923
rect 27728 13889 27762 13923
rect 27762 13889 27764 13923
rect 27712 13880 27764 13889
rect 20076 13676 20128 13728
rect 20352 13676 20404 13728
rect 26424 13744 26476 13796
rect 28540 13812 28592 13864
rect 28724 13812 28776 13864
rect 30472 13812 30524 13864
rect 32864 13923 32916 13932
rect 32864 13889 32873 13923
rect 32873 13889 32907 13923
rect 32907 13889 32916 13923
rect 32864 13880 32916 13889
rect 37372 13948 37424 14000
rect 39396 13948 39448 14000
rect 42708 13948 42760 14000
rect 32680 13812 32732 13864
rect 27252 13744 27304 13796
rect 23480 13676 23532 13728
rect 24676 13676 24728 13728
rect 26792 13676 26844 13728
rect 27528 13676 27580 13728
rect 28080 13676 28132 13728
rect 28172 13676 28224 13728
rect 28540 13676 28592 13728
rect 29368 13676 29420 13728
rect 29460 13719 29512 13728
rect 29460 13685 29469 13719
rect 29469 13685 29503 13719
rect 29503 13685 29512 13719
rect 32864 13744 32916 13796
rect 35256 13812 35308 13864
rect 29460 13676 29512 13685
rect 32404 13676 32456 13728
rect 38568 13880 38620 13932
rect 39028 13923 39080 13932
rect 39028 13889 39037 13923
rect 39037 13889 39071 13923
rect 39071 13889 39080 13923
rect 39028 13880 39080 13889
rect 40408 13880 40460 13932
rect 40592 13880 40644 13932
rect 43352 13923 43404 13932
rect 43352 13889 43361 13923
rect 43361 13889 43395 13923
rect 43395 13889 43404 13923
rect 43352 13880 43404 13889
rect 47768 13880 47820 13932
rect 40684 13812 40736 13864
rect 45928 13855 45980 13864
rect 45928 13821 45937 13855
rect 45937 13821 45971 13855
rect 45971 13821 45980 13855
rect 45928 13812 45980 13821
rect 49148 13855 49200 13864
rect 49148 13821 49157 13855
rect 49157 13821 49191 13855
rect 49191 13821 49200 13855
rect 49148 13812 49200 13821
rect 37648 13676 37700 13728
rect 40776 13719 40828 13728
rect 40776 13685 40785 13719
rect 40785 13685 40819 13719
rect 40819 13685 40828 13719
rect 40776 13676 40828 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 20352 13472 20404 13524
rect 20076 13311 20128 13320
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 18604 13175 18656 13184
rect 18604 13141 18613 13175
rect 18613 13141 18647 13175
rect 18647 13141 18656 13175
rect 18604 13132 18656 13141
rect 24952 13515 25004 13524
rect 24952 13481 24961 13515
rect 24961 13481 24995 13515
rect 24995 13481 25004 13515
rect 24952 13472 25004 13481
rect 26332 13472 26384 13524
rect 26792 13472 26844 13524
rect 28448 13472 28500 13524
rect 29644 13472 29696 13524
rect 31024 13472 31076 13524
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 26424 13404 26476 13456
rect 27528 13404 27580 13456
rect 30012 13404 30064 13456
rect 25504 13379 25556 13388
rect 25504 13345 25513 13379
rect 25513 13345 25547 13379
rect 25547 13345 25556 13379
rect 25504 13336 25556 13345
rect 28080 13336 28132 13388
rect 30380 13336 30432 13388
rect 30840 13379 30892 13388
rect 30840 13345 30849 13379
rect 30849 13345 30883 13379
rect 30883 13345 30892 13379
rect 30840 13336 30892 13345
rect 26792 13268 26844 13320
rect 26884 13268 26936 13320
rect 30656 13268 30708 13320
rect 32312 13472 32364 13524
rect 37096 13472 37148 13524
rect 37188 13472 37240 13524
rect 38660 13472 38712 13524
rect 48780 13472 48832 13524
rect 35624 13404 35676 13456
rect 44640 13404 44692 13456
rect 23296 13200 23348 13252
rect 24860 13200 24912 13252
rect 27804 13200 27856 13252
rect 31760 13268 31812 13320
rect 32404 13379 32456 13388
rect 32404 13345 32413 13379
rect 32413 13345 32447 13379
rect 32447 13345 32456 13379
rect 32404 13336 32456 13345
rect 32864 13336 32916 13388
rect 36268 13336 36320 13388
rect 39028 13336 39080 13388
rect 33416 13268 33468 13320
rect 24032 13132 24084 13184
rect 25412 13175 25464 13184
rect 25412 13141 25421 13175
rect 25421 13141 25455 13175
rect 25455 13141 25464 13175
rect 25412 13132 25464 13141
rect 26424 13132 26476 13184
rect 26700 13132 26752 13184
rect 26976 13175 27028 13184
rect 26976 13141 26985 13175
rect 26985 13141 27019 13175
rect 27019 13141 27028 13175
rect 26976 13132 27028 13141
rect 28080 13132 28132 13184
rect 35164 13268 35216 13320
rect 35808 13268 35860 13320
rect 39488 13311 39540 13320
rect 39488 13277 39497 13311
rect 39497 13277 39531 13311
rect 39531 13277 39540 13311
rect 39488 13268 39540 13277
rect 42340 13336 42392 13388
rect 44732 13336 44784 13388
rect 40500 13268 40552 13320
rect 44364 13268 44416 13320
rect 47860 13268 47912 13320
rect 28264 13132 28316 13184
rect 29644 13132 29696 13184
rect 30380 13175 30432 13184
rect 30380 13141 30389 13175
rect 30389 13141 30423 13175
rect 30423 13141 30432 13175
rect 30380 13132 30432 13141
rect 34888 13200 34940 13252
rect 35992 13200 36044 13252
rect 33784 13132 33836 13184
rect 37280 13200 37332 13252
rect 49148 13243 49200 13252
rect 49148 13209 49157 13243
rect 49157 13209 49191 13243
rect 49191 13209 49200 13243
rect 49148 13200 49200 13209
rect 37740 13132 37792 13184
rect 39212 13132 39264 13184
rect 40500 13132 40552 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 17224 12928 17276 12980
rect 21456 12928 21508 12980
rect 23388 12928 23440 12980
rect 23296 12903 23348 12912
rect 23296 12869 23305 12903
rect 23305 12869 23339 12903
rect 23339 12869 23348 12903
rect 23296 12860 23348 12869
rect 25320 12928 25372 12980
rect 27344 12928 27396 12980
rect 30380 12928 30432 12980
rect 24860 12860 24912 12912
rect 29092 12860 29144 12912
rect 31576 12928 31628 12980
rect 32772 12971 32824 12980
rect 32772 12937 32781 12971
rect 32781 12937 32815 12971
rect 32815 12937 32824 12971
rect 32772 12928 32824 12937
rect 31024 12860 31076 12912
rect 32312 12860 32364 12912
rect 35348 12903 35400 12912
rect 35348 12869 35357 12903
rect 35357 12869 35391 12903
rect 35391 12869 35400 12903
rect 35348 12860 35400 12869
rect 36820 12860 36872 12912
rect 27252 12792 27304 12844
rect 23480 12767 23532 12776
rect 23480 12733 23489 12767
rect 23489 12733 23523 12767
rect 23523 12733 23532 12767
rect 23480 12724 23532 12733
rect 24768 12724 24820 12776
rect 24860 12724 24912 12776
rect 25136 12724 25188 12776
rect 26700 12724 26752 12776
rect 27896 12724 27948 12776
rect 29920 12792 29972 12844
rect 28080 12724 28132 12776
rect 26608 12656 26660 12708
rect 26976 12656 27028 12708
rect 29368 12767 29420 12776
rect 29368 12733 29377 12767
rect 29377 12733 29411 12767
rect 29411 12733 29420 12767
rect 29368 12724 29420 12733
rect 29736 12724 29788 12776
rect 30380 12724 30432 12776
rect 34060 12792 34112 12844
rect 48596 12928 48648 12980
rect 33968 12724 34020 12776
rect 25504 12588 25556 12640
rect 27804 12588 27856 12640
rect 28356 12588 28408 12640
rect 28632 12588 28684 12640
rect 29000 12588 29052 12640
rect 33876 12656 33928 12708
rect 34704 12656 34756 12708
rect 31760 12631 31812 12640
rect 31760 12597 31769 12631
rect 31769 12597 31803 12631
rect 31803 12597 31812 12631
rect 31760 12588 31812 12597
rect 32312 12631 32364 12640
rect 32312 12597 32321 12631
rect 32321 12597 32355 12631
rect 32355 12597 32364 12631
rect 32312 12588 32364 12597
rect 33692 12631 33744 12640
rect 33692 12597 33701 12631
rect 33701 12597 33735 12631
rect 33735 12597 33744 12631
rect 33692 12588 33744 12597
rect 34796 12631 34848 12640
rect 34796 12597 34805 12631
rect 34805 12597 34839 12631
rect 34839 12597 34848 12631
rect 34796 12588 34848 12597
rect 34980 12656 35032 12708
rect 38660 12792 38712 12844
rect 39028 12792 39080 12844
rect 40592 12792 40644 12844
rect 40868 12792 40920 12844
rect 40776 12724 40828 12776
rect 37648 12631 37700 12640
rect 37648 12597 37657 12631
rect 37657 12597 37691 12631
rect 37691 12597 37700 12631
rect 37648 12588 37700 12597
rect 40224 12588 40276 12640
rect 40684 12588 40736 12640
rect 44180 12588 44232 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 25412 12384 25464 12436
rect 27068 12384 27120 12436
rect 24768 12316 24820 12368
rect 25044 12291 25096 12300
rect 25044 12257 25053 12291
rect 25053 12257 25087 12291
rect 25087 12257 25096 12291
rect 25044 12248 25096 12257
rect 24584 12180 24636 12232
rect 27620 12316 27672 12368
rect 29552 12384 29604 12436
rect 31852 12384 31904 12436
rect 32496 12384 32548 12436
rect 33508 12384 33560 12436
rect 28172 12316 28224 12368
rect 28724 12316 28776 12368
rect 31760 12316 31812 12368
rect 28448 12248 28500 12300
rect 30288 12291 30340 12300
rect 30288 12257 30297 12291
rect 30297 12257 30331 12291
rect 30331 12257 30340 12291
rect 30288 12248 30340 12257
rect 28724 12180 28776 12232
rect 30104 12223 30156 12232
rect 30104 12189 30113 12223
rect 30113 12189 30147 12223
rect 30147 12189 30156 12223
rect 32220 12248 32272 12300
rect 32496 12291 32548 12300
rect 32496 12257 32505 12291
rect 32505 12257 32539 12291
rect 32539 12257 32548 12291
rect 32496 12248 32548 12257
rect 36176 12384 36228 12436
rect 37188 12384 37240 12436
rect 37740 12384 37792 12436
rect 35164 12248 35216 12300
rect 30104 12180 30156 12189
rect 28264 12112 28316 12164
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 26148 12044 26200 12096
rect 33692 12112 33744 12164
rect 33876 12112 33928 12164
rect 36268 12291 36320 12300
rect 36268 12257 36277 12291
rect 36277 12257 36311 12291
rect 36311 12257 36320 12291
rect 36268 12248 36320 12257
rect 39304 12223 39356 12232
rect 39304 12189 39313 12223
rect 39313 12189 39347 12223
rect 39347 12189 39356 12223
rect 39304 12180 39356 12189
rect 41052 12180 41104 12232
rect 45928 12180 45980 12232
rect 49148 12223 49200 12232
rect 49148 12189 49157 12223
rect 49157 12189 49191 12223
rect 49191 12189 49200 12223
rect 49148 12180 49200 12189
rect 36636 12112 36688 12164
rect 37280 12112 37332 12164
rect 37832 12112 37884 12164
rect 43352 12112 43404 12164
rect 30196 12087 30248 12096
rect 30196 12053 30205 12087
rect 30205 12053 30239 12087
rect 30239 12053 30248 12087
rect 30196 12044 30248 12053
rect 30380 12044 30432 12096
rect 30656 12044 30708 12096
rect 31116 12044 31168 12096
rect 38292 12044 38344 12096
rect 38476 12087 38528 12096
rect 38476 12053 38485 12087
rect 38485 12053 38519 12087
rect 38519 12053 38528 12087
rect 38476 12044 38528 12053
rect 40868 12044 40920 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 23480 11840 23532 11892
rect 26516 11840 26568 11892
rect 28356 11883 28408 11892
rect 28356 11849 28365 11883
rect 28365 11849 28399 11883
rect 28399 11849 28408 11883
rect 28356 11840 28408 11849
rect 28724 11883 28776 11892
rect 28724 11849 28733 11883
rect 28733 11849 28767 11883
rect 28767 11849 28776 11883
rect 28724 11840 28776 11849
rect 29828 11840 29880 11892
rect 27252 11772 27304 11824
rect 29552 11772 29604 11824
rect 25136 11704 25188 11756
rect 26608 11704 26660 11756
rect 23756 11679 23808 11688
rect 23756 11645 23765 11679
rect 23765 11645 23799 11679
rect 23799 11645 23808 11679
rect 23756 11636 23808 11645
rect 24032 11679 24084 11688
rect 24032 11645 24041 11679
rect 24041 11645 24075 11679
rect 24075 11645 24084 11679
rect 24032 11636 24084 11645
rect 24676 11636 24728 11688
rect 29276 11704 29328 11756
rect 29092 11636 29144 11688
rect 29368 11636 29420 11688
rect 29184 11568 29236 11620
rect 30380 11772 30432 11824
rect 31668 11840 31720 11892
rect 33876 11840 33928 11892
rect 34796 11840 34848 11892
rect 37832 11840 37884 11892
rect 39304 11840 39356 11892
rect 40592 11883 40644 11892
rect 40592 11849 40601 11883
rect 40601 11849 40635 11883
rect 40635 11849 40644 11883
rect 40592 11840 40644 11849
rect 34704 11772 34756 11824
rect 30288 11747 30340 11756
rect 30288 11713 30297 11747
rect 30297 11713 30331 11747
rect 30331 11713 30340 11747
rect 30288 11704 30340 11713
rect 30380 11679 30432 11688
rect 30380 11645 30389 11679
rect 30389 11645 30423 11679
rect 30423 11645 30432 11679
rect 31760 11704 31812 11756
rect 36820 11772 36872 11824
rect 38292 11815 38344 11824
rect 38292 11781 38301 11815
rect 38301 11781 38335 11815
rect 38335 11781 38344 11815
rect 38292 11772 38344 11781
rect 38476 11772 38528 11824
rect 30380 11636 30432 11645
rect 33508 11636 33560 11688
rect 35256 11568 35308 11620
rect 24768 11500 24820 11552
rect 27620 11500 27672 11552
rect 32496 11500 32548 11552
rect 36268 11747 36320 11756
rect 36268 11713 36277 11747
rect 36277 11713 36311 11747
rect 36311 11713 36320 11747
rect 36268 11704 36320 11713
rect 37740 11704 37792 11756
rect 37924 11636 37976 11688
rect 38568 11704 38620 11756
rect 39120 11747 39172 11756
rect 39120 11713 39129 11747
rect 39129 11713 39163 11747
rect 39163 11713 39172 11747
rect 39120 11704 39172 11713
rect 42432 11704 42484 11756
rect 40684 11679 40736 11688
rect 40684 11645 40693 11679
rect 40693 11645 40727 11679
rect 40727 11645 40736 11679
rect 40684 11636 40736 11645
rect 38936 11500 38988 11552
rect 43720 11636 43772 11688
rect 42800 11568 42852 11620
rect 49148 11679 49200 11688
rect 49148 11645 49157 11679
rect 49157 11645 49191 11679
rect 49191 11645 49200 11679
rect 49148 11636 49200 11645
rect 45192 11500 45244 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 13360 11296 13412 11348
rect 24584 11296 24636 11348
rect 24860 11296 24912 11348
rect 19984 11228 20036 11280
rect 28816 11296 28868 11348
rect 29644 11296 29696 11348
rect 29920 11296 29972 11348
rect 32128 11339 32180 11348
rect 32128 11305 32137 11339
rect 32137 11305 32171 11339
rect 32171 11305 32180 11339
rect 32128 11296 32180 11305
rect 29092 11228 29144 11280
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 26240 11160 26292 11212
rect 28632 11160 28684 11212
rect 29828 11160 29880 11212
rect 32312 11228 32364 11280
rect 32588 11228 32640 11280
rect 34520 11228 34572 11280
rect 31576 11203 31628 11212
rect 31576 11169 31585 11203
rect 31585 11169 31619 11203
rect 31619 11169 31628 11203
rect 31576 11160 31628 11169
rect 32772 11203 32824 11212
rect 32772 11169 32781 11203
rect 32781 11169 32815 11203
rect 32815 11169 32824 11203
rect 32772 11160 32824 11169
rect 35164 11160 35216 11212
rect 29644 11092 29696 11144
rect 30564 11092 30616 11144
rect 31116 11092 31168 11144
rect 31392 11092 31444 11144
rect 32312 11092 32364 11144
rect 35900 11092 35952 11144
rect 26608 11024 26660 11076
rect 29920 11024 29972 11076
rect 31944 11024 31996 11076
rect 32588 11067 32640 11076
rect 32588 11033 32597 11067
rect 32597 11033 32631 11067
rect 32631 11033 32640 11067
rect 32588 11024 32640 11033
rect 34060 11024 34112 11076
rect 35256 11067 35308 11076
rect 35256 11033 35265 11067
rect 35265 11033 35299 11067
rect 35299 11033 35308 11067
rect 35256 11024 35308 11033
rect 35348 11067 35400 11076
rect 35348 11033 35357 11067
rect 35357 11033 35391 11067
rect 35391 11033 35400 11067
rect 35348 11024 35400 11033
rect 37004 11067 37056 11076
rect 37004 11033 37013 11067
rect 37013 11033 37047 11067
rect 37047 11033 37056 11067
rect 37004 11024 37056 11033
rect 44364 11296 44416 11348
rect 37924 11228 37976 11280
rect 38844 11228 38896 11280
rect 39488 11160 39540 11212
rect 40960 11160 41012 11212
rect 37832 11135 37884 11144
rect 37832 11101 37841 11135
rect 37841 11101 37875 11135
rect 37875 11101 37884 11135
rect 37832 11092 37884 11101
rect 38660 11135 38712 11144
rect 38660 11101 38669 11135
rect 38669 11101 38703 11135
rect 38703 11101 38712 11135
rect 38660 11092 38712 11101
rect 38936 11092 38988 11144
rect 38844 11067 38896 11076
rect 38844 11033 38853 11067
rect 38853 11033 38887 11067
rect 38887 11033 38896 11067
rect 38844 11024 38896 11033
rect 29000 10956 29052 11008
rect 31116 10956 31168 11008
rect 31576 10956 31628 11008
rect 32128 10956 32180 11008
rect 37556 10956 37608 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 27160 10752 27212 10804
rect 29552 10795 29604 10804
rect 29552 10761 29561 10795
rect 29561 10761 29595 10795
rect 29595 10761 29604 10795
rect 29552 10752 29604 10761
rect 30104 10752 30156 10804
rect 31024 10752 31076 10804
rect 31392 10752 31444 10804
rect 30012 10684 30064 10736
rect 28724 10659 28776 10668
rect 28724 10625 28733 10659
rect 28733 10625 28767 10659
rect 28767 10625 28776 10659
rect 28724 10616 28776 10625
rect 28816 10591 28868 10600
rect 28816 10557 28825 10591
rect 28825 10557 28859 10591
rect 28859 10557 28868 10591
rect 28816 10548 28868 10557
rect 28448 10480 28500 10532
rect 29368 10548 29420 10600
rect 32128 10616 32180 10668
rect 40132 10752 40184 10804
rect 35716 10684 35768 10736
rect 36084 10727 36136 10736
rect 36084 10693 36093 10727
rect 36093 10693 36127 10727
rect 36127 10693 36136 10727
rect 36084 10684 36136 10693
rect 30748 10548 30800 10600
rect 30932 10548 30984 10600
rect 31208 10591 31260 10600
rect 31208 10557 31217 10591
rect 31217 10557 31251 10591
rect 31251 10557 31260 10591
rect 31208 10548 31260 10557
rect 30196 10480 30248 10532
rect 31116 10480 31168 10532
rect 32772 10548 32824 10600
rect 28908 10412 28960 10464
rect 31024 10412 31076 10464
rect 33416 10591 33468 10600
rect 33416 10557 33425 10591
rect 33425 10557 33459 10591
rect 33459 10557 33468 10591
rect 33416 10548 33468 10557
rect 34152 10548 34204 10600
rect 40316 10616 40368 10668
rect 42800 10659 42852 10668
rect 42800 10625 42809 10659
rect 42809 10625 42843 10659
rect 42843 10625 42852 10659
rect 42800 10616 42852 10625
rect 45560 10616 45612 10668
rect 34704 10480 34756 10532
rect 35072 10480 35124 10532
rect 37004 10548 37056 10600
rect 40684 10548 40736 10600
rect 49148 10591 49200 10600
rect 49148 10557 49157 10591
rect 49157 10557 49191 10591
rect 49191 10557 49200 10591
rect 49148 10548 49200 10557
rect 38752 10480 38804 10532
rect 34796 10412 34848 10464
rect 36360 10412 36412 10464
rect 37832 10412 37884 10464
rect 44088 10412 44140 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 28724 10208 28776 10260
rect 29828 10140 29880 10192
rect 32404 10251 32456 10260
rect 32404 10217 32413 10251
rect 32413 10217 32447 10251
rect 32447 10217 32456 10251
rect 32404 10208 32456 10217
rect 32680 10208 32732 10260
rect 33324 10208 33376 10260
rect 34152 10208 34204 10260
rect 36636 10208 36688 10260
rect 25320 10072 25372 10124
rect 25780 10115 25832 10124
rect 25780 10081 25789 10115
rect 25789 10081 25823 10115
rect 25823 10081 25832 10115
rect 25780 10072 25832 10081
rect 29460 10072 29512 10124
rect 29736 10072 29788 10124
rect 35348 10140 35400 10192
rect 32312 10072 32364 10124
rect 32772 10072 32824 10124
rect 34888 10004 34940 10056
rect 37004 10072 37056 10124
rect 37188 10004 37240 10056
rect 38660 10004 38712 10056
rect 26608 9936 26660 9988
rect 30932 9979 30984 9988
rect 30932 9945 30941 9979
rect 30941 9945 30975 9979
rect 30975 9945 30984 9979
rect 30932 9936 30984 9945
rect 31392 9936 31444 9988
rect 32220 9936 32272 9988
rect 27528 9911 27580 9920
rect 27528 9877 27537 9911
rect 27537 9877 27571 9911
rect 27571 9877 27580 9911
rect 27528 9868 27580 9877
rect 29552 9868 29604 9920
rect 31024 9868 31076 9920
rect 33232 9911 33284 9920
rect 33232 9877 33241 9911
rect 33241 9877 33275 9911
rect 33275 9877 33284 9911
rect 33232 9868 33284 9877
rect 33324 9911 33376 9920
rect 33324 9877 33333 9911
rect 33333 9877 33367 9911
rect 33367 9877 33376 9911
rect 33324 9868 33376 9877
rect 34612 9936 34664 9988
rect 35072 9936 35124 9988
rect 35716 9936 35768 9988
rect 44640 10004 44692 10056
rect 46940 10004 46992 10056
rect 44180 9936 44232 9988
rect 46296 9979 46348 9988
rect 46296 9945 46305 9979
rect 46305 9945 46339 9979
rect 46339 9945 46348 9979
rect 46296 9936 46348 9945
rect 47032 9979 47084 9988
rect 47032 9945 47041 9979
rect 47041 9945 47075 9979
rect 47075 9945 47084 9979
rect 47032 9936 47084 9945
rect 49148 9979 49200 9988
rect 49148 9945 49157 9979
rect 49157 9945 49191 9979
rect 49191 9945 49200 9979
rect 49148 9936 49200 9945
rect 40408 9868 40460 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 3424 9596 3476 9648
rect 24400 9596 24452 9648
rect 22744 9528 22796 9580
rect 30288 9596 30340 9648
rect 31484 9664 31536 9716
rect 32588 9664 32640 9716
rect 33232 9664 33284 9716
rect 39120 9664 39172 9716
rect 30656 9596 30708 9648
rect 34796 9596 34848 9648
rect 38384 9596 38436 9648
rect 38752 9639 38804 9648
rect 38752 9605 38761 9639
rect 38761 9605 38795 9639
rect 38795 9605 38804 9639
rect 38752 9596 38804 9605
rect 39028 9596 39080 9648
rect 29092 9528 29144 9580
rect 25136 9460 25188 9512
rect 23940 9392 23992 9444
rect 29000 9392 29052 9444
rect 23296 9367 23348 9376
rect 23296 9333 23305 9367
rect 23305 9333 23339 9367
rect 23339 9333 23348 9367
rect 23296 9324 23348 9333
rect 26424 9367 26476 9376
rect 26424 9333 26433 9367
rect 26433 9333 26467 9367
rect 26467 9333 26476 9367
rect 26424 9324 26476 9333
rect 28816 9367 28868 9376
rect 28816 9333 28825 9367
rect 28825 9333 28859 9367
rect 28859 9333 28868 9367
rect 28816 9324 28868 9333
rect 29276 9435 29328 9444
rect 29276 9401 29285 9435
rect 29285 9401 29319 9435
rect 29319 9401 29328 9435
rect 29276 9392 29328 9401
rect 30012 9460 30064 9512
rect 30564 9460 30616 9512
rect 31116 9528 31168 9580
rect 33232 9503 33284 9512
rect 30380 9392 30432 9444
rect 30472 9435 30524 9444
rect 30472 9401 30481 9435
rect 30481 9401 30515 9435
rect 30515 9401 30524 9435
rect 30472 9392 30524 9401
rect 33232 9469 33241 9503
rect 33241 9469 33275 9503
rect 33275 9469 33284 9503
rect 33232 9460 33284 9469
rect 34520 9460 34572 9512
rect 31668 9392 31720 9444
rect 35072 9571 35124 9580
rect 35072 9537 35081 9571
rect 35081 9537 35115 9571
rect 35115 9537 35124 9571
rect 35072 9528 35124 9537
rect 37004 9528 37056 9580
rect 43720 9571 43772 9580
rect 43720 9537 43729 9571
rect 43729 9537 43763 9571
rect 43763 9537 43772 9571
rect 43720 9528 43772 9537
rect 44088 9528 44140 9580
rect 36452 9460 36504 9512
rect 36728 9460 36780 9512
rect 40040 9460 40092 9512
rect 32772 9367 32824 9376
rect 32772 9333 32781 9367
rect 32781 9333 32815 9367
rect 32815 9333 32824 9367
rect 32772 9324 32824 9333
rect 36268 9367 36320 9376
rect 36268 9333 36277 9367
rect 36277 9333 36311 9367
rect 36311 9333 36320 9367
rect 36268 9324 36320 9333
rect 37464 9324 37516 9376
rect 39120 9324 39172 9376
rect 40224 9367 40276 9376
rect 40224 9333 40233 9367
rect 40233 9333 40267 9367
rect 40267 9333 40276 9367
rect 40224 9324 40276 9333
rect 45468 9324 45520 9376
rect 47860 9324 47912 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 22744 9163 22796 9172
rect 22744 9129 22753 9163
rect 22753 9129 22787 9163
rect 22787 9129 22796 9163
rect 22744 9120 22796 9129
rect 34704 9120 34756 9172
rect 35716 9120 35768 9172
rect 27068 9095 27120 9104
rect 27068 9061 27077 9095
rect 27077 9061 27111 9095
rect 27111 9061 27120 9095
rect 27068 9052 27120 9061
rect 24124 8984 24176 9036
rect 27528 8984 27580 9036
rect 28356 9052 28408 9104
rect 31944 9095 31996 9104
rect 31944 9061 31953 9095
rect 31953 9061 31987 9095
rect 31987 9061 31996 9095
rect 31944 9052 31996 9061
rect 37280 9052 37332 9104
rect 29736 9027 29788 9036
rect 29736 8993 29745 9027
rect 29745 8993 29779 9027
rect 29779 8993 29788 9027
rect 29736 8984 29788 8993
rect 31852 8984 31904 9036
rect 32128 8984 32180 9036
rect 32588 9027 32640 9036
rect 32588 8993 32597 9027
rect 32597 8993 32631 9027
rect 32631 8993 32640 9027
rect 32588 8984 32640 8993
rect 32772 8984 32824 9036
rect 45560 9120 45612 9172
rect 46940 9120 46992 9172
rect 40040 9052 40092 9104
rect 2596 8780 2648 8832
rect 24768 8916 24820 8968
rect 28816 8959 28868 8968
rect 28816 8925 28825 8959
rect 28825 8925 28859 8959
rect 28859 8925 28868 8959
rect 28816 8916 28868 8925
rect 31392 8916 31444 8968
rect 34428 8916 34480 8968
rect 34888 8959 34940 8968
rect 34888 8925 34897 8959
rect 34897 8925 34931 8959
rect 34931 8925 34940 8959
rect 34888 8916 34940 8925
rect 36176 8916 36228 8968
rect 37004 8916 37056 8968
rect 23296 8848 23348 8900
rect 26608 8848 26660 8900
rect 23480 8780 23532 8832
rect 35164 8891 35216 8900
rect 35164 8857 35173 8891
rect 35173 8857 35207 8891
rect 35207 8857 35216 8891
rect 35164 8848 35216 8857
rect 31484 8823 31536 8832
rect 31484 8789 31493 8823
rect 31493 8789 31527 8823
rect 31527 8789 31536 8823
rect 31484 8780 31536 8789
rect 32588 8780 32640 8832
rect 33140 8780 33192 8832
rect 33416 8780 33468 8832
rect 38660 8959 38712 8968
rect 38660 8925 38669 8959
rect 38669 8925 38703 8959
rect 38703 8925 38712 8959
rect 38660 8916 38712 8925
rect 38936 8916 38988 8968
rect 40316 8916 40368 8968
rect 37464 8891 37516 8900
rect 37464 8857 37473 8891
rect 37473 8857 37507 8891
rect 37507 8857 37516 8891
rect 37464 8848 37516 8857
rect 38476 8848 38528 8900
rect 39028 8848 39080 8900
rect 37280 8780 37332 8832
rect 44180 8916 44232 8968
rect 45284 8891 45336 8900
rect 45284 8857 45293 8891
rect 45293 8857 45327 8891
rect 45327 8857 45336 8891
rect 45284 8848 45336 8857
rect 49148 8891 49200 8900
rect 49148 8857 49157 8891
rect 49157 8857 49191 8891
rect 49191 8857 49200 8891
rect 49148 8848 49200 8857
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 23480 8619 23532 8628
rect 23480 8585 23489 8619
rect 23489 8585 23523 8619
rect 23523 8585 23532 8619
rect 23480 8576 23532 8585
rect 23940 8619 23992 8628
rect 23940 8585 23949 8619
rect 23949 8585 23983 8619
rect 23983 8585 23992 8619
rect 23940 8576 23992 8585
rect 18512 8508 18564 8560
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 25780 8508 25832 8560
rect 27528 8508 27580 8560
rect 26424 8483 26476 8492
rect 26424 8449 26433 8483
rect 26433 8449 26467 8483
rect 26467 8449 26476 8483
rect 26424 8440 26476 8449
rect 26608 8440 26660 8492
rect 32312 8619 32364 8628
rect 32312 8585 32321 8619
rect 32321 8585 32355 8619
rect 32355 8585 32364 8619
rect 32312 8576 32364 8585
rect 34428 8576 34480 8628
rect 34520 8576 34572 8628
rect 35256 8576 35308 8628
rect 32312 8440 32364 8492
rect 32680 8440 32732 8492
rect 24124 8415 24176 8424
rect 24124 8381 24133 8415
rect 24133 8381 24167 8415
rect 24167 8381 24176 8415
rect 24124 8372 24176 8381
rect 22008 8304 22060 8356
rect 26240 8372 26292 8424
rect 26700 8415 26752 8424
rect 26700 8381 26709 8415
rect 26709 8381 26743 8415
rect 26743 8381 26752 8415
rect 26700 8372 26752 8381
rect 27620 8415 27672 8424
rect 27620 8381 27636 8415
rect 27636 8381 27670 8415
rect 27670 8381 27672 8415
rect 27620 8372 27672 8381
rect 30932 8372 30984 8424
rect 31668 8372 31720 8424
rect 35716 8576 35768 8628
rect 36452 8576 36504 8628
rect 40316 8619 40368 8628
rect 40316 8585 40325 8619
rect 40325 8585 40359 8619
rect 40359 8585 40368 8619
rect 40316 8576 40368 8585
rect 36176 8508 36228 8560
rect 36728 8551 36780 8560
rect 36728 8517 36737 8551
rect 36737 8517 36771 8551
rect 36771 8517 36780 8551
rect 36728 8508 36780 8517
rect 37188 8508 37240 8560
rect 38476 8508 38528 8560
rect 40132 8508 40184 8560
rect 45192 8508 45244 8560
rect 34060 8483 34112 8492
rect 34060 8449 34069 8483
rect 34069 8449 34103 8483
rect 34103 8449 34112 8483
rect 34060 8440 34112 8449
rect 36360 8440 36412 8492
rect 40224 8440 40276 8492
rect 35808 8372 35860 8424
rect 47860 8440 47912 8492
rect 49148 8415 49200 8424
rect 49148 8381 49157 8415
rect 49157 8381 49191 8415
rect 49191 8381 49200 8415
rect 49148 8372 49200 8381
rect 26148 8236 26200 8288
rect 30656 8304 30708 8356
rect 35348 8304 35400 8356
rect 41236 8304 41288 8356
rect 46848 8347 46900 8356
rect 46848 8313 46857 8347
rect 46857 8313 46891 8347
rect 46891 8313 46900 8347
rect 46848 8304 46900 8313
rect 27896 8279 27948 8288
rect 27896 8245 27920 8279
rect 27920 8245 27948 8279
rect 27896 8236 27948 8245
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 27896 8032 27948 8084
rect 29000 8032 29052 8084
rect 32312 8075 32364 8084
rect 32312 8041 32321 8075
rect 32321 8041 32355 8075
rect 32355 8041 32364 8075
rect 32312 8032 32364 8041
rect 35164 8032 35216 8084
rect 44180 8032 44232 8084
rect 30012 7964 30064 8016
rect 31668 7964 31720 8016
rect 34612 7964 34664 8016
rect 45284 7964 45336 8016
rect 25780 7896 25832 7948
rect 27068 7896 27120 7948
rect 28632 7896 28684 7948
rect 31484 7896 31536 7948
rect 32588 7896 32640 7948
rect 37740 7896 37792 7948
rect 28816 7828 28868 7880
rect 31668 7828 31720 7880
rect 32404 7828 32456 7880
rect 35716 7828 35768 7880
rect 35808 7871 35860 7880
rect 35808 7837 35817 7871
rect 35817 7837 35851 7871
rect 35851 7837 35860 7871
rect 35808 7828 35860 7837
rect 37188 7828 37240 7880
rect 26792 7760 26844 7812
rect 23848 7692 23900 7744
rect 35532 7760 35584 7812
rect 33416 7692 33468 7744
rect 40224 7871 40276 7880
rect 40224 7837 40233 7871
rect 40233 7837 40267 7871
rect 40267 7837 40276 7871
rect 40224 7828 40276 7837
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 28540 7420 28592 7472
rect 32496 7463 32548 7472
rect 32496 7429 32505 7463
rect 32505 7429 32539 7463
rect 32539 7429 32548 7463
rect 32496 7420 32548 7429
rect 34888 7488 34940 7540
rect 35808 7488 35860 7540
rect 34704 7420 34756 7472
rect 35256 7420 35308 7472
rect 35716 7463 35768 7472
rect 35716 7429 35725 7463
rect 35725 7429 35759 7463
rect 35759 7429 35768 7463
rect 35716 7420 35768 7429
rect 46296 7420 46348 7472
rect 35532 7352 35584 7404
rect 41236 7352 41288 7404
rect 45468 7352 45520 7404
rect 34152 7284 34204 7336
rect 29276 7216 29328 7268
rect 34612 7284 34664 7336
rect 49148 7327 49200 7336
rect 49148 7293 49157 7327
rect 49157 7293 49191 7327
rect 49191 7293 49200 7327
rect 49148 7284 49200 7293
rect 40224 7216 40276 7268
rect 34428 7148 34480 7200
rect 39028 7148 39080 7200
rect 45468 7148 45520 7200
rect 46940 7191 46992 7200
rect 46940 7157 46949 7191
rect 46949 7157 46983 7191
rect 46983 7157 46992 7191
rect 46940 7148 46992 7157
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 31484 6944 31536 6996
rect 36452 6944 36504 6996
rect 29736 6851 29788 6860
rect 29736 6817 29745 6851
rect 29745 6817 29779 6851
rect 29779 6817 29788 6851
rect 29736 6808 29788 6817
rect 32312 6808 32364 6860
rect 34060 6808 34112 6860
rect 35808 6808 35860 6860
rect 37740 6808 37792 6860
rect 34244 6740 34296 6792
rect 36360 6740 36412 6792
rect 39028 6783 39080 6792
rect 39028 6749 39037 6783
rect 39037 6749 39071 6783
rect 39071 6749 39080 6783
rect 39028 6740 39080 6749
rect 39120 6783 39172 6792
rect 39120 6749 39129 6783
rect 39129 6749 39163 6783
rect 39163 6749 39172 6783
rect 39120 6740 39172 6749
rect 40040 6740 40092 6792
rect 47032 6740 47084 6792
rect 31392 6672 31444 6724
rect 32220 6715 32272 6724
rect 32220 6681 32229 6715
rect 32229 6681 32263 6715
rect 32263 6681 32272 6715
rect 32220 6672 32272 6681
rect 34704 6672 34756 6724
rect 35624 6672 35676 6724
rect 37188 6672 37240 6724
rect 32588 6604 32640 6656
rect 38936 6672 38988 6724
rect 49148 6715 49200 6724
rect 49148 6681 49157 6715
rect 49157 6681 49191 6715
rect 49191 6681 49200 6715
rect 49148 6672 49200 6681
rect 40592 6604 40644 6656
rect 44088 6604 44140 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 31392 6400 31444 6452
rect 32588 6375 32640 6384
rect 32588 6341 32597 6375
rect 32597 6341 32631 6375
rect 32631 6341 32640 6375
rect 32588 6332 32640 6341
rect 34152 6400 34204 6452
rect 34704 6332 34756 6384
rect 37556 6375 37608 6384
rect 37556 6341 37565 6375
rect 37565 6341 37599 6375
rect 37599 6341 37608 6375
rect 37556 6332 37608 6341
rect 38292 6375 38344 6384
rect 38292 6341 38301 6375
rect 38301 6341 38335 6375
rect 38335 6341 38344 6375
rect 38292 6332 38344 6341
rect 39488 6375 39540 6384
rect 39488 6341 39497 6375
rect 39497 6341 39531 6375
rect 39531 6341 39540 6375
rect 39488 6332 39540 6341
rect 32312 6307 32364 6316
rect 32312 6273 32321 6307
rect 32321 6273 32355 6307
rect 32355 6273 32364 6307
rect 32312 6264 32364 6273
rect 37188 6264 37240 6316
rect 40040 6196 40092 6248
rect 45192 6264 45244 6316
rect 48504 6196 48556 6248
rect 49240 6196 49292 6248
rect 39488 6128 39540 6180
rect 42616 6060 42668 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 33416 5856 33468 5908
rect 40224 5856 40276 5908
rect 45192 5899 45244 5908
rect 45192 5865 45201 5899
rect 45201 5865 45235 5899
rect 45235 5865 45244 5899
rect 45192 5856 45244 5865
rect 43352 5788 43404 5840
rect 46848 5788 46900 5840
rect 32220 5720 32272 5772
rect 40132 5720 40184 5772
rect 40408 5720 40460 5772
rect 29184 5652 29236 5704
rect 32404 5695 32456 5704
rect 32404 5661 32413 5695
rect 32413 5661 32447 5695
rect 32447 5661 32456 5695
rect 32404 5652 32456 5661
rect 37372 5652 37424 5704
rect 39212 5652 39264 5704
rect 30012 5584 30064 5636
rect 36820 5584 36872 5636
rect 40592 5652 40644 5704
rect 45468 5652 45520 5704
rect 27528 5516 27580 5568
rect 42800 5584 42852 5636
rect 47032 5627 47084 5636
rect 47032 5593 47041 5627
rect 47041 5593 47075 5627
rect 47075 5593 47084 5627
rect 47032 5584 47084 5593
rect 49148 5627 49200 5636
rect 49148 5593 49157 5627
rect 49157 5593 49191 5627
rect 49191 5593 49200 5627
rect 49148 5584 49200 5593
rect 40500 5516 40552 5568
rect 45468 5516 45520 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 36636 5244 36688 5296
rect 40868 5287 40920 5296
rect 40868 5253 40877 5287
rect 40877 5253 40911 5287
rect 40911 5253 40920 5287
rect 40868 5244 40920 5253
rect 44088 5176 44140 5228
rect 46940 5176 46992 5228
rect 47768 5108 47820 5160
rect 49148 5151 49200 5160
rect 49148 5117 49157 5151
rect 49157 5117 49191 5151
rect 49191 5117 49200 5151
rect 49148 5108 49200 5117
rect 42708 5040 42760 5092
rect 24676 4972 24728 5024
rect 37648 4972 37700 5024
rect 47952 4972 48004 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 10600 4768 10652 4820
rect 26884 4768 26936 4820
rect 31300 4768 31352 4820
rect 46388 4768 46440 4820
rect 13452 4700 13504 4752
rect 24032 4700 24084 4752
rect 47860 4632 47912 4684
rect 11704 4539 11756 4548
rect 11704 4505 11713 4539
rect 11713 4505 11747 4539
rect 11747 4505 11756 4539
rect 11704 4496 11756 4505
rect 13452 4539 13504 4548
rect 13452 4505 13461 4539
rect 13461 4505 13495 4539
rect 13495 4505 13504 4539
rect 13452 4496 13504 4505
rect 24768 4564 24820 4616
rect 46112 4607 46164 4616
rect 46112 4573 46121 4607
rect 46121 4573 46155 4607
rect 46155 4573 46164 4607
rect 46112 4564 46164 4573
rect 47952 4607 48004 4616
rect 47952 4573 47961 4607
rect 47961 4573 47995 4607
rect 47995 4573 48004 4607
rect 47952 4564 48004 4573
rect 26792 4496 26844 4548
rect 48688 4496 48740 4548
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 35348 4088 35400 4140
rect 38936 4088 38988 4140
rect 42800 4088 42852 4140
rect 45468 4088 45520 4140
rect 47032 4088 47084 4140
rect 33876 4020 33928 4072
rect 39028 4020 39080 4072
rect 44180 4020 44232 4072
rect 49148 4063 49200 4072
rect 49148 4029 49157 4063
rect 49157 4029 49191 4063
rect 49191 4029 49200 4063
rect 49148 4020 49200 4029
rect 46296 3927 46348 3936
rect 46296 3893 46305 3927
rect 46305 3893 46339 3927
rect 46339 3893 46348 3927
rect 46296 3884 46348 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 20904 3680 20956 3732
rect 32128 3680 32180 3732
rect 48504 3723 48556 3732
rect 48504 3689 48513 3723
rect 48513 3689 48547 3723
rect 48547 3689 48556 3723
rect 48504 3680 48556 3689
rect 14372 3612 14424 3664
rect 20260 3587 20312 3596
rect 20260 3553 20269 3587
rect 20269 3553 20303 3587
rect 20303 3553 20312 3587
rect 20260 3544 20312 3553
rect 24308 3544 24360 3596
rect 16948 3476 17000 3528
rect 19892 3476 19944 3528
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 3976 3408 4028 3460
rect 23664 3408 23716 3460
rect 28816 3340 28868 3392
rect 33324 3612 33376 3664
rect 29460 3408 29512 3460
rect 30932 3544 30984 3596
rect 34612 3544 34664 3596
rect 36084 3544 36136 3596
rect 39764 3544 39816 3596
rect 41236 3544 41288 3596
rect 44916 3544 44968 3596
rect 30748 3340 30800 3392
rect 34428 3476 34480 3528
rect 38568 3476 38620 3528
rect 40040 3519 40092 3528
rect 40040 3485 40049 3519
rect 40049 3485 40083 3519
rect 40083 3485 40092 3519
rect 40040 3476 40092 3485
rect 40132 3476 40184 3528
rect 42708 3476 42760 3528
rect 47124 3408 47176 3460
rect 35992 3340 36044 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 3976 3179 4028 3188
rect 3976 3145 3985 3179
rect 3985 3145 4019 3179
rect 4019 3145 4028 3179
rect 3976 3136 4028 3145
rect 22008 3136 22060 3188
rect 18604 3068 18656 3120
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 3700 3000 3752 3052
rect 6644 3000 6696 3052
rect 8852 3000 8904 3052
rect 11060 3000 11112 3052
rect 13360 3000 13412 3052
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 22376 3000 22428 3052
rect 33508 3136 33560 3188
rect 2228 2932 2280 2984
rect 12532 2932 12584 2984
rect 14004 2932 14056 2984
rect 17684 2932 17736 2984
rect 19156 2932 19208 2984
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 22100 2932 22152 2984
rect 30564 3068 30616 3120
rect 25320 3043 25372 3052
rect 25320 3009 25329 3043
rect 25329 3009 25363 3043
rect 25363 3009 25372 3043
rect 25320 3000 25372 3009
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 29552 3000 29604 3052
rect 33968 3000 34020 3052
rect 34980 3000 35032 3052
rect 38844 3000 38896 3052
rect 44548 3068 44600 3120
rect 49148 3111 49200 3120
rect 49148 3077 49157 3111
rect 49157 3077 49191 3111
rect 49191 3077 49200 3111
rect 49148 3068 49200 3077
rect 42616 3043 42668 3052
rect 42616 3009 42625 3043
rect 42625 3009 42659 3043
rect 42659 3009 42668 3043
rect 42616 3000 42668 3009
rect 43352 3000 43404 3052
rect 46296 3000 46348 3052
rect 25044 2932 25096 2984
rect 27252 2932 27304 2984
rect 28724 2932 28776 2984
rect 31668 2932 31720 2984
rect 22376 2864 22428 2916
rect 31116 2864 31168 2916
rect 32404 2864 32456 2916
rect 36820 2932 36872 2984
rect 37556 2864 37608 2916
rect 41972 2932 42024 2984
rect 42708 2864 42760 2916
rect 27804 2796 27856 2848
rect 28356 2796 28408 2848
rect 30380 2796 30432 2848
rect 45652 2796 45704 2848
rect 48320 2796 48372 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 11704 2592 11756 2644
rect 30840 2592 30892 2644
rect 19800 2524 19852 2576
rect 10600 2499 10652 2508
rect 10600 2465 10609 2499
rect 10609 2465 10643 2499
rect 10643 2465 10652 2499
rect 10600 2456 10652 2465
rect 13268 2456 13320 2508
rect 1492 2388 1544 2440
rect 2964 2388 3016 2440
rect 7380 2388 7432 2440
rect 4436 2320 4488 2372
rect 5172 2320 5224 2372
rect 5540 2363 5592 2372
rect 5540 2329 5549 2363
rect 5549 2329 5583 2363
rect 5583 2329 5592 2363
rect 5540 2320 5592 2329
rect 5908 2320 5960 2372
rect 8300 2363 8352 2372
rect 8300 2329 8309 2363
rect 8309 2329 8343 2363
rect 8343 2329 8352 2363
rect 8300 2320 8352 2329
rect 9588 2320 9640 2372
rect 9864 2363 9916 2372
rect 9864 2329 9873 2363
rect 9873 2329 9907 2363
rect 9907 2329 9916 2363
rect 9864 2320 9916 2329
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 11796 2388 11848 2440
rect 14740 2388 14792 2440
rect 15476 2388 15528 2440
rect 16488 2388 16540 2440
rect 18420 2456 18472 2508
rect 24584 2524 24636 2576
rect 29000 2524 29052 2576
rect 19984 2388 20036 2440
rect 22836 2388 22888 2440
rect 23572 2388 23624 2440
rect 21180 2320 21232 2372
rect 21364 2320 21416 2372
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 7472 2295 7524 2304
rect 7472 2261 7481 2295
rect 7481 2261 7515 2295
rect 7515 2261 7524 2295
rect 7472 2252 7524 2261
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 16120 2295 16172 2304
rect 16120 2261 16129 2295
rect 16129 2261 16163 2295
rect 16163 2261 16172 2295
rect 16120 2252 16172 2261
rect 17316 2252 17368 2304
rect 22284 2252 22336 2304
rect 24584 2252 24636 2304
rect 25780 2499 25832 2508
rect 25780 2465 25789 2499
rect 25789 2465 25823 2499
rect 25823 2465 25832 2499
rect 25780 2456 25832 2465
rect 26516 2456 26568 2508
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 33600 2524 33652 2576
rect 30380 2499 30432 2508
rect 30380 2465 30389 2499
rect 30389 2465 30423 2499
rect 30423 2465 30432 2499
rect 30380 2456 30432 2465
rect 29276 2388 29328 2440
rect 30196 2388 30248 2440
rect 35348 2456 35400 2508
rect 33784 2388 33836 2440
rect 36268 2388 36320 2440
rect 36360 2388 36412 2440
rect 45376 2592 45428 2644
rect 40224 2524 40276 2576
rect 40592 2456 40644 2508
rect 30656 2320 30708 2372
rect 29368 2252 29420 2304
rect 33140 2252 33192 2304
rect 39488 2320 39540 2372
rect 43444 2456 43496 2508
rect 48320 2499 48372 2508
rect 48320 2465 48329 2499
rect 48329 2465 48363 2499
rect 48363 2465 48372 2499
rect 48320 2456 48372 2465
rect 47768 2431 47820 2440
rect 47768 2397 47777 2431
rect 47777 2397 47811 2431
rect 47811 2397 47820 2431
rect 47768 2388 47820 2397
rect 38292 2252 38344 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
rect 7472 2048 7524 2100
rect 17224 2048 17276 2100
rect 17316 2048 17368 2100
rect 23848 2048 23900 2100
rect 3424 1980 3476 2032
rect 41604 1980 41656 2032
rect 4712 1912 4764 1964
rect 17224 1912 17276 1964
rect 5540 1844 5592 1896
rect 11888 1776 11940 1828
rect 18512 1844 18564 1896
rect 21180 1912 21232 1964
rect 27712 1912 27764 1964
rect 24952 1844 25004 1896
rect 22284 1776 22336 1828
rect 31576 1776 31628 1828
rect 16120 1708 16172 1760
rect 26240 1708 26292 1760
rect 17224 1640 17276 1692
rect 25688 1640 25740 1692
rect 6736 1504 6788 1556
rect 23388 1504 23440 1556
<< metal2 >>
rect 1398 56200 1454 57000
rect 4066 56200 4122 57000
rect 6734 56200 6790 57000
rect 9402 56200 9458 57000
rect 12070 56200 12126 57000
rect 12176 56222 12388 56250
rect 1412 54126 1440 56200
rect 4080 54126 4108 56200
rect 6748 54210 6776 56200
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8392 54256 8444 54262
rect 6748 54182 7052 54210
rect 8392 54198 8444 54204
rect 7024 54126 7052 54182
rect 7104 54188 7156 54194
rect 7104 54130 7156 54136
rect 1400 54120 1452 54126
rect 1400 54062 1452 54068
rect 4068 54120 4120 54126
rect 4068 54062 4120 54068
rect 7012 54120 7064 54126
rect 7012 54062 7064 54068
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 7116 52154 7144 54130
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 8404 53242 8432 54198
rect 9416 54126 9444 56200
rect 12084 56114 12112 56200
rect 12176 56114 12204 56222
rect 12084 56086 12204 56114
rect 9588 54188 9640 54194
rect 9588 54130 9640 54136
rect 12256 54188 12308 54194
rect 12256 54130 12308 54136
rect 9404 54120 9456 54126
rect 9404 54062 9456 54068
rect 8392 53236 8444 53242
rect 8392 53178 8444 53184
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7104 52148 7156 52154
rect 7104 52090 7156 52096
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 9600 51270 9628 54130
rect 12268 51542 12296 54130
rect 12360 54126 12388 56222
rect 14738 56200 14794 57000
rect 17406 56200 17462 57000
rect 17512 56222 17908 56250
rect 14752 54126 14780 56200
rect 17420 56114 17448 56200
rect 17512 56114 17540 56222
rect 17420 56086 17540 56114
rect 15016 54188 15068 54194
rect 15016 54130 15068 54136
rect 17684 54188 17736 54194
rect 17684 54130 17736 54136
rect 12348 54120 12400 54126
rect 12348 54062 12400 54068
rect 14740 54120 14792 54126
rect 14740 54062 14792 54068
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 13728 53100 13780 53106
rect 13728 53042 13780 53048
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12256 51536 12308 51542
rect 12256 51478 12308 51484
rect 9588 51264 9640 51270
rect 9588 51206 9640 51212
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 13740 50454 13768 53042
rect 15028 51610 15056 54130
rect 15200 54052 15252 54058
rect 15200 53994 15252 54000
rect 15016 51604 15068 51610
rect 15016 51546 15068 51552
rect 15212 50522 15240 53994
rect 17500 51400 17552 51406
rect 17500 51342 17552 51348
rect 15200 50516 15252 50522
rect 15200 50458 15252 50464
rect 16120 50516 16172 50522
rect 16120 50458 16172 50464
rect 13728 50448 13780 50454
rect 13728 50390 13780 50396
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 16132 48278 16160 50458
rect 17316 50448 17368 50454
rect 17316 50390 17368 50396
rect 16120 48272 16172 48278
rect 16120 48214 16172 48220
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 17328 47598 17356 50390
rect 17316 47592 17368 47598
rect 17316 47534 17368 47540
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 17328 46034 17356 47534
rect 17512 46170 17540 51342
rect 17696 50522 17724 54130
rect 17880 54126 17908 56222
rect 20074 56200 20130 57000
rect 22742 56200 22798 57000
rect 25410 56200 25466 57000
rect 28078 56200 28134 57000
rect 28184 56222 28396 56250
rect 20088 55214 20116 56200
rect 20088 55186 20208 55214
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 20180 54126 20208 55186
rect 20260 54188 20312 54194
rect 20260 54130 20312 54136
rect 17868 54120 17920 54126
rect 17868 54062 17920 54068
rect 20168 54120 20220 54126
rect 20168 54062 20220 54068
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 19800 52012 19852 52018
rect 19800 51954 19852 51960
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17684 50516 17736 50522
rect 17684 50458 17736 50464
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 19432 48204 19484 48210
rect 19432 48146 19484 48152
rect 18328 48068 18380 48074
rect 18328 48010 18380 48016
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17500 46164 17552 46170
rect 17500 46106 17552 46112
rect 17316 46028 17368 46034
rect 17316 45970 17368 45976
rect 17132 45960 17184 45966
rect 17132 45902 17184 45908
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 17144 37126 17172 45902
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 18340 44742 18368 48010
rect 19444 44878 19472 48146
rect 19524 48000 19576 48006
rect 19524 47942 19576 47948
rect 19536 47598 19564 47942
rect 19812 47802 19840 51954
rect 20272 49434 20300 54130
rect 22756 54126 22784 56200
rect 25424 54194 25452 56200
rect 28092 56114 28120 56200
rect 28184 56114 28212 56222
rect 28092 56086 28212 56114
rect 27950 54428 28258 54437
rect 27950 54426 27956 54428
rect 28012 54426 28036 54428
rect 28092 54426 28116 54428
rect 28172 54426 28196 54428
rect 28252 54426 28258 54428
rect 28012 54374 28014 54426
rect 28194 54374 28196 54426
rect 27950 54372 27956 54374
rect 28012 54372 28036 54374
rect 28092 54372 28116 54374
rect 28172 54372 28196 54374
rect 28252 54372 28258 54374
rect 27950 54363 28258 54372
rect 28368 54194 28396 56222
rect 30746 56200 30802 57000
rect 33414 56200 33470 57000
rect 36082 56200 36138 57000
rect 38750 56200 38806 57000
rect 41418 56200 41474 57000
rect 44086 56200 44142 57000
rect 46754 56200 46810 57000
rect 48410 56264 48466 56273
rect 29552 54324 29604 54330
rect 29552 54266 29604 54272
rect 22836 54188 22888 54194
rect 22836 54130 22888 54136
rect 25412 54188 25464 54194
rect 25412 54130 25464 54136
rect 28356 54188 28408 54194
rect 28356 54130 28408 54136
rect 22744 54120 22796 54126
rect 22744 54062 22796 54068
rect 20536 53984 20588 53990
rect 20536 53926 20588 53932
rect 20548 50318 20576 53926
rect 21640 51468 21692 51474
rect 21640 51410 21692 51416
rect 20536 50312 20588 50318
rect 20536 50254 20588 50260
rect 20260 49428 20312 49434
rect 20260 49370 20312 49376
rect 19800 47796 19852 47802
rect 19800 47738 19852 47744
rect 19524 47592 19576 47598
rect 19524 47534 19576 47540
rect 19812 47054 19840 47738
rect 20548 47734 20576 50254
rect 20628 50244 20680 50250
rect 20628 50186 20680 50192
rect 20536 47728 20588 47734
rect 20536 47670 20588 47676
rect 19800 47048 19852 47054
rect 19800 46990 19852 46996
rect 19432 44872 19484 44878
rect 19432 44814 19484 44820
rect 18328 44736 18380 44742
rect 18328 44678 18380 44684
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 19444 41682 19472 44814
rect 19812 44402 19840 46990
rect 20548 46714 20576 47670
rect 20536 46708 20588 46714
rect 20536 46650 20588 46656
rect 20548 45966 20576 46650
rect 20536 45960 20588 45966
rect 20536 45902 20588 45908
rect 20640 44538 20668 50186
rect 21456 49156 21508 49162
rect 21456 49098 21508 49104
rect 21180 47592 21232 47598
rect 21180 47534 21232 47540
rect 20996 46096 21048 46102
rect 20996 46038 21048 46044
rect 20628 44532 20680 44538
rect 20628 44474 20680 44480
rect 19800 44396 19852 44402
rect 19800 44338 19852 44344
rect 19984 44328 20036 44334
rect 19984 44270 20036 44276
rect 19432 41676 19484 41682
rect 19432 41618 19484 41624
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17132 37120 17184 37126
rect 17132 37062 17184 37068
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 19996 34202 20024 44270
rect 21008 42226 21036 46038
rect 21192 45082 21220 47534
rect 21180 45076 21232 45082
rect 21180 45018 21232 45024
rect 21468 42362 21496 49098
rect 21652 46170 21680 51410
rect 22744 51332 22796 51338
rect 22744 51274 22796 51280
rect 22008 47456 22060 47462
rect 22008 47398 22060 47404
rect 22020 46510 22048 47398
rect 22468 46708 22520 46714
rect 22468 46650 22520 46656
rect 22008 46504 22060 46510
rect 22008 46446 22060 46452
rect 21548 46164 21600 46170
rect 21548 46106 21600 46112
rect 21640 46164 21692 46170
rect 21640 46106 21692 46112
rect 21560 44946 21588 46106
rect 21548 44940 21600 44946
rect 21548 44882 21600 44888
rect 21456 42356 21508 42362
rect 21456 42298 21508 42304
rect 20996 42220 21048 42226
rect 20996 42162 21048 42168
rect 20812 42152 20864 42158
rect 20812 42094 20864 42100
rect 19984 34196 20036 34202
rect 19984 34138 20036 34144
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 20824 30938 20852 42094
rect 21560 41818 21588 44882
rect 22480 44402 22508 46650
rect 22756 45554 22784 51274
rect 22848 49434 22876 54130
rect 24400 53984 24452 53990
rect 24400 53926 24452 53932
rect 25688 53984 25740 53990
rect 25688 53926 25740 53932
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22836 49428 22888 49434
rect 22836 49370 22888 49376
rect 23296 49156 23348 49162
rect 23296 49098 23348 49104
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22756 45526 22876 45554
rect 22848 45490 22876 45526
rect 22836 45484 22888 45490
rect 22836 45426 22888 45432
rect 22848 44538 22876 45426
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22836 44532 22888 44538
rect 22836 44474 22888 44480
rect 22468 44396 22520 44402
rect 22468 44338 22520 44344
rect 22560 44192 22612 44198
rect 22560 44134 22612 44140
rect 21548 41812 21600 41818
rect 21548 41754 21600 41760
rect 22572 41478 22600 44134
rect 22652 42220 22704 42226
rect 22652 42162 22704 42168
rect 22560 41472 22612 41478
rect 22560 41414 22612 41420
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 20812 30932 20864 30938
rect 20812 30874 20864 30880
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 22480 18970 22508 30670
rect 22572 28218 22600 37198
rect 22664 30938 22692 42162
rect 22848 42158 22876 44474
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 23308 42362 23336 49098
rect 24412 46646 24440 53926
rect 25700 47122 25728 53926
rect 27950 53340 28258 53349
rect 27950 53338 27956 53340
rect 28012 53338 28036 53340
rect 28092 53338 28116 53340
rect 28172 53338 28196 53340
rect 28252 53338 28258 53340
rect 28012 53286 28014 53338
rect 28194 53286 28196 53338
rect 27950 53284 27956 53286
rect 28012 53284 28036 53286
rect 28092 53284 28116 53286
rect 28172 53284 28196 53286
rect 28252 53284 28258 53286
rect 27950 53275 28258 53284
rect 27950 52252 28258 52261
rect 27950 52250 27956 52252
rect 28012 52250 28036 52252
rect 28092 52250 28116 52252
rect 28172 52250 28196 52252
rect 28252 52250 28258 52252
rect 28012 52198 28014 52250
rect 28194 52198 28196 52250
rect 27950 52196 27956 52198
rect 28012 52196 28036 52198
rect 28092 52196 28116 52198
rect 28172 52196 28196 52198
rect 28252 52196 28258 52198
rect 27950 52187 28258 52196
rect 27950 51164 28258 51173
rect 27950 51162 27956 51164
rect 28012 51162 28036 51164
rect 28092 51162 28116 51164
rect 28172 51162 28196 51164
rect 28252 51162 28258 51164
rect 28012 51110 28014 51162
rect 28194 51110 28196 51162
rect 27950 51108 27956 51110
rect 28012 51108 28036 51110
rect 28092 51108 28116 51110
rect 28172 51108 28196 51110
rect 28252 51108 28258 51110
rect 27950 51099 28258 51108
rect 27950 50076 28258 50085
rect 27950 50074 27956 50076
rect 28012 50074 28036 50076
rect 28092 50074 28116 50076
rect 28172 50074 28196 50076
rect 28252 50074 28258 50076
rect 28012 50022 28014 50074
rect 28194 50022 28196 50074
rect 27950 50020 27956 50022
rect 28012 50020 28036 50022
rect 28092 50020 28116 50022
rect 28172 50020 28196 50022
rect 28252 50020 28258 50022
rect 27950 50011 28258 50020
rect 27950 48988 28258 48997
rect 27950 48986 27956 48988
rect 28012 48986 28036 48988
rect 28092 48986 28116 48988
rect 28172 48986 28196 48988
rect 28252 48986 28258 48988
rect 28012 48934 28014 48986
rect 28194 48934 28196 48986
rect 27950 48932 27956 48934
rect 28012 48932 28036 48934
rect 28092 48932 28116 48934
rect 28172 48932 28196 48934
rect 28252 48932 28258 48934
rect 27950 48923 28258 48932
rect 27950 47900 28258 47909
rect 27950 47898 27956 47900
rect 28012 47898 28036 47900
rect 28092 47898 28116 47900
rect 28172 47898 28196 47900
rect 28252 47898 28258 47900
rect 28012 47846 28014 47898
rect 28194 47846 28196 47898
rect 27950 47844 27956 47846
rect 28012 47844 28036 47846
rect 28092 47844 28116 47846
rect 28172 47844 28196 47846
rect 28252 47844 28258 47846
rect 27950 47835 28258 47844
rect 25688 47116 25740 47122
rect 25688 47058 25740 47064
rect 27528 46980 27580 46986
rect 27528 46922 27580 46928
rect 24400 46640 24452 46646
rect 24400 46582 24452 46588
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 23388 44804 23440 44810
rect 23388 44746 23440 44752
rect 23296 42356 23348 42362
rect 23296 42298 23348 42304
rect 22836 42152 22888 42158
rect 22836 42094 22888 42100
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 23400 41682 23428 44746
rect 22836 41676 22888 41682
rect 22836 41618 22888 41624
rect 23388 41676 23440 41682
rect 23388 41618 23440 41624
rect 22848 34542 22876 41618
rect 24308 41608 24360 41614
rect 24308 41550 24360 41556
rect 23388 41540 23440 41546
rect 23388 41482 23440 41488
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23400 34746 23428 41482
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 24320 34610 24348 41550
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 22836 34536 22888 34542
rect 22836 34478 22888 34484
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 22560 28212 22612 28218
rect 22560 28154 22612 28160
rect 22756 26234 22784 33934
rect 22848 29646 22876 34478
rect 24216 34400 24268 34406
rect 24216 34342 24268 34348
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22756 26206 22876 26234
rect 22848 24410 22876 26206
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22836 24404 22888 24410
rect 22836 24346 22888 24352
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23400 19514 23428 30670
rect 24228 28014 24256 34342
rect 24216 28008 24268 28014
rect 24216 27950 24268 27956
rect 24228 27334 24256 27950
rect 24320 27402 24348 34546
rect 24780 31890 24808 46446
rect 27540 33862 27568 46922
rect 27950 46812 28258 46821
rect 27950 46810 27956 46812
rect 28012 46810 28036 46812
rect 28092 46810 28116 46812
rect 28172 46810 28196 46812
rect 28252 46810 28258 46812
rect 28012 46758 28014 46810
rect 28194 46758 28196 46810
rect 27950 46756 27956 46758
rect 28012 46756 28036 46758
rect 28092 46756 28116 46758
rect 28172 46756 28196 46758
rect 28252 46756 28258 46758
rect 27950 46747 28258 46756
rect 28908 46028 28960 46034
rect 28908 45970 28960 45976
rect 27950 45724 28258 45733
rect 27950 45722 27956 45724
rect 28012 45722 28036 45724
rect 28092 45722 28116 45724
rect 28172 45722 28196 45724
rect 28252 45722 28258 45724
rect 28012 45670 28014 45722
rect 28194 45670 28196 45722
rect 27950 45668 27956 45670
rect 28012 45668 28036 45670
rect 28092 45668 28116 45670
rect 28172 45668 28196 45670
rect 28252 45668 28258 45670
rect 27950 45659 28258 45668
rect 27950 44636 28258 44645
rect 27950 44634 27956 44636
rect 28012 44634 28036 44636
rect 28092 44634 28116 44636
rect 28172 44634 28196 44636
rect 28252 44634 28258 44636
rect 28012 44582 28014 44634
rect 28194 44582 28196 44634
rect 27950 44580 27956 44582
rect 28012 44580 28036 44582
rect 28092 44580 28116 44582
rect 28172 44580 28196 44582
rect 28252 44580 28258 44582
rect 27950 44571 28258 44580
rect 27950 43548 28258 43557
rect 27950 43546 27956 43548
rect 28012 43546 28036 43548
rect 28092 43546 28116 43548
rect 28172 43546 28196 43548
rect 28252 43546 28258 43548
rect 28012 43494 28014 43546
rect 28194 43494 28196 43546
rect 27950 43492 27956 43494
rect 28012 43492 28036 43494
rect 28092 43492 28116 43494
rect 28172 43492 28196 43494
rect 28252 43492 28258 43494
rect 27950 43483 28258 43492
rect 27950 42460 28258 42469
rect 27950 42458 27956 42460
rect 28012 42458 28036 42460
rect 28092 42458 28116 42460
rect 28172 42458 28196 42460
rect 28252 42458 28258 42460
rect 28012 42406 28014 42458
rect 28194 42406 28196 42458
rect 27950 42404 27956 42406
rect 28012 42404 28036 42406
rect 28092 42404 28116 42406
rect 28172 42404 28196 42406
rect 28252 42404 28258 42406
rect 27950 42395 28258 42404
rect 27950 41372 28258 41381
rect 27950 41370 27956 41372
rect 28012 41370 28036 41372
rect 28092 41370 28116 41372
rect 28172 41370 28196 41372
rect 28252 41370 28258 41372
rect 28012 41318 28014 41370
rect 28194 41318 28196 41370
rect 27950 41316 27956 41318
rect 28012 41316 28036 41318
rect 28092 41316 28116 41318
rect 28172 41316 28196 41318
rect 28252 41316 28258 41318
rect 27950 41307 28258 41316
rect 27950 40284 28258 40293
rect 27950 40282 27956 40284
rect 28012 40282 28036 40284
rect 28092 40282 28116 40284
rect 28172 40282 28196 40284
rect 28252 40282 28258 40284
rect 28012 40230 28014 40282
rect 28194 40230 28196 40282
rect 27950 40228 27956 40230
rect 28012 40228 28036 40230
rect 28092 40228 28116 40230
rect 28172 40228 28196 40230
rect 28252 40228 28258 40230
rect 27950 40219 28258 40228
rect 27950 39196 28258 39205
rect 27950 39194 27956 39196
rect 28012 39194 28036 39196
rect 28092 39194 28116 39196
rect 28172 39194 28196 39196
rect 28252 39194 28258 39196
rect 28012 39142 28014 39194
rect 28194 39142 28196 39194
rect 27950 39140 27956 39142
rect 28012 39140 28036 39142
rect 28092 39140 28116 39142
rect 28172 39140 28196 39142
rect 28252 39140 28258 39142
rect 27950 39131 28258 39140
rect 27950 38108 28258 38117
rect 27950 38106 27956 38108
rect 28012 38106 28036 38108
rect 28092 38106 28116 38108
rect 28172 38106 28196 38108
rect 28252 38106 28258 38108
rect 28012 38054 28014 38106
rect 28194 38054 28196 38106
rect 27950 38052 27956 38054
rect 28012 38052 28036 38054
rect 28092 38052 28116 38054
rect 28172 38052 28196 38054
rect 28252 38052 28258 38054
rect 27950 38043 28258 38052
rect 27950 37020 28258 37029
rect 27950 37018 27956 37020
rect 28012 37018 28036 37020
rect 28092 37018 28116 37020
rect 28172 37018 28196 37020
rect 28252 37018 28258 37020
rect 28012 36966 28014 37018
rect 28194 36966 28196 37018
rect 27950 36964 27956 36966
rect 28012 36964 28036 36966
rect 28092 36964 28116 36966
rect 28172 36964 28196 36966
rect 28252 36964 28258 36966
rect 27950 36955 28258 36964
rect 27950 35932 28258 35941
rect 27950 35930 27956 35932
rect 28012 35930 28036 35932
rect 28092 35930 28116 35932
rect 28172 35930 28196 35932
rect 28252 35930 28258 35932
rect 28012 35878 28014 35930
rect 28194 35878 28196 35930
rect 27950 35876 27956 35878
rect 28012 35876 28036 35878
rect 28092 35876 28116 35878
rect 28172 35876 28196 35878
rect 28252 35876 28258 35878
rect 27950 35867 28258 35876
rect 27950 34844 28258 34853
rect 27950 34842 27956 34844
rect 28012 34842 28036 34844
rect 28092 34842 28116 34844
rect 28172 34842 28196 34844
rect 28252 34842 28258 34844
rect 28012 34790 28014 34842
rect 28194 34790 28196 34842
rect 27950 34788 27956 34790
rect 28012 34788 28036 34790
rect 28092 34788 28116 34790
rect 28172 34788 28196 34790
rect 28252 34788 28258 34790
rect 27950 34779 28258 34788
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27540 33697 27568 33798
rect 27950 33756 28258 33765
rect 27950 33754 27956 33756
rect 28012 33754 28036 33756
rect 28092 33754 28116 33756
rect 28172 33754 28196 33756
rect 28252 33754 28258 33756
rect 28012 33702 28014 33754
rect 28194 33702 28196 33754
rect 27950 33700 27956 33702
rect 28012 33700 28036 33702
rect 28092 33700 28116 33702
rect 28172 33700 28196 33702
rect 28252 33700 28258 33702
rect 27526 33688 27582 33697
rect 27950 33691 28258 33700
rect 27526 33623 27582 33632
rect 28920 33289 28948 45970
rect 29564 45490 29592 54266
rect 30760 54194 30788 56200
rect 33428 54194 33456 56200
rect 36096 54262 36124 56200
rect 37950 54428 38258 54437
rect 37950 54426 37956 54428
rect 38012 54426 38036 54428
rect 38092 54426 38116 54428
rect 38172 54426 38196 54428
rect 38252 54426 38258 54428
rect 38012 54374 38014 54426
rect 38194 54374 38196 54426
rect 37950 54372 37956 54374
rect 38012 54372 38036 54374
rect 38092 54372 38116 54374
rect 38172 54372 38196 54374
rect 38252 54372 38258 54374
rect 37950 54363 38258 54372
rect 36084 54256 36136 54262
rect 36084 54198 36136 54204
rect 38764 54194 38792 56200
rect 41432 54194 41460 56200
rect 44100 54194 44128 56200
rect 46768 54262 46796 56200
rect 48410 56199 48466 56208
rect 49422 56200 49478 57000
rect 48226 55448 48282 55457
rect 48226 55383 48282 55392
rect 48240 54618 48268 55383
rect 48240 54590 48360 54618
rect 47950 54428 48258 54437
rect 47950 54426 47956 54428
rect 48012 54426 48036 54428
rect 48092 54426 48116 54428
rect 48172 54426 48196 54428
rect 48252 54426 48258 54428
rect 48012 54374 48014 54426
rect 48194 54374 48196 54426
rect 47950 54372 47956 54374
rect 48012 54372 48036 54374
rect 48092 54372 48116 54374
rect 48172 54372 48196 54374
rect 48252 54372 48258 54374
rect 47950 54363 48258 54372
rect 46756 54256 46808 54262
rect 46756 54198 46808 54204
rect 48332 54194 48360 54590
rect 30748 54188 30800 54194
rect 30748 54130 30800 54136
rect 33416 54188 33468 54194
rect 33416 54130 33468 54136
rect 38752 54188 38804 54194
rect 38752 54130 38804 54136
rect 41420 54188 41472 54194
rect 41420 54130 41472 54136
rect 44088 54188 44140 54194
rect 44088 54130 44140 54136
rect 48320 54188 48372 54194
rect 48320 54130 48372 54136
rect 30840 53984 30892 53990
rect 30840 53926 30892 53932
rect 39028 53984 39080 53990
rect 39028 53926 39080 53932
rect 41696 53984 41748 53990
rect 41696 53926 41748 53932
rect 44364 53984 44416 53990
rect 44364 53926 44416 53932
rect 46940 53984 46992 53990
rect 46940 53926 46992 53932
rect 30852 46102 30880 53926
rect 32950 53884 33258 53893
rect 32950 53882 32956 53884
rect 33012 53882 33036 53884
rect 33092 53882 33116 53884
rect 33172 53882 33196 53884
rect 33252 53882 33258 53884
rect 33012 53830 33014 53882
rect 33194 53830 33196 53882
rect 32950 53828 32956 53830
rect 33012 53828 33036 53830
rect 33092 53828 33116 53830
rect 33172 53828 33196 53830
rect 33252 53828 33258 53830
rect 32950 53819 33258 53828
rect 37950 53340 38258 53349
rect 37950 53338 37956 53340
rect 38012 53338 38036 53340
rect 38092 53338 38116 53340
rect 38172 53338 38196 53340
rect 38252 53338 38258 53340
rect 38012 53286 38014 53338
rect 38194 53286 38196 53338
rect 37950 53284 37956 53286
rect 38012 53284 38036 53286
rect 38092 53284 38116 53286
rect 38172 53284 38196 53286
rect 38252 53284 38258 53286
rect 37950 53275 38258 53284
rect 34704 52896 34756 52902
rect 34704 52838 34756 52844
rect 32950 52796 33258 52805
rect 32950 52794 32956 52796
rect 33012 52794 33036 52796
rect 33092 52794 33116 52796
rect 33172 52794 33196 52796
rect 33252 52794 33258 52796
rect 33012 52742 33014 52794
rect 33194 52742 33196 52794
rect 32950 52740 32956 52742
rect 33012 52740 33036 52742
rect 33092 52740 33116 52742
rect 33172 52740 33196 52742
rect 33252 52740 33258 52742
rect 32950 52731 33258 52740
rect 32950 51708 33258 51717
rect 32950 51706 32956 51708
rect 33012 51706 33036 51708
rect 33092 51706 33116 51708
rect 33172 51706 33196 51708
rect 33252 51706 33258 51708
rect 33012 51654 33014 51706
rect 33194 51654 33196 51706
rect 32950 51652 32956 51654
rect 33012 51652 33036 51654
rect 33092 51652 33116 51654
rect 33172 51652 33196 51654
rect 33252 51652 33258 51654
rect 32950 51643 33258 51652
rect 32950 50620 33258 50629
rect 32950 50618 32956 50620
rect 33012 50618 33036 50620
rect 33092 50618 33116 50620
rect 33172 50618 33196 50620
rect 33252 50618 33258 50620
rect 33012 50566 33014 50618
rect 33194 50566 33196 50618
rect 32950 50564 32956 50566
rect 33012 50564 33036 50566
rect 33092 50564 33116 50566
rect 33172 50564 33196 50566
rect 33252 50564 33258 50566
rect 32950 50555 33258 50564
rect 32950 49532 33258 49541
rect 32950 49530 32956 49532
rect 33012 49530 33036 49532
rect 33092 49530 33116 49532
rect 33172 49530 33196 49532
rect 33252 49530 33258 49532
rect 33012 49478 33014 49530
rect 33194 49478 33196 49530
rect 32950 49476 32956 49478
rect 33012 49476 33036 49478
rect 33092 49476 33116 49478
rect 33172 49476 33196 49478
rect 33252 49476 33258 49478
rect 32950 49467 33258 49476
rect 32950 48444 33258 48453
rect 32950 48442 32956 48444
rect 33012 48442 33036 48444
rect 33092 48442 33116 48444
rect 33172 48442 33196 48444
rect 33252 48442 33258 48444
rect 33012 48390 33014 48442
rect 33194 48390 33196 48442
rect 32950 48388 32956 48390
rect 33012 48388 33036 48390
rect 33092 48388 33116 48390
rect 33172 48388 33196 48390
rect 33252 48388 33258 48390
rect 32950 48379 33258 48388
rect 33692 48000 33744 48006
rect 33692 47942 33744 47948
rect 32950 47356 33258 47365
rect 32950 47354 32956 47356
rect 33012 47354 33036 47356
rect 33092 47354 33116 47356
rect 33172 47354 33196 47356
rect 33252 47354 33258 47356
rect 33012 47302 33014 47354
rect 33194 47302 33196 47354
rect 32950 47300 32956 47302
rect 33012 47300 33036 47302
rect 33092 47300 33116 47302
rect 33172 47300 33196 47302
rect 33252 47300 33258 47302
rect 32950 47291 33258 47300
rect 32950 46268 33258 46277
rect 32950 46266 32956 46268
rect 33012 46266 33036 46268
rect 33092 46266 33116 46268
rect 33172 46266 33196 46268
rect 33252 46266 33258 46268
rect 33012 46214 33014 46266
rect 33194 46214 33196 46266
rect 32950 46212 32956 46214
rect 33012 46212 33036 46214
rect 33092 46212 33116 46214
rect 33172 46212 33196 46214
rect 33252 46212 33258 46214
rect 32950 46203 33258 46212
rect 30840 46096 30892 46102
rect 30840 46038 30892 46044
rect 29552 45484 29604 45490
rect 29552 45426 29604 45432
rect 31392 45416 31444 45422
rect 31392 45358 31444 45364
rect 31404 33386 31432 45358
rect 32950 45180 33258 45189
rect 32950 45178 32956 45180
rect 33012 45178 33036 45180
rect 33092 45178 33116 45180
rect 33172 45178 33196 45180
rect 33252 45178 33258 45180
rect 33012 45126 33014 45178
rect 33194 45126 33196 45178
rect 32950 45124 32956 45126
rect 33012 45124 33036 45126
rect 33092 45124 33116 45126
rect 33172 45124 33196 45126
rect 33252 45124 33258 45126
rect 32950 45115 33258 45124
rect 32950 44092 33258 44101
rect 32950 44090 32956 44092
rect 33012 44090 33036 44092
rect 33092 44090 33116 44092
rect 33172 44090 33196 44092
rect 33252 44090 33258 44092
rect 33012 44038 33014 44090
rect 33194 44038 33196 44090
rect 32950 44036 32956 44038
rect 33012 44036 33036 44038
rect 33092 44036 33116 44038
rect 33172 44036 33196 44038
rect 33252 44036 33258 44038
rect 32950 44027 33258 44036
rect 32950 43004 33258 43013
rect 32950 43002 32956 43004
rect 33012 43002 33036 43004
rect 33092 43002 33116 43004
rect 33172 43002 33196 43004
rect 33252 43002 33258 43004
rect 33012 42950 33014 43002
rect 33194 42950 33196 43002
rect 32950 42948 32956 42950
rect 33012 42948 33036 42950
rect 33092 42948 33116 42950
rect 33172 42948 33196 42950
rect 33252 42948 33258 42950
rect 32950 42939 33258 42948
rect 32950 41916 33258 41925
rect 32950 41914 32956 41916
rect 33012 41914 33036 41916
rect 33092 41914 33116 41916
rect 33172 41914 33196 41916
rect 33252 41914 33258 41916
rect 33012 41862 33014 41914
rect 33194 41862 33196 41914
rect 32950 41860 32956 41862
rect 33012 41860 33036 41862
rect 33092 41860 33116 41862
rect 33172 41860 33196 41862
rect 33252 41860 33258 41862
rect 32950 41851 33258 41860
rect 32950 40828 33258 40837
rect 32950 40826 32956 40828
rect 33012 40826 33036 40828
rect 33092 40826 33116 40828
rect 33172 40826 33196 40828
rect 33252 40826 33258 40828
rect 33012 40774 33014 40826
rect 33194 40774 33196 40826
rect 32950 40772 32956 40774
rect 33012 40772 33036 40774
rect 33092 40772 33116 40774
rect 33172 40772 33196 40774
rect 33252 40772 33258 40774
rect 32950 40763 33258 40772
rect 32950 39740 33258 39749
rect 32950 39738 32956 39740
rect 33012 39738 33036 39740
rect 33092 39738 33116 39740
rect 33172 39738 33196 39740
rect 33252 39738 33258 39740
rect 33012 39686 33014 39738
rect 33194 39686 33196 39738
rect 32950 39684 32956 39686
rect 33012 39684 33036 39686
rect 33092 39684 33116 39686
rect 33172 39684 33196 39686
rect 33252 39684 33258 39686
rect 32950 39675 33258 39684
rect 32950 38652 33258 38661
rect 32950 38650 32956 38652
rect 33012 38650 33036 38652
rect 33092 38650 33116 38652
rect 33172 38650 33196 38652
rect 33252 38650 33258 38652
rect 33012 38598 33014 38650
rect 33194 38598 33196 38650
rect 32950 38596 32956 38598
rect 33012 38596 33036 38598
rect 33092 38596 33116 38598
rect 33172 38596 33196 38598
rect 33252 38596 33258 38598
rect 32950 38587 33258 38596
rect 32950 37564 33258 37573
rect 32950 37562 32956 37564
rect 33012 37562 33036 37564
rect 33092 37562 33116 37564
rect 33172 37562 33196 37564
rect 33252 37562 33258 37564
rect 33012 37510 33014 37562
rect 33194 37510 33196 37562
rect 32950 37508 32956 37510
rect 33012 37508 33036 37510
rect 33092 37508 33116 37510
rect 33172 37508 33196 37510
rect 33252 37508 33258 37510
rect 32950 37499 33258 37508
rect 32950 36476 33258 36485
rect 32950 36474 32956 36476
rect 33012 36474 33036 36476
rect 33092 36474 33116 36476
rect 33172 36474 33196 36476
rect 33252 36474 33258 36476
rect 33012 36422 33014 36474
rect 33194 36422 33196 36474
rect 32950 36420 32956 36422
rect 33012 36420 33036 36422
rect 33092 36420 33116 36422
rect 33172 36420 33196 36422
rect 33252 36420 33258 36422
rect 32950 36411 33258 36420
rect 33704 35894 33732 47942
rect 33704 35866 34100 35894
rect 32950 35388 33258 35397
rect 32950 35386 32956 35388
rect 33012 35386 33036 35388
rect 33092 35386 33116 35388
rect 33172 35386 33196 35388
rect 33252 35386 33258 35388
rect 33012 35334 33014 35386
rect 33194 35334 33196 35386
rect 32950 35332 32956 35334
rect 33012 35332 33036 35334
rect 33092 35332 33116 35334
rect 33172 35332 33196 35334
rect 33252 35332 33258 35334
rect 32950 35323 33258 35332
rect 32950 34300 33258 34309
rect 32950 34298 32956 34300
rect 33012 34298 33036 34300
rect 33092 34298 33116 34300
rect 33172 34298 33196 34300
rect 33252 34298 33258 34300
rect 33012 34246 33014 34298
rect 33194 34246 33196 34298
rect 32950 34244 32956 34246
rect 33012 34244 33036 34246
rect 33092 34244 33116 34246
rect 33172 34244 33196 34246
rect 33252 34244 33258 34246
rect 32950 34235 33258 34244
rect 31392 33380 31444 33386
rect 31392 33322 31444 33328
rect 28906 33280 28962 33289
rect 28906 33215 28962 33224
rect 32950 33212 33258 33221
rect 32950 33210 32956 33212
rect 33012 33210 33036 33212
rect 33092 33210 33116 33212
rect 33172 33210 33196 33212
rect 33252 33210 33258 33212
rect 33012 33158 33014 33210
rect 33194 33158 33196 33210
rect 32950 33156 32956 33158
rect 33012 33156 33036 33158
rect 33092 33156 33116 33158
rect 33172 33156 33196 33158
rect 33252 33156 33258 33158
rect 32950 33147 33258 33156
rect 27950 32668 28258 32677
rect 27950 32666 27956 32668
rect 28012 32666 28036 32668
rect 28092 32666 28116 32668
rect 28172 32666 28196 32668
rect 28252 32666 28258 32668
rect 28012 32614 28014 32666
rect 28194 32614 28196 32666
rect 27950 32612 27956 32614
rect 28012 32612 28036 32614
rect 28092 32612 28116 32614
rect 28172 32612 28196 32614
rect 28252 32612 28258 32614
rect 27950 32603 28258 32612
rect 32950 32124 33258 32133
rect 32950 32122 32956 32124
rect 33012 32122 33036 32124
rect 33092 32122 33116 32124
rect 33172 32122 33196 32124
rect 33252 32122 33258 32124
rect 33012 32070 33014 32122
rect 33194 32070 33196 32122
rect 32950 32068 32956 32070
rect 33012 32068 33036 32070
rect 33092 32068 33116 32070
rect 33172 32068 33196 32070
rect 33252 32068 33258 32070
rect 32950 32059 33258 32068
rect 24400 31884 24452 31890
rect 24400 31826 24452 31832
rect 24768 31884 24820 31890
rect 24768 31826 24820 31832
rect 24308 27396 24360 27402
rect 24308 27338 24360 27344
rect 24216 27328 24268 27334
rect 24216 27270 24268 27276
rect 24032 23316 24084 23322
rect 24032 23258 24084 23264
rect 24044 20398 24072 23258
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 23768 19922 23796 20334
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2596 8832 2648 8838
rect 3436 8809 3464 9590
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 2596 8774 2648 8780
rect 3422 8800 3478 8809
rect 2608 3058 2636 8774
rect 3422 8735 3478 8744
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 3988 3194 4016 3402
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1504 800 1532 2382
rect 2240 800 2268 2926
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2976 800 3004 2382
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 3436 1873 3464 1974
rect 3422 1864 3478 1873
rect 3422 1799 3478 1808
rect 3712 800 3740 2994
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 4448 800 4476 2314
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 4724 1970 4752 2246
rect 4712 1964 4764 1970
rect 4712 1906 4764 1912
rect 5184 800 5212 2314
rect 5552 1902 5580 2314
rect 5540 1896 5592 1902
rect 5540 1838 5592 1844
rect 5920 800 5948 2314
rect 6656 800 6684 2994
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6748 1562 6776 2246
rect 6736 1556 6788 1562
rect 6736 1498 6788 1504
rect 7392 800 7420 2382
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7484 2106 7512 2246
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 8312 1442 8340 2314
rect 8128 1414 8340 1442
rect 8128 800 8156 1414
rect 8864 800 8892 2994
rect 10612 2514 10640 4762
rect 11704 4548 11756 4554
rect 11704 4490 11756 4496
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10324 2440 10376 2446
rect 9862 2408 9918 2417
rect 9588 2372 9640 2378
rect 10324 2382 10376 2388
rect 9862 2343 9864 2352
rect 9588 2314 9640 2320
rect 9916 2343 9918 2352
rect 9864 2314 9916 2320
rect 9600 800 9628 2314
rect 10336 800 10364 2382
rect 11072 800 11100 2994
rect 11716 2650 11744 4490
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13372 3058 13400 11290
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13464 4554 13492 4694
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14384 3058 14412 3606
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11808 800 11836 2382
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 1834 11928 2246
rect 11888 1828 11940 1834
rect 11888 1770 11940 1776
rect 12544 800 12572 2926
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13280 800 13308 2450
rect 14016 800 14044 2926
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 14752 800 14780 2382
rect 15488 800 15516 2382
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16132 1766 16160 2246
rect 16120 1760 16172 1766
rect 16120 1702 16172 1708
rect 16224 870 16344 898
rect 16224 800 16252 870
rect 1490 0 1546 800
rect 2226 0 2282 800
rect 2962 0 3018 800
rect 3698 0 3754 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7378 0 7434 800
rect 8114 0 8170 800
rect 8850 0 8906 800
rect 9586 0 9642 800
rect 10322 0 10378 800
rect 11058 0 11114 800
rect 11794 0 11850 800
rect 12530 0 12586 800
rect 13266 0 13322 800
rect 14002 0 14058 800
rect 14738 0 14794 800
rect 15474 0 15530 800
rect 16210 0 16266 800
rect 16316 762 16344 870
rect 16500 762 16528 2382
rect 16960 800 16988 3470
rect 17236 2106 17264 12922
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 2106 17356 2246
rect 17224 2100 17276 2106
rect 17224 2042 17276 2048
rect 17316 2100 17368 2106
rect 17316 2042 17368 2048
rect 17224 1964 17276 1970
rect 17224 1906 17276 1912
rect 17236 1698 17264 1906
rect 17224 1692 17276 1698
rect 17224 1634 17276 1640
rect 17696 800 17724 2926
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18432 800 18460 2450
rect 18524 1902 18552 8502
rect 18616 3126 18644 13126
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 18512 1896 18564 1902
rect 18512 1838 18564 1844
rect 19168 800 19196 2926
rect 19812 2582 19840 17070
rect 21008 16794 21036 17138
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23308 15706 23336 19314
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23584 16046 23612 16594
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20088 13326 20116 13670
rect 20364 13530 20392 13670
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 21468 12986 21496 13330
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 23308 12918 23336 13194
rect 23400 12986 23428 15370
rect 23584 15094 23612 15982
rect 23572 15088 23624 15094
rect 23492 15048 23572 15076
rect 23492 14074 23520 15048
rect 23572 15030 23624 15036
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23308 12434 23336 12854
rect 23492 12782 23520 13670
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23308 12406 23428 12434
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19800 2576 19852 2582
rect 19800 2518 19852 2524
rect 19904 800 19932 3470
rect 19996 2446 20024 11222
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22756 9178 22784 9522
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 23308 8906 23336 9318
rect 23296 8900 23348 8906
rect 23296 8842 23348 8848
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 20258 3632 20314 3641
rect 20258 3567 20260 3576
rect 20312 3567 20314 3576
rect 20260 3538 20312 3544
rect 20916 2990 20944 3674
rect 22020 3194 22048 8298
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 20640 800 20668 2926
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21192 1970 21220 2314
rect 21180 1964 21232 1970
rect 21180 1906 21232 1912
rect 21376 800 21404 2314
rect 22112 800 22140 2926
rect 22388 2922 22416 2994
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 22284 2304 22336 2310
rect 22284 2246 22336 2252
rect 22296 1834 22324 2246
rect 22284 1828 22336 1834
rect 22284 1770 22336 1776
rect 22848 800 22876 2382
rect 23400 1562 23428 12406
rect 23492 11898 23520 12718
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23492 8634 23520 8774
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23676 3466 23704 18226
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23860 15570 23888 16730
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23860 14482 23888 15506
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23860 14074 23888 14418
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23768 11694 23796 14010
rect 24044 13190 24072 20334
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24136 16454 24164 19246
rect 24124 16448 24176 16454
rect 24124 16390 24176 16396
rect 24136 16182 24164 16390
rect 24124 16176 24176 16182
rect 24124 16118 24176 16124
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 23940 9444 23992 9450
rect 23940 9386 23992 9392
rect 23952 8634 23980 9386
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23664 3460 23716 3466
rect 23664 3402 23716 3408
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23388 1556 23440 1562
rect 23388 1498 23440 1504
rect 23584 800 23612 2382
rect 23860 2106 23888 7686
rect 24044 4758 24072 11630
rect 24412 9654 24440 31826
rect 27950 31580 28258 31589
rect 27950 31578 27956 31580
rect 28012 31578 28036 31580
rect 28092 31578 28116 31580
rect 28172 31578 28196 31580
rect 28252 31578 28258 31580
rect 28012 31526 28014 31578
rect 28194 31526 28196 31578
rect 27950 31524 27956 31526
rect 28012 31524 28036 31526
rect 28092 31524 28116 31526
rect 28172 31524 28196 31526
rect 28252 31524 28258 31526
rect 27950 31515 28258 31524
rect 31484 31204 31536 31210
rect 31484 31146 31536 31152
rect 27950 30492 28258 30501
rect 27950 30490 27956 30492
rect 28012 30490 28036 30492
rect 28092 30490 28116 30492
rect 28172 30490 28196 30492
rect 28252 30490 28258 30492
rect 28012 30438 28014 30490
rect 28194 30438 28196 30490
rect 27950 30436 27956 30438
rect 28012 30436 28036 30438
rect 28092 30436 28116 30438
rect 28172 30436 28196 30438
rect 28252 30436 28258 30438
rect 27950 30427 28258 30436
rect 27950 29404 28258 29413
rect 27950 29402 27956 29404
rect 28012 29402 28036 29404
rect 28092 29402 28116 29404
rect 28172 29402 28196 29404
rect 28252 29402 28258 29404
rect 28012 29350 28014 29402
rect 28194 29350 28196 29402
rect 27950 29348 27956 29350
rect 28012 29348 28036 29350
rect 28092 29348 28116 29350
rect 28172 29348 28196 29350
rect 28252 29348 28258 29350
rect 27950 29339 28258 29348
rect 31392 29300 31444 29306
rect 31392 29242 31444 29248
rect 30288 29096 30340 29102
rect 30288 29038 30340 29044
rect 27950 28316 28258 28325
rect 27950 28314 27956 28316
rect 28012 28314 28036 28316
rect 28092 28314 28116 28316
rect 28172 28314 28196 28316
rect 28252 28314 28258 28316
rect 28012 28262 28014 28314
rect 28194 28262 28196 28314
rect 27950 28260 27956 28262
rect 28012 28260 28036 28262
rect 28092 28260 28116 28262
rect 28172 28260 28196 28262
rect 28252 28260 28258 28262
rect 27950 28251 28258 28260
rect 25596 28144 25648 28150
rect 25596 28086 25648 28092
rect 28816 28144 28868 28150
rect 28816 28086 28868 28092
rect 30104 28144 30156 28150
rect 30104 28086 30156 28092
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 24768 27396 24820 27402
rect 24768 27338 24820 27344
rect 24780 26790 24808 27338
rect 24768 26784 24820 26790
rect 24768 26726 24820 26732
rect 25228 26308 25280 26314
rect 25228 26250 25280 26256
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24872 23186 24900 25434
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 24596 22166 24624 23054
rect 24584 22160 24636 22166
rect 24584 22102 24636 22108
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 24964 20942 24992 21286
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 24768 16516 24820 16522
rect 24768 16458 24820 16464
rect 24780 16046 24808 16458
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24504 15570 24532 15982
rect 24492 15564 24544 15570
rect 24492 15506 24544 15512
rect 24780 15026 24808 15982
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24780 14006 24808 14962
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24596 11354 24624 12174
rect 24688 11694 24716 13670
rect 24780 13138 24808 13942
rect 24872 13258 24900 17070
rect 24964 13530 24992 18566
rect 25056 18358 25084 20742
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 25148 17338 25176 21286
rect 25240 21010 25268 26250
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25424 22094 25452 23122
rect 25332 22066 25452 22094
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25332 20584 25360 22066
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 25424 20942 25452 21966
rect 25516 21690 25544 28018
rect 25608 23866 25636 28086
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 27528 28008 27580 28014
rect 27528 27950 27580 27956
rect 26148 27668 26200 27674
rect 26148 27610 26200 27616
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 26160 23662 26188 27610
rect 27344 26580 27396 26586
rect 27344 26522 27396 26528
rect 26424 25832 26476 25838
rect 26424 25774 26476 25780
rect 26056 23656 26108 23662
rect 26056 23598 26108 23604
rect 26148 23656 26200 23662
rect 26148 23598 26200 23604
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25412 20936 25464 20942
rect 25412 20878 25464 20884
rect 25240 20556 25360 20584
rect 25240 18222 25268 20556
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25332 19786 25360 20402
rect 25424 20398 25452 20878
rect 25412 20392 25464 20398
rect 25412 20334 25464 20340
rect 25424 19922 25452 20334
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25320 19780 25372 19786
rect 25320 19722 25372 19728
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25240 17814 25268 18158
rect 25228 17808 25280 17814
rect 25228 17750 25280 17756
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25228 16788 25280 16794
rect 25228 16730 25280 16736
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 24780 13110 24900 13138
rect 24872 12918 24900 13110
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24872 12782 24900 12854
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24780 12374 24808 12718
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24780 11642 24808 12310
rect 25056 12306 25084 14826
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24780 11614 24900 11642
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 24136 8430 24164 8978
rect 24780 8974 24808 11494
rect 24872 11354 24900 11614
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 23848 2100 23900 2106
rect 23848 2042 23900 2048
rect 24320 800 24348 3538
rect 24688 3534 24716 4966
rect 24780 4622 24808 8910
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24584 2576 24636 2582
rect 24584 2518 24636 2524
rect 24596 2310 24624 2518
rect 24584 2304 24636 2310
rect 24584 2246 24636 2252
rect 24964 1902 24992 12038
rect 25148 11762 25176 12718
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 25148 8566 25176 9454
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24952 1896 25004 1902
rect 24952 1838 25004 1844
rect 25056 800 25084 2926
rect 25240 2446 25268 16730
rect 25332 14618 25360 19314
rect 25424 17746 25452 19858
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25412 17740 25464 17746
rect 25412 17682 25464 17688
rect 25516 15434 25544 18770
rect 26068 18426 26096 23598
rect 26160 23322 26188 23598
rect 26148 23316 26200 23322
rect 26148 23258 26200 23264
rect 26160 21486 26188 23258
rect 26436 22094 26464 25774
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 27080 23866 27108 24550
rect 27160 24336 27212 24342
rect 27160 24278 27212 24284
rect 27068 23860 27120 23866
rect 27068 23802 27120 23808
rect 26608 23044 26660 23050
rect 26608 22986 26660 22992
rect 26700 23044 26752 23050
rect 26700 22986 26752 22992
rect 26344 22066 26464 22094
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26252 19718 26280 20198
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26252 18834 26280 19654
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 26344 18714 26372 22066
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26436 21010 26464 21830
rect 26620 21690 26648 22986
rect 26608 21684 26660 21690
rect 26608 21626 26660 21632
rect 26712 21570 26740 22986
rect 26792 22092 26844 22098
rect 26792 22034 26844 22040
rect 26620 21542 26740 21570
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26424 21004 26476 21010
rect 26424 20946 26476 20952
rect 26252 18686 26372 18714
rect 26056 18420 26108 18426
rect 26056 18362 26108 18368
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25596 18080 25648 18086
rect 25596 18022 25648 18028
rect 25608 17338 25636 18022
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25700 16658 25728 17818
rect 25976 17338 26004 18226
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 26252 17202 26280 18686
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 25504 15428 25556 15434
rect 25504 15370 25556 15376
rect 25516 15162 25544 15370
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25504 14952 25556 14958
rect 25504 14894 25556 14900
rect 25320 14612 25372 14618
rect 25320 14554 25372 14560
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 25332 12986 25360 13942
rect 25516 13394 25544 14894
rect 25504 13388 25556 13394
rect 25504 13330 25556 13336
rect 25412 13184 25464 13190
rect 25412 13126 25464 13132
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25332 11218 25360 12922
rect 25424 12442 25452 13126
rect 25516 12646 25544 13330
rect 25504 12640 25556 12646
rect 25504 12582 25556 12588
rect 25412 12436 25464 12442
rect 25792 12434 25820 16526
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25884 14074 25912 15302
rect 26252 15094 26280 15506
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26252 14074 26280 14350
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 26240 14068 26292 14074
rect 26240 14010 26292 14016
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 25412 12378 25464 12384
rect 25700 12406 25820 12434
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25332 10130 25360 11154
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25318 5128 25374 5137
rect 25318 5063 25374 5072
rect 25332 3058 25360 5063
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25700 1698 25728 12406
rect 26148 12096 26200 12102
rect 26148 12038 26200 12044
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 25792 8566 25820 10066
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25792 7954 25820 8502
rect 26160 8294 26188 12038
rect 26252 11218 26280 13874
rect 26344 13530 26372 18566
rect 26436 13802 26464 18566
rect 26528 16590 26556 21422
rect 26620 20330 26648 21542
rect 26700 21412 26752 21418
rect 26700 21354 26752 21360
rect 26608 20324 26660 20330
rect 26608 20266 26660 20272
rect 26620 19718 26648 20266
rect 26608 19712 26660 19718
rect 26608 19654 26660 19660
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26620 16266 26648 19654
rect 26712 16454 26740 21354
rect 26804 16522 26832 22034
rect 27068 21956 27120 21962
rect 27068 21898 27120 21904
rect 27080 21706 27108 21898
rect 26896 21690 27108 21706
rect 26884 21684 27108 21690
rect 26936 21678 27108 21684
rect 26884 21626 26936 21632
rect 26896 20874 26924 21626
rect 26976 21616 27028 21622
rect 26976 21558 27028 21564
rect 26884 20868 26936 20874
rect 26884 20810 26936 20816
rect 26896 20466 26924 20810
rect 26884 20460 26936 20466
rect 26884 20402 26936 20408
rect 26792 16516 26844 16522
rect 26792 16458 26844 16464
rect 26700 16448 26752 16454
rect 26700 16390 26752 16396
rect 26620 16238 26740 16266
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26424 13796 26476 13802
rect 26424 13738 26476 13744
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26424 13456 26476 13462
rect 26424 13398 26476 13404
rect 26436 13190 26464 13398
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26528 11898 26556 14214
rect 26620 12714 26648 14214
rect 26712 13190 26740 16238
rect 26988 15706 27016 21558
rect 27172 17270 27200 24278
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 27264 18766 27292 22918
rect 27356 21418 27384 26522
rect 27436 26444 27488 26450
rect 27436 26386 27488 26392
rect 27448 25974 27476 26386
rect 27436 25968 27488 25974
rect 27436 25910 27488 25916
rect 27540 25838 27568 27950
rect 28460 27538 28488 28018
rect 28448 27532 28500 27538
rect 28448 27474 28500 27480
rect 27950 27228 28258 27237
rect 27950 27226 27956 27228
rect 28012 27226 28036 27228
rect 28092 27226 28116 27228
rect 28172 27226 28196 27228
rect 28252 27226 28258 27228
rect 28012 27174 28014 27226
rect 28194 27174 28196 27226
rect 27950 27172 27956 27174
rect 28012 27172 28036 27174
rect 28092 27172 28116 27174
rect 28172 27172 28196 27174
rect 28252 27172 28258 27174
rect 27950 27163 28258 27172
rect 28460 26994 28488 27474
rect 28448 26988 28500 26994
rect 28448 26930 28500 26936
rect 27712 26852 27764 26858
rect 27712 26794 27764 26800
rect 27724 26314 27752 26794
rect 28172 26784 28224 26790
rect 28172 26726 28224 26732
rect 28184 26330 28212 26726
rect 28460 26450 28488 26930
rect 28448 26444 28500 26450
rect 28448 26386 28500 26392
rect 28184 26314 28580 26330
rect 27712 26308 27764 26314
rect 27712 26250 27764 26256
rect 28172 26308 28580 26314
rect 28224 26302 28580 26308
rect 28172 26250 28224 26256
rect 27950 26140 28258 26149
rect 27950 26138 27956 26140
rect 28012 26138 28036 26140
rect 28092 26138 28116 26140
rect 28172 26138 28196 26140
rect 28252 26138 28258 26140
rect 28012 26086 28014 26138
rect 28194 26086 28196 26138
rect 27950 26084 27956 26086
rect 28012 26084 28036 26086
rect 28092 26084 28116 26086
rect 28172 26084 28196 26086
rect 28252 26084 28258 26086
rect 27950 26075 28258 26084
rect 28552 25906 28580 26302
rect 28540 25900 28592 25906
rect 28540 25842 28592 25848
rect 27528 25832 27580 25838
rect 27528 25774 27580 25780
rect 27950 25052 28258 25061
rect 27950 25050 27956 25052
rect 28012 25050 28036 25052
rect 28092 25050 28116 25052
rect 28172 25050 28196 25052
rect 28252 25050 28258 25052
rect 28012 24998 28014 25050
rect 28194 24998 28196 25050
rect 27950 24996 27956 24998
rect 28012 24996 28036 24998
rect 28092 24996 28116 24998
rect 28172 24996 28196 24998
rect 28252 24996 28258 24998
rect 27950 24987 28258 24996
rect 27528 24268 27580 24274
rect 27528 24210 27580 24216
rect 27540 21894 27568 24210
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27344 21412 27396 21418
rect 27344 21354 27396 21360
rect 27540 21146 27568 21490
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27528 20528 27580 20534
rect 27528 20470 27580 20476
rect 27540 19718 27568 20470
rect 27632 19786 27660 22714
rect 27816 21894 27844 24074
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 28552 23730 28580 25842
rect 28724 25764 28776 25770
rect 28724 25706 28776 25712
rect 28736 25498 28764 25706
rect 28828 25702 28856 28086
rect 28908 27872 28960 27878
rect 28908 27814 28960 27820
rect 28816 25696 28868 25702
rect 28816 25638 28868 25644
rect 28724 25492 28776 25498
rect 28724 25434 28776 25440
rect 28828 24342 28856 25638
rect 28816 24336 28868 24342
rect 28816 24278 28868 24284
rect 28920 24274 28948 27814
rect 30116 27062 30144 28086
rect 30300 27878 30328 29038
rect 30656 28620 30708 28626
rect 30656 28562 30708 28568
rect 30472 28484 30524 28490
rect 30472 28426 30524 28432
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30300 27130 30328 27814
rect 30288 27124 30340 27130
rect 30288 27066 30340 27072
rect 30104 27056 30156 27062
rect 30104 26998 30156 27004
rect 30104 26852 30156 26858
rect 30104 26794 30156 26800
rect 29000 25696 29052 25702
rect 29000 25638 29052 25644
rect 29012 24614 29040 25638
rect 29460 24744 29512 24750
rect 29460 24686 29512 24692
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 28908 24268 28960 24274
rect 28908 24210 28960 24216
rect 28632 24064 28684 24070
rect 28632 24006 28684 24012
rect 29368 24064 29420 24070
rect 29368 24006 29420 24012
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28552 23594 28580 23666
rect 28540 23588 28592 23594
rect 28540 23530 28592 23536
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27804 21888 27856 21894
rect 27804 21830 27856 21836
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27528 19712 27580 19718
rect 27528 19654 27580 19660
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 27448 18698 27476 19314
rect 27436 18692 27488 18698
rect 27436 18634 27488 18640
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27160 17264 27212 17270
rect 27160 17206 27212 17212
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 26804 13734 26832 14418
rect 26976 14408 27028 14414
rect 26974 14376 26976 14385
rect 27028 14376 27030 14385
rect 26974 14311 27030 14320
rect 26884 14272 26936 14278
rect 26884 14214 26936 14220
rect 26792 13728 26844 13734
rect 26792 13670 26844 13676
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26804 13326 26832 13466
rect 26896 13326 26924 14214
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 26700 13184 26752 13190
rect 26700 13126 26752 13132
rect 26700 12776 26752 12782
rect 26700 12718 26752 12724
rect 26608 12708 26660 12714
rect 26608 12650 26660 12656
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26608 11756 26660 11762
rect 26608 11698 26660 11704
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 26620 11082 26648 11698
rect 26608 11076 26660 11082
rect 26608 11018 26660 11024
rect 26620 9994 26648 11018
rect 26608 9988 26660 9994
rect 26608 9930 26660 9936
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26436 8498 26464 9318
rect 26620 8906 26648 9930
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 26620 8498 26648 8842
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26608 8492 26660 8498
rect 26608 8434 26660 8440
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 25688 1692 25740 1698
rect 25688 1634 25740 1640
rect 25792 800 25820 2450
rect 26252 1766 26280 8366
rect 26620 8242 26648 8434
rect 26712 8430 26740 12718
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 26620 8214 26832 8242
rect 26804 7818 26832 8214
rect 26792 7812 26844 7818
rect 26792 7754 26844 7760
rect 26804 4554 26832 7754
rect 26896 4826 26924 13262
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 26988 12714 27016 13126
rect 26976 12708 27028 12714
rect 26976 12650 27028 12656
rect 27080 12442 27108 16390
rect 27068 12436 27120 12442
rect 27068 12378 27120 12384
rect 27172 10810 27200 16594
rect 27356 16522 27384 17546
rect 27344 16516 27396 16522
rect 27344 16458 27396 16464
rect 27356 16182 27384 16458
rect 27344 16176 27396 16182
rect 27344 16118 27396 16124
rect 27356 15434 27384 16118
rect 27344 15428 27396 15434
rect 27344 15370 27396 15376
rect 27448 15026 27476 18634
rect 27632 17882 27660 19722
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27632 16776 27660 17682
rect 27724 17542 27752 20810
rect 27816 19922 27844 21422
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27804 19916 27856 19922
rect 27804 19858 27856 19864
rect 27816 19446 27844 19858
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27804 19440 27856 19446
rect 27804 19382 27856 19388
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 28644 18426 28672 24006
rect 29380 23662 29408 24006
rect 29368 23656 29420 23662
rect 29368 23598 29420 23604
rect 29472 23594 29500 24686
rect 29736 24200 29788 24206
rect 29736 24142 29788 24148
rect 29748 23866 29776 24142
rect 29736 23860 29788 23866
rect 29736 23802 29788 23808
rect 29000 23588 29052 23594
rect 29000 23530 29052 23536
rect 29460 23588 29512 23594
rect 29460 23530 29512 23536
rect 28908 23520 28960 23526
rect 28908 23462 28960 23468
rect 28920 23186 28948 23462
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 29012 21622 29040 23530
rect 29184 22160 29236 22166
rect 29184 22102 29236 22108
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 28724 21480 28776 21486
rect 28724 21422 28776 21428
rect 28736 20602 28764 21422
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 28736 19242 28764 20538
rect 29196 20058 29224 22102
rect 29276 20800 29328 20806
rect 29276 20742 29328 20748
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 28908 19916 28960 19922
rect 28908 19858 28960 19864
rect 28920 19514 28948 19858
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 28816 19372 28868 19378
rect 28816 19314 28868 19320
rect 28724 19236 28776 19242
rect 28724 19178 28776 19184
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 28632 18420 28684 18426
rect 28632 18362 28684 18368
rect 28448 18284 28500 18290
rect 28448 18226 28500 18232
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 27724 17066 27752 17478
rect 27816 17134 27844 18158
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27804 17128 27856 17134
rect 27804 17070 27856 17076
rect 27712 17060 27764 17066
rect 27712 17002 27764 17008
rect 27540 16748 27752 16776
rect 27540 16658 27568 16748
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27540 15026 27568 15982
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27448 14414 27476 14962
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27344 14340 27396 14346
rect 27344 14282 27396 14288
rect 27252 13796 27304 13802
rect 27252 13738 27304 13744
rect 27264 12850 27292 13738
rect 27356 12986 27384 14282
rect 27540 13938 27568 14962
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27528 13728 27580 13734
rect 27528 13670 27580 13676
rect 27540 13462 27568 13670
rect 27528 13456 27580 13462
rect 27528 13398 27580 13404
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27264 11830 27292 12786
rect 27632 12481 27660 16594
rect 27724 16250 27752 16748
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 27712 16040 27764 16046
rect 27712 15982 27764 15988
rect 27724 14482 27752 15982
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27724 13938 27752 14418
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27816 13818 27844 17070
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 28276 15570 28304 16186
rect 28264 15564 28316 15570
rect 28264 15506 28316 15512
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 28264 14816 28316 14822
rect 28262 14784 28264 14793
rect 28316 14784 28318 14793
rect 28262 14719 28318 14728
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 28172 14068 28224 14074
rect 28172 14010 28224 14016
rect 27724 13790 27844 13818
rect 27618 12472 27674 12481
rect 27618 12407 27674 12416
rect 27620 12368 27672 12374
rect 27620 12310 27672 12316
rect 27252 11824 27304 11830
rect 27252 11766 27304 11772
rect 27632 11558 27660 12310
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27160 10804 27212 10810
rect 27160 10746 27212 10752
rect 27528 9920 27580 9926
rect 27528 9862 27580 9868
rect 27068 9104 27120 9110
rect 27068 9046 27120 9052
rect 27080 7954 27108 9046
rect 27540 9042 27568 9862
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27528 8560 27580 8566
rect 27580 8508 27660 8514
rect 27528 8502 27660 8508
rect 27540 8486 27660 8502
rect 27632 8430 27660 8486
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 27068 7948 27120 7954
rect 27068 7890 27120 7896
rect 27528 5568 27580 5574
rect 27528 5510 27580 5516
rect 26884 4820 26936 4826
rect 26884 4762 26936 4768
rect 26792 4548 26844 4554
rect 26792 4490 26844 4496
rect 27540 3058 27568 5510
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 27252 2984 27304 2990
rect 27252 2926 27304 2932
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26240 1760 26292 1766
rect 26240 1702 26292 1708
rect 26528 800 26556 2450
rect 27264 800 27292 2926
rect 27724 1970 27752 13790
rect 28184 13734 28212 14010
rect 28080 13728 28132 13734
rect 28080 13670 28132 13676
rect 28172 13728 28224 13734
rect 28172 13670 28224 13676
rect 28092 13394 28120 13670
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 28092 13246 28304 13274
rect 27816 12646 27844 13194
rect 28092 13190 28120 13246
rect 28276 13190 28304 13246
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 28368 12866 28396 17478
rect 28460 14618 28488 18226
rect 28736 17678 28764 18702
rect 28724 17672 28776 17678
rect 28724 17614 28776 17620
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28552 17338 28580 17478
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 28540 17128 28592 17134
rect 28540 17070 28592 17076
rect 28632 17128 28684 17134
rect 28632 17070 28684 17076
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28448 14408 28500 14414
rect 28448 14350 28500 14356
rect 28460 13530 28488 14350
rect 28552 13870 28580 17070
rect 28644 16658 28672 17070
rect 28724 17060 28776 17066
rect 28724 17002 28776 17008
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28736 16046 28764 17002
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28736 15502 28764 15982
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28736 14328 28764 15438
rect 28828 14414 28856 19314
rect 29196 18222 29224 19994
rect 29184 18216 29236 18222
rect 29184 18158 29236 18164
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28920 16046 28948 17818
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 29012 16590 29040 17614
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 29092 16992 29144 16998
rect 29092 16934 29144 16940
rect 29104 16726 29132 16934
rect 29196 16794 29224 17206
rect 29184 16788 29236 16794
rect 29184 16730 29236 16736
rect 29092 16720 29144 16726
rect 29092 16662 29144 16668
rect 29000 16584 29052 16590
rect 29000 16526 29052 16532
rect 29288 16454 29316 20742
rect 29368 18896 29420 18902
rect 29368 18838 29420 18844
rect 29276 16448 29328 16454
rect 29276 16390 29328 16396
rect 28908 16040 28960 16046
rect 28908 15982 28960 15988
rect 28920 14482 28948 15982
rect 28908 14476 28960 14482
rect 28908 14418 28960 14424
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28644 14300 28764 14328
rect 28540 13864 28592 13870
rect 28540 13806 28592 13812
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 28276 12838 28396 12866
rect 27896 12776 27948 12782
rect 28080 12776 28132 12782
rect 27948 12724 28080 12730
rect 27896 12718 28132 12724
rect 27908 12702 28120 12718
rect 27804 12640 27856 12646
rect 27804 12582 27856 12588
rect 27802 12472 27858 12481
rect 27802 12407 27858 12416
rect 27816 2854 27844 12407
rect 28172 12368 28224 12374
rect 28170 12336 28172 12345
rect 28224 12336 28226 12345
rect 28170 12271 28226 12280
rect 28276 12170 28304 12838
rect 28356 12640 28408 12646
rect 28356 12582 28408 12588
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 28368 11898 28396 12582
rect 28448 12300 28500 12306
rect 28448 12242 28500 12248
rect 28356 11892 28408 11898
rect 28356 11834 28408 11840
rect 28354 11792 28410 11801
rect 28354 11727 28410 11736
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 28368 9110 28396 11727
rect 28460 10538 28488 12242
rect 28448 10532 28500 10538
rect 28448 10474 28500 10480
rect 28356 9104 28408 9110
rect 28356 9046 28408 9052
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27896 8288 27948 8294
rect 27896 8230 27948 8236
rect 27908 8090 27936 8230
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 28552 7478 28580 13670
rect 28644 12646 28672 14300
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28644 11218 28672 12582
rect 28736 12374 28764 13806
rect 28724 12368 28776 12374
rect 28724 12310 28776 12316
rect 28724 12232 28776 12238
rect 28724 12174 28776 12180
rect 28736 11898 28764 12174
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28828 11354 28856 14214
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28630 10704 28686 10713
rect 28630 10639 28686 10648
rect 28724 10668 28776 10674
rect 28644 7954 28672 10639
rect 28724 10610 28776 10616
rect 28736 10266 28764 10610
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28724 10260 28776 10266
rect 28724 10202 28776 10208
rect 28828 9466 28856 10542
rect 28920 10470 28948 14214
rect 29380 13734 29408 18838
rect 29472 17202 29500 23530
rect 29748 22030 29776 23802
rect 30116 23118 30144 26794
rect 30484 26586 30512 28426
rect 30668 28218 30696 28562
rect 30656 28212 30708 28218
rect 30656 28154 30708 28160
rect 30668 27538 30696 28154
rect 30656 27532 30708 27538
rect 30656 27474 30708 27480
rect 30668 27282 30696 27474
rect 30576 27254 30696 27282
rect 30840 27328 30892 27334
rect 30840 27270 30892 27276
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 30484 25430 30512 26522
rect 30576 26450 30604 27254
rect 30656 26784 30708 26790
rect 30656 26726 30708 26732
rect 30564 26444 30616 26450
rect 30564 26386 30616 26392
rect 30472 25424 30524 25430
rect 30472 25366 30524 25372
rect 30668 25362 30696 26726
rect 30852 26450 30880 27270
rect 31404 27130 31432 29242
rect 31496 28218 31524 31146
rect 32950 31036 33258 31045
rect 32950 31034 32956 31036
rect 33012 31034 33036 31036
rect 33092 31034 33116 31036
rect 33172 31034 33196 31036
rect 33252 31034 33258 31036
rect 33012 30982 33014 31034
rect 33194 30982 33196 31034
rect 32950 30980 32956 30982
rect 33012 30980 33036 30982
rect 33092 30980 33116 30982
rect 33172 30980 33196 30982
rect 33252 30980 33258 30982
rect 32950 30971 33258 30980
rect 32864 30660 32916 30666
rect 32864 30602 32916 30608
rect 33508 30660 33560 30666
rect 33508 30602 33560 30608
rect 32680 29640 32732 29646
rect 32680 29582 32732 29588
rect 31668 29504 31720 29510
rect 31668 29446 31720 29452
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 31484 28212 31536 28218
rect 31484 28154 31536 28160
rect 31588 27130 31616 28970
rect 31680 28014 31708 29446
rect 31944 28484 31996 28490
rect 31944 28426 31996 28432
rect 31956 28150 31984 28426
rect 32036 28416 32088 28422
rect 32036 28358 32088 28364
rect 31944 28144 31996 28150
rect 31944 28086 31996 28092
rect 31668 28008 31720 28014
rect 31668 27950 31720 27956
rect 31956 27452 31984 28086
rect 32048 27674 32076 28358
rect 32692 27674 32720 29582
rect 32876 28490 32904 30602
rect 32950 29948 33258 29957
rect 32950 29946 32956 29948
rect 33012 29946 33036 29948
rect 33092 29946 33116 29948
rect 33172 29946 33196 29948
rect 33252 29946 33258 29948
rect 33012 29894 33014 29946
rect 33194 29894 33196 29946
rect 32950 29892 32956 29894
rect 33012 29892 33036 29894
rect 33092 29892 33116 29894
rect 33172 29892 33196 29894
rect 33252 29892 33258 29894
rect 32950 29883 33258 29892
rect 33520 29714 33548 30602
rect 33508 29708 33560 29714
rect 33508 29650 33560 29656
rect 33324 29572 33376 29578
rect 33324 29514 33376 29520
rect 32950 28860 33258 28869
rect 32950 28858 32956 28860
rect 33012 28858 33036 28860
rect 33092 28858 33116 28860
rect 33172 28858 33196 28860
rect 33252 28858 33258 28860
rect 33012 28806 33014 28858
rect 33194 28806 33196 28858
rect 32950 28804 32956 28806
rect 33012 28804 33036 28806
rect 33092 28804 33116 28806
rect 33172 28804 33196 28806
rect 33252 28804 33258 28806
rect 32950 28795 33258 28804
rect 32864 28484 32916 28490
rect 32864 28426 32916 28432
rect 32876 28218 32904 28426
rect 32864 28212 32916 28218
rect 32864 28154 32916 28160
rect 32036 27668 32088 27674
rect 32036 27610 32088 27616
rect 32680 27668 32732 27674
rect 32680 27610 32732 27616
rect 32220 27600 32272 27606
rect 32220 27542 32272 27548
rect 32128 27464 32180 27470
rect 31956 27424 32128 27452
rect 32128 27406 32180 27412
rect 31392 27124 31444 27130
rect 31392 27066 31444 27072
rect 31576 27124 31628 27130
rect 31576 27066 31628 27072
rect 31484 26580 31536 26586
rect 31484 26522 31536 26528
rect 30840 26444 30892 26450
rect 30840 26386 30892 26392
rect 30656 25356 30708 25362
rect 30656 25298 30708 25304
rect 30380 25220 30432 25226
rect 30380 25162 30432 25168
rect 31300 25220 31352 25226
rect 31300 25162 31352 25168
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 29736 22024 29788 22030
rect 29736 21966 29788 21972
rect 29748 20942 29776 21966
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29644 20528 29696 20534
rect 29644 20470 29696 20476
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29656 16658 29684 20470
rect 29748 20398 29776 20878
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29748 19310 29776 20334
rect 30116 19514 30144 22918
rect 30196 22228 30248 22234
rect 30196 22170 30248 22176
rect 30208 21350 30236 22170
rect 30392 21690 30420 25162
rect 30564 25152 30616 25158
rect 30564 25094 30616 25100
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 30472 21616 30524 21622
rect 30472 21558 30524 21564
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30104 19508 30156 19514
rect 30104 19450 30156 19456
rect 29736 19304 29788 19310
rect 29736 19246 29788 19252
rect 29748 18834 29776 19246
rect 29736 18828 29788 18834
rect 29736 18770 29788 18776
rect 29748 18222 29776 18770
rect 30208 18358 30236 21286
rect 30288 21140 30340 21146
rect 30288 21082 30340 21088
rect 30300 20534 30328 21082
rect 30288 20528 30340 20534
rect 30288 20470 30340 20476
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30392 18358 30420 19110
rect 30196 18352 30248 18358
rect 30196 18294 30248 18300
rect 30380 18352 30432 18358
rect 30380 18294 30432 18300
rect 29920 18284 29972 18290
rect 29920 18226 29972 18232
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29748 16658 29776 18158
rect 29644 16652 29696 16658
rect 29644 16594 29696 16600
rect 29736 16652 29788 16658
rect 29736 16594 29788 16600
rect 29644 16516 29696 16522
rect 29644 16458 29696 16464
rect 29656 16182 29684 16458
rect 29644 16176 29696 16182
rect 29644 16118 29696 16124
rect 29552 15428 29604 15434
rect 29552 15370 29604 15376
rect 29368 13728 29420 13734
rect 29368 13670 29420 13676
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 29092 12912 29144 12918
rect 29090 12880 29092 12889
rect 29144 12880 29146 12889
rect 29090 12815 29146 12824
rect 29368 12776 29420 12782
rect 29368 12718 29420 12724
rect 29000 12640 29052 12646
rect 29000 12582 29052 12588
rect 29012 11014 29040 12582
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 29092 11688 29144 11694
rect 29092 11630 29144 11636
rect 29104 11286 29132 11630
rect 29184 11620 29236 11626
rect 29184 11562 29236 11568
rect 29092 11280 29144 11286
rect 29092 11222 29144 11228
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 28908 10464 28960 10470
rect 28908 10406 28960 10412
rect 29092 9580 29144 9586
rect 29092 9522 29144 9528
rect 28828 9438 28948 9466
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28828 8974 28856 9318
rect 28816 8968 28868 8974
rect 28816 8910 28868 8916
rect 28632 7948 28684 7954
rect 28632 7890 28684 7896
rect 28816 7880 28868 7886
rect 28920 7868 28948 9438
rect 29000 9444 29052 9450
rect 29000 9386 29052 9392
rect 29012 8090 29040 9386
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 28868 7840 28948 7868
rect 28816 7822 28868 7828
rect 28540 7472 28592 7478
rect 28540 7414 28592 7420
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 28828 3398 28856 7822
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 27712 1964 27764 1970
rect 27712 1906 27764 1912
rect 28000 870 28120 898
rect 28000 800 28028 870
rect 16316 734 16528 762
rect 16946 0 17002 800
rect 17682 0 17738 800
rect 18418 0 18474 800
rect 19154 0 19210 800
rect 19890 0 19946 800
rect 20626 0 20682 800
rect 21362 0 21418 800
rect 22098 0 22154 800
rect 22834 0 22890 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25042 0 25098 800
rect 25778 0 25834 800
rect 26514 0 26570 800
rect 27250 0 27306 800
rect 27986 0 28042 800
rect 28092 762 28120 870
rect 28368 762 28396 2790
rect 28736 800 28764 2926
rect 29104 2774 29132 9522
rect 29196 5710 29224 11562
rect 29288 9450 29316 11698
rect 29380 11694 29408 12718
rect 29368 11688 29420 11694
rect 29368 11630 29420 11636
rect 29368 10600 29420 10606
rect 29368 10542 29420 10548
rect 29276 9444 29328 9450
rect 29276 9386 29328 9392
rect 29276 7268 29328 7274
rect 29276 7210 29328 7216
rect 29184 5704 29236 5710
rect 29184 5646 29236 5652
rect 29012 2746 29132 2774
rect 29012 2582 29040 2746
rect 29000 2576 29052 2582
rect 29000 2518 29052 2524
rect 29288 2446 29316 7210
rect 29276 2440 29328 2446
rect 29276 2382 29328 2388
rect 29380 2310 29408 10542
rect 29472 10130 29500 13670
rect 29564 12442 29592 15370
rect 29656 14006 29684 16118
rect 29828 15360 29880 15366
rect 29828 15302 29880 15308
rect 29644 14000 29696 14006
rect 29644 13942 29696 13948
rect 29656 13530 29684 13942
rect 29644 13524 29696 13530
rect 29644 13466 29696 13472
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 29552 12436 29604 12442
rect 29552 12378 29604 12384
rect 29552 11824 29604 11830
rect 29552 11766 29604 11772
rect 29564 10810 29592 11766
rect 29656 11354 29684 13126
rect 29736 12776 29788 12782
rect 29736 12718 29788 12724
rect 29644 11348 29696 11354
rect 29644 11290 29696 11296
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29656 10985 29684 11086
rect 29642 10976 29698 10985
rect 29642 10911 29698 10920
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29748 10130 29776 12718
rect 29840 11898 29868 15302
rect 29932 14074 29960 18226
rect 30392 17134 30420 18294
rect 30484 18086 30512 21558
rect 30576 21078 30604 25094
rect 31024 24608 31076 24614
rect 31024 24550 31076 24556
rect 31116 24608 31168 24614
rect 31116 24550 31168 24556
rect 30932 23520 30984 23526
rect 30932 23462 30984 23468
rect 30944 21962 30972 23462
rect 30932 21956 30984 21962
rect 30932 21898 30984 21904
rect 30840 21888 30892 21894
rect 30840 21830 30892 21836
rect 30852 21690 30880 21830
rect 30840 21684 30892 21690
rect 30840 21626 30892 21632
rect 30564 21072 30616 21078
rect 30564 21014 30616 21020
rect 30944 20874 30972 21898
rect 31036 21690 31064 24550
rect 31128 23118 31156 24550
rect 31208 24268 31260 24274
rect 31208 24210 31260 24216
rect 31220 23662 31248 24210
rect 31208 23656 31260 23662
rect 31208 23598 31260 23604
rect 31116 23112 31168 23118
rect 31116 23054 31168 23060
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 31220 21486 31248 23598
rect 31208 21480 31260 21486
rect 31208 21422 31260 21428
rect 31024 21412 31076 21418
rect 31024 21354 31076 21360
rect 31036 21010 31064 21354
rect 31024 21004 31076 21010
rect 31024 20946 31076 20952
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 30944 20534 30972 20810
rect 30932 20528 30984 20534
rect 30932 20470 30984 20476
rect 30944 19446 30972 20470
rect 30932 19440 30984 19446
rect 30932 19382 30984 19388
rect 31024 18352 31076 18358
rect 31024 18294 31076 18300
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30930 17232 30986 17241
rect 30748 17196 30800 17202
rect 30930 17167 30932 17176
rect 30748 17138 30800 17144
rect 30984 17167 30986 17176
rect 30932 17138 30984 17144
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30380 16448 30432 16454
rect 30380 16390 30432 16396
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30300 14618 30328 14894
rect 30288 14612 30340 14618
rect 30288 14554 30340 14560
rect 30196 14544 30248 14550
rect 30196 14486 30248 14492
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 30012 13456 30064 13462
rect 30012 13398 30064 13404
rect 29920 12844 29972 12850
rect 29920 12786 29972 12792
rect 29828 11892 29880 11898
rect 29828 11834 29880 11840
rect 29932 11354 29960 12786
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 29918 11248 29974 11257
rect 29828 11212 29880 11218
rect 29918 11183 29974 11192
rect 29828 11154 29880 11160
rect 29840 10198 29868 11154
rect 29932 11082 29960 11183
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 30024 10742 30052 13398
rect 30104 12232 30156 12238
rect 30104 12174 30156 12180
rect 30116 10810 30144 12174
rect 30208 12102 30236 14486
rect 30392 13394 30420 16390
rect 30472 16040 30524 16046
rect 30472 15982 30524 15988
rect 30484 13870 30512 15982
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 30668 15162 30696 15438
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30472 13864 30524 13870
rect 30472 13806 30524 13812
rect 30380 13388 30432 13394
rect 30380 13330 30432 13336
rect 30380 13184 30432 13190
rect 30380 13126 30432 13132
rect 30392 12986 30420 13126
rect 30380 12980 30432 12986
rect 30380 12922 30432 12928
rect 30470 12880 30526 12889
rect 30470 12815 30526 12824
rect 30380 12776 30432 12782
rect 30380 12718 30432 12724
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30012 10736 30064 10742
rect 30012 10678 30064 10684
rect 29828 10192 29880 10198
rect 29828 10134 29880 10140
rect 29460 10124 29512 10130
rect 29460 10066 29512 10072
rect 29736 10124 29788 10130
rect 29736 10066 29788 10072
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29460 3460 29512 3466
rect 29460 3402 29512 3408
rect 29368 2304 29420 2310
rect 29368 2246 29420 2252
rect 29472 800 29500 3402
rect 29564 3058 29592 9862
rect 29748 9042 29776 10066
rect 30024 9518 30052 10678
rect 30208 10538 30236 12038
rect 30300 11914 30328 12242
rect 30392 12102 30420 12718
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30300 11886 30420 11914
rect 30392 11830 30420 11886
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30196 10532 30248 10538
rect 30196 10474 30248 10480
rect 30300 9654 30328 11698
rect 30380 11688 30432 11694
rect 30380 11630 30432 11636
rect 30288 9648 30340 9654
rect 30288 9590 30340 9596
rect 30012 9512 30064 9518
rect 30300 9489 30328 9590
rect 30012 9454 30064 9460
rect 30286 9480 30342 9489
rect 30392 9450 30420 11630
rect 30484 9450 30512 12815
rect 30576 11257 30604 14894
rect 30760 14822 30788 17138
rect 31036 16590 31064 18294
rect 31024 16584 31076 16590
rect 31024 16526 31076 16532
rect 31036 16182 31064 16526
rect 31024 16176 31076 16182
rect 31024 16118 31076 16124
rect 30840 15428 30892 15434
rect 30840 15370 30892 15376
rect 30748 14816 30800 14822
rect 30748 14758 30800 14764
rect 30852 13394 30880 15370
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 30944 14278 30972 14350
rect 30932 14272 30984 14278
rect 30932 14214 30984 14220
rect 30840 13388 30892 13394
rect 30840 13330 30892 13336
rect 30656 13320 30708 13326
rect 30708 13280 30788 13308
rect 30656 13262 30708 13268
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30562 11248 30618 11257
rect 30562 11183 30618 11192
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30576 9518 30604 11086
rect 30668 9654 30696 12038
rect 30760 10713 30788 13280
rect 30746 10704 30802 10713
rect 30746 10639 30802 10648
rect 30748 10600 30800 10606
rect 30748 10542 30800 10548
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30286 9415 30342 9424
rect 30380 9444 30432 9450
rect 30380 9386 30432 9392
rect 30472 9444 30524 9450
rect 30472 9386 30524 9392
rect 29736 9036 29788 9042
rect 29736 8978 29788 8984
rect 29748 6866 29776 8978
rect 30012 8016 30064 8022
rect 30012 7958 30064 7964
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 30024 5642 30052 7958
rect 30012 5636 30064 5642
rect 30012 5578 30064 5584
rect 30576 3126 30604 9454
rect 30656 8356 30708 8362
rect 30656 8298 30708 8304
rect 30564 3120 30616 3126
rect 30564 3062 30616 3068
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30392 2514 30420 2790
rect 30380 2508 30432 2514
rect 30380 2450 30432 2456
rect 30196 2440 30248 2446
rect 30196 2382 30248 2388
rect 30208 800 30236 2382
rect 30668 2378 30696 8298
rect 30760 3398 30788 10542
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 30852 2650 30880 13330
rect 30944 10606 30972 14214
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 31036 12918 31064 13466
rect 31024 12912 31076 12918
rect 31024 12854 31076 12860
rect 31036 10810 31064 12854
rect 31116 12096 31168 12102
rect 31116 12038 31168 12044
rect 31128 11150 31156 12038
rect 31116 11144 31168 11150
rect 31116 11086 31168 11092
rect 31116 11008 31168 11014
rect 31116 10950 31168 10956
rect 31024 10804 31076 10810
rect 31024 10746 31076 10752
rect 30932 10600 30984 10606
rect 30932 10542 30984 10548
rect 31128 10538 31156 10950
rect 31208 10600 31260 10606
rect 31208 10542 31260 10548
rect 31116 10532 31168 10538
rect 31116 10474 31168 10480
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 30932 9988 30984 9994
rect 30932 9930 30984 9936
rect 30944 8430 30972 9930
rect 31036 9926 31064 10406
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 31220 9602 31248 10542
rect 31128 9586 31248 9602
rect 31116 9580 31248 9586
rect 31168 9574 31248 9580
rect 31116 9522 31168 9528
rect 30932 8424 30984 8430
rect 30932 8366 30984 8372
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30840 2644 30892 2650
rect 30840 2586 30892 2592
rect 30656 2372 30708 2378
rect 30656 2314 30708 2320
rect 30944 800 30972 3538
rect 31128 2922 31156 9522
rect 31312 4826 31340 25162
rect 31496 24818 31524 26522
rect 32140 26314 32168 27406
rect 32128 26308 32180 26314
rect 32128 26250 32180 26256
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 31852 25968 31904 25974
rect 31852 25910 31904 25916
rect 31864 24993 31892 25910
rect 31850 24984 31906 24993
rect 31850 24919 31906 24928
rect 31484 24812 31536 24818
rect 31484 24754 31536 24760
rect 31392 24132 31444 24138
rect 31392 24074 31444 24080
rect 31404 23798 31432 24074
rect 32048 23798 32076 25978
rect 32140 24138 32168 26250
rect 32128 24132 32180 24138
rect 32128 24074 32180 24080
rect 31392 23792 31444 23798
rect 31392 23734 31444 23740
rect 32036 23792 32088 23798
rect 32036 23734 32088 23740
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31680 21418 31708 21830
rect 31668 21412 31720 21418
rect 31668 21354 31720 21360
rect 31760 21004 31812 21010
rect 31760 20946 31812 20952
rect 31772 20602 31800 20946
rect 31760 20596 31812 20602
rect 31760 20538 31812 20544
rect 31772 19310 31800 20538
rect 31760 19304 31812 19310
rect 31760 19246 31812 19252
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31576 18352 31628 18358
rect 31576 18294 31628 18300
rect 31588 15706 31616 18294
rect 31576 15700 31628 15706
rect 31576 15642 31628 15648
rect 31680 15570 31708 18702
rect 32048 17746 32076 23734
rect 32232 22982 32260 27542
rect 32772 26920 32824 26926
rect 32772 26862 32824 26868
rect 32680 26852 32732 26858
rect 32680 26794 32732 26800
rect 32496 25492 32548 25498
rect 32496 25434 32548 25440
rect 32404 24608 32456 24614
rect 32324 24556 32404 24562
rect 32324 24550 32456 24556
rect 32324 24534 32444 24550
rect 32324 24138 32352 24534
rect 32312 24132 32364 24138
rect 32312 24074 32364 24080
rect 32404 23860 32456 23866
rect 32404 23802 32456 23808
rect 32220 22976 32272 22982
rect 32220 22918 32272 22924
rect 32220 19236 32272 19242
rect 32220 19178 32272 19184
rect 32128 19168 32180 19174
rect 32128 19110 32180 19116
rect 32140 18902 32168 19110
rect 32128 18896 32180 18902
rect 32128 18838 32180 18844
rect 32128 18080 32180 18086
rect 32128 18022 32180 18028
rect 32036 17740 32088 17746
rect 32036 17682 32088 17688
rect 32034 17640 32090 17649
rect 32034 17575 32090 17584
rect 31760 17332 31812 17338
rect 31760 17274 31812 17280
rect 31772 17082 31800 17274
rect 32048 17270 32076 17575
rect 32036 17264 32088 17270
rect 32036 17206 32088 17212
rect 32140 17202 32168 18022
rect 32128 17196 32180 17202
rect 32128 17138 32180 17144
rect 31772 17054 31984 17082
rect 31760 16992 31812 16998
rect 31760 16934 31812 16940
rect 31772 16250 31800 16934
rect 31956 16794 31984 17054
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 31944 16652 31996 16658
rect 31944 16594 31996 16600
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 31668 15564 31720 15570
rect 31668 15506 31720 15512
rect 31956 15094 31984 16594
rect 32140 16522 32168 17138
rect 32128 16516 32180 16522
rect 32128 16458 32180 16464
rect 32036 16040 32088 16046
rect 32036 15982 32088 15988
rect 31944 15088 31996 15094
rect 31944 15030 31996 15036
rect 31852 14952 31904 14958
rect 31852 14894 31904 14900
rect 31484 14612 31536 14618
rect 31484 14554 31536 14560
rect 31496 14482 31524 14554
rect 31484 14476 31536 14482
rect 31484 14418 31536 14424
rect 31496 12434 31524 14418
rect 31864 14346 31892 14894
rect 32048 14414 32076 15982
rect 32128 15020 32180 15026
rect 32128 14962 32180 14968
rect 32140 14618 32168 14962
rect 32128 14612 32180 14618
rect 32128 14554 32180 14560
rect 32036 14408 32088 14414
rect 32036 14350 32088 14356
rect 31852 14340 31904 14346
rect 31852 14282 31904 14288
rect 31576 14272 31628 14278
rect 31576 14214 31628 14220
rect 31588 12986 31616 14214
rect 32128 14068 32180 14074
rect 32128 14010 32180 14016
rect 31760 13320 31812 13326
rect 31680 13268 31760 13274
rect 31680 13262 31812 13268
rect 31680 13246 31800 13262
rect 31576 12980 31628 12986
rect 31576 12922 31628 12928
rect 31496 12406 31616 12434
rect 31390 11248 31446 11257
rect 31588 11218 31616 12406
rect 31680 12345 31708 13246
rect 31760 12640 31812 12646
rect 31760 12582 31812 12588
rect 31772 12434 31800 12582
rect 31852 12436 31904 12442
rect 31772 12406 31852 12434
rect 31852 12378 31904 12384
rect 31760 12368 31812 12374
rect 31666 12336 31722 12345
rect 31760 12310 31812 12316
rect 31666 12271 31722 12280
rect 31668 11892 31720 11898
rect 31668 11834 31720 11840
rect 31390 11183 31446 11192
rect 31576 11212 31628 11218
rect 31404 11150 31432 11183
rect 31576 11154 31628 11160
rect 31392 11144 31444 11150
rect 31588 11098 31616 11154
rect 31392 11086 31444 11092
rect 31496 11070 31616 11098
rect 31392 10804 31444 10810
rect 31392 10746 31444 10752
rect 31404 9994 31432 10746
rect 31392 9988 31444 9994
rect 31392 9930 31444 9936
rect 31404 8974 31432 9930
rect 31496 9722 31524 11070
rect 31576 11008 31628 11014
rect 31680 10996 31708 11834
rect 31772 11762 31800 12310
rect 31760 11756 31812 11762
rect 31760 11698 31812 11704
rect 31628 10968 31708 10996
rect 31576 10950 31628 10956
rect 31484 9716 31536 9722
rect 31484 9658 31536 9664
rect 31392 8968 31444 8974
rect 31392 8910 31444 8916
rect 31404 6730 31432 8910
rect 31484 8832 31536 8838
rect 31484 8774 31536 8780
rect 31496 7954 31524 8774
rect 31484 7948 31536 7954
rect 31484 7890 31536 7896
rect 31496 7002 31524 7890
rect 31484 6996 31536 7002
rect 31484 6938 31536 6944
rect 31392 6724 31444 6730
rect 31392 6666 31444 6672
rect 31404 6458 31432 6666
rect 31392 6452 31444 6458
rect 31392 6394 31444 6400
rect 31300 4820 31352 4826
rect 31300 4762 31352 4768
rect 31116 2916 31168 2922
rect 31116 2858 31168 2864
rect 31588 1834 31616 10950
rect 31668 9444 31720 9450
rect 31668 9386 31720 9392
rect 31680 8430 31708 9386
rect 31864 9042 31892 12378
rect 32140 11354 32168 14010
rect 32232 12306 32260 19178
rect 32416 18698 32444 23802
rect 32508 23610 32536 25434
rect 32692 24954 32720 26794
rect 32784 25362 32812 26862
rect 32772 25356 32824 25362
rect 32772 25298 32824 25304
rect 32680 24948 32732 24954
rect 32680 24890 32732 24896
rect 32588 24744 32640 24750
rect 32586 24712 32588 24721
rect 32640 24712 32642 24721
rect 32586 24647 32642 24656
rect 32784 24154 32812 25298
rect 32876 25158 32904 28154
rect 32950 27772 33258 27781
rect 32950 27770 32956 27772
rect 33012 27770 33036 27772
rect 33092 27770 33116 27772
rect 33172 27770 33196 27772
rect 33252 27770 33258 27772
rect 33012 27718 33014 27770
rect 33194 27718 33196 27770
rect 32950 27716 32956 27718
rect 33012 27716 33036 27718
rect 33092 27716 33116 27718
rect 33172 27716 33196 27718
rect 33252 27716 33258 27718
rect 32950 27707 33258 27716
rect 33232 27328 33284 27334
rect 33232 27270 33284 27276
rect 33244 26874 33272 27270
rect 33336 27130 33364 29514
rect 33416 28484 33468 28490
rect 33416 28426 33468 28432
rect 33324 27124 33376 27130
rect 33324 27066 33376 27072
rect 33244 26846 33364 26874
rect 32950 26684 33258 26693
rect 32950 26682 32956 26684
rect 33012 26682 33036 26684
rect 33092 26682 33116 26684
rect 33172 26682 33196 26684
rect 33252 26682 33258 26684
rect 33012 26630 33014 26682
rect 33194 26630 33196 26682
rect 32950 26628 32956 26630
rect 33012 26628 33036 26630
rect 33092 26628 33116 26630
rect 33172 26628 33196 26630
rect 33252 26628 33258 26630
rect 32950 26619 33258 26628
rect 33048 25968 33100 25974
rect 33048 25910 33100 25916
rect 33060 25809 33088 25910
rect 33046 25800 33102 25809
rect 33046 25735 33102 25744
rect 32950 25596 33258 25605
rect 32950 25594 32956 25596
rect 33012 25594 33036 25596
rect 33092 25594 33116 25596
rect 33172 25594 33196 25596
rect 33252 25594 33258 25596
rect 33012 25542 33014 25594
rect 33194 25542 33196 25594
rect 32950 25540 32956 25542
rect 33012 25540 33036 25542
rect 33092 25540 33116 25542
rect 33172 25540 33196 25542
rect 33252 25540 33258 25542
rect 32950 25531 33258 25540
rect 33336 25362 33364 26846
rect 32956 25356 33008 25362
rect 32956 25298 33008 25304
rect 33324 25356 33376 25362
rect 33324 25298 33376 25304
rect 32864 25152 32916 25158
rect 32864 25094 32916 25100
rect 32600 24126 32812 24154
rect 32600 24070 32628 24126
rect 32588 24064 32640 24070
rect 32588 24006 32640 24012
rect 32876 23866 32904 25094
rect 32968 24750 32996 25298
rect 33428 24954 33456 28426
rect 33520 28150 33548 29650
rect 33600 29504 33652 29510
rect 33600 29446 33652 29452
rect 33508 28144 33560 28150
rect 33508 28086 33560 28092
rect 33508 28008 33560 28014
rect 33508 27950 33560 27956
rect 33520 26450 33548 27950
rect 33612 27402 33640 29446
rect 33600 27396 33652 27402
rect 33600 27338 33652 27344
rect 33600 27124 33652 27130
rect 33600 27066 33652 27072
rect 33508 26444 33560 26450
rect 33508 26386 33560 26392
rect 33612 26330 33640 27066
rect 33520 26302 33640 26330
rect 33416 24948 33468 24954
rect 33416 24890 33468 24896
rect 33520 24800 33548 26302
rect 33600 25696 33652 25702
rect 33600 25638 33652 25644
rect 33336 24772 33548 24800
rect 32956 24744 33008 24750
rect 32956 24686 33008 24692
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32956 24064 33008 24070
rect 32956 24006 33008 24012
rect 32864 23860 32916 23866
rect 32864 23802 32916 23808
rect 32508 23582 32812 23610
rect 32680 23520 32732 23526
rect 32680 23462 32732 23468
rect 32496 22976 32548 22982
rect 32496 22918 32548 22924
rect 32508 19446 32536 22918
rect 32692 21146 32720 23462
rect 32784 21690 32812 23582
rect 32968 23526 32996 24006
rect 32956 23520 33008 23526
rect 32956 23462 33008 23468
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32864 22976 32916 22982
rect 32864 22918 32916 22924
rect 32876 22098 32904 22918
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33336 22166 33364 24772
rect 33612 24750 33640 25638
rect 33600 24744 33652 24750
rect 33600 24686 33652 24692
rect 33876 24744 33928 24750
rect 33876 24686 33928 24692
rect 33508 24676 33560 24682
rect 33508 24618 33560 24624
rect 33520 24342 33548 24618
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33612 24274 33640 24686
rect 33600 24268 33652 24274
rect 33600 24210 33652 24216
rect 33416 23180 33468 23186
rect 33416 23122 33468 23128
rect 33428 22778 33456 23122
rect 33508 23044 33560 23050
rect 33508 22986 33560 22992
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33324 22160 33376 22166
rect 33324 22102 33376 22108
rect 32864 22092 32916 22098
rect 32864 22034 32916 22040
rect 32772 21684 32824 21690
rect 32772 21626 32824 21632
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32680 21140 32732 21146
rect 32680 21082 32732 21088
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32588 19848 32640 19854
rect 32588 19790 32640 19796
rect 32496 19440 32548 19446
rect 32496 19382 32548 19388
rect 32600 18834 32628 19790
rect 32772 19372 32824 19378
rect 32772 19314 32824 19320
rect 32588 18828 32640 18834
rect 32588 18770 32640 18776
rect 32404 18692 32456 18698
rect 32404 18634 32456 18640
rect 32312 18420 32364 18426
rect 32312 18362 32364 18368
rect 32324 14890 32352 18362
rect 32312 14884 32364 14890
rect 32312 14826 32364 14832
rect 32416 14822 32444 18634
rect 32588 18080 32640 18086
rect 32588 18022 32640 18028
rect 32404 14816 32456 14822
rect 32404 14758 32456 14764
rect 32404 13728 32456 13734
rect 32404 13670 32456 13676
rect 32312 13524 32364 13530
rect 32312 13466 32364 13472
rect 32324 12918 32352 13466
rect 32416 13394 32444 13670
rect 32404 13388 32456 13394
rect 32404 13330 32456 13336
rect 32312 12912 32364 12918
rect 32312 12854 32364 12860
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32220 12300 32272 12306
rect 32220 12242 32272 12248
rect 32324 11370 32352 12582
rect 32128 11348 32180 11354
rect 32128 11290 32180 11296
rect 32232 11342 32352 11370
rect 31944 11076 31996 11082
rect 31944 11018 31996 11024
rect 31956 9110 31984 11018
rect 32128 11008 32180 11014
rect 32128 10950 32180 10956
rect 32140 10674 32168 10950
rect 32128 10668 32180 10674
rect 32128 10610 32180 10616
rect 32232 9994 32260 11342
rect 32312 11280 32364 11286
rect 32312 11222 32364 11228
rect 32324 11150 32352 11222
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32416 10266 32444 13330
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32508 12306 32536 12378
rect 32496 12300 32548 12306
rect 32496 12242 32548 12248
rect 32600 11642 32628 18022
rect 32680 13864 32732 13870
rect 32680 13806 32732 13812
rect 32508 11614 32628 11642
rect 32508 11558 32536 11614
rect 32496 11552 32548 11558
rect 32496 11494 32548 11500
rect 32404 10260 32456 10266
rect 32404 10202 32456 10208
rect 32312 10124 32364 10130
rect 32312 10066 32364 10072
rect 32220 9988 32272 9994
rect 32220 9930 32272 9936
rect 31944 9104 31996 9110
rect 31944 9046 31996 9052
rect 32126 9072 32182 9081
rect 31852 9036 31904 9042
rect 32126 9007 32128 9016
rect 31852 8978 31904 8984
rect 32180 9007 32182 9016
rect 32128 8978 32180 8984
rect 31668 8424 31720 8430
rect 31668 8366 31720 8372
rect 31668 8016 31720 8022
rect 31668 7958 31720 7964
rect 31680 7886 31708 7958
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 32140 3738 32168 8978
rect 32324 8634 32352 10066
rect 32312 8628 32364 8634
rect 32312 8570 32364 8576
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32324 8090 32352 8434
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32312 6860 32364 6866
rect 32312 6802 32364 6808
rect 32220 6724 32272 6730
rect 32220 6666 32272 6672
rect 32232 5778 32260 6666
rect 32324 6322 32352 6802
rect 32312 6316 32364 6322
rect 32312 6258 32364 6264
rect 32220 5772 32272 5778
rect 32220 5714 32272 5720
rect 32416 5710 32444 7822
rect 32508 7478 32536 11494
rect 32588 11280 32640 11286
rect 32588 11222 32640 11228
rect 32600 11121 32628 11222
rect 32586 11112 32642 11121
rect 32586 11047 32588 11056
rect 32640 11047 32642 11056
rect 32588 11018 32640 11024
rect 32692 10266 32720 13806
rect 32784 12986 32812 19314
rect 32864 19168 32916 19174
rect 32864 19110 32916 19116
rect 32876 18834 32904 19110
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32864 18828 32916 18834
rect 32864 18770 32916 18776
rect 32876 18698 32904 18770
rect 32864 18692 32916 18698
rect 32864 18634 32916 18640
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 33428 17762 33456 22578
rect 33520 22506 33548 22986
rect 33508 22500 33560 22506
rect 33508 22442 33560 22448
rect 33508 22160 33560 22166
rect 33508 22102 33560 22108
rect 33520 19514 33548 22102
rect 33612 21010 33640 24210
rect 33784 24064 33836 24070
rect 33784 24006 33836 24012
rect 33600 21004 33652 21010
rect 33600 20946 33652 20952
rect 33796 20942 33824 24006
rect 33888 23662 33916 24686
rect 33876 23656 33928 23662
rect 33928 23604 34008 23610
rect 33876 23598 34008 23604
rect 33888 23582 34008 23598
rect 33980 22574 34008 23582
rect 34072 22982 34100 35866
rect 34716 31754 34744 52838
rect 37950 52252 38258 52261
rect 37950 52250 37956 52252
rect 38012 52250 38036 52252
rect 38092 52250 38116 52252
rect 38172 52250 38196 52252
rect 38252 52250 38258 52252
rect 38012 52198 38014 52250
rect 38194 52198 38196 52250
rect 37950 52196 37956 52198
rect 38012 52196 38036 52198
rect 38092 52196 38116 52198
rect 38172 52196 38196 52198
rect 38252 52196 38258 52198
rect 37950 52187 38258 52196
rect 37950 51164 38258 51173
rect 37950 51162 37956 51164
rect 38012 51162 38036 51164
rect 38092 51162 38116 51164
rect 38172 51162 38196 51164
rect 38252 51162 38258 51164
rect 38012 51110 38014 51162
rect 38194 51110 38196 51162
rect 37950 51108 37956 51110
rect 38012 51108 38036 51110
rect 38092 51108 38116 51110
rect 38172 51108 38196 51110
rect 38252 51108 38258 51110
rect 37950 51099 38258 51108
rect 35716 50720 35768 50726
rect 35716 50662 35768 50668
rect 34980 43648 35032 43654
rect 34980 43590 35032 43596
rect 34716 31726 34836 31754
rect 34336 31680 34388 31686
rect 34336 31622 34388 31628
rect 34348 31346 34376 31622
rect 34336 31340 34388 31346
rect 34336 31282 34388 31288
rect 34348 28966 34376 31282
rect 34704 30048 34756 30054
rect 34704 29990 34756 29996
rect 34520 29776 34572 29782
rect 34520 29718 34572 29724
rect 34532 29306 34560 29718
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34520 29300 34572 29306
rect 34520 29242 34572 29248
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34532 29073 34560 29106
rect 34518 29064 34574 29073
rect 34518 28999 34574 29008
rect 34336 28960 34388 28966
rect 34336 28902 34388 28908
rect 34152 26444 34204 26450
rect 34152 26386 34204 26392
rect 34164 25362 34192 26386
rect 34152 25356 34204 25362
rect 34152 25298 34204 25304
rect 34060 22976 34112 22982
rect 34060 22918 34112 22924
rect 33968 22568 34020 22574
rect 33968 22510 34020 22516
rect 34072 22094 34100 22918
rect 34072 22066 34284 22094
rect 33784 20936 33836 20942
rect 33784 20878 33836 20884
rect 34152 19780 34204 19786
rect 34152 19722 34204 19728
rect 33508 19508 33560 19514
rect 33508 19450 33560 19456
rect 33968 19440 34020 19446
rect 33968 19382 34020 19388
rect 33876 19236 33928 19242
rect 33876 19178 33928 19184
rect 33336 17734 33456 17762
rect 33336 17610 33364 17734
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33324 17604 33376 17610
rect 33324 17546 33376 17552
rect 33428 17338 33456 17614
rect 33416 17332 33468 17338
rect 33416 17274 33468 17280
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33324 16584 33376 16590
rect 32876 16532 33324 16538
rect 32876 16526 33376 16532
rect 32876 16510 33364 16526
rect 32876 16454 32904 16510
rect 32864 16448 32916 16454
rect 32864 16390 32916 16396
rect 32956 16448 33008 16454
rect 32956 16390 33008 16396
rect 32968 16046 32996 16390
rect 32956 16040 33008 16046
rect 32956 15982 33008 15988
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32864 15156 32916 15162
rect 32864 15098 32916 15104
rect 32876 13938 32904 15098
rect 33336 15094 33364 16510
rect 33888 16454 33916 19178
rect 33980 17241 34008 19382
rect 34164 18698 34192 19722
rect 34152 18692 34204 18698
rect 34152 18634 34204 18640
rect 34152 17808 34204 17814
rect 34152 17750 34204 17756
rect 34060 17604 34112 17610
rect 34060 17546 34112 17552
rect 33966 17232 34022 17241
rect 33966 17167 34022 17176
rect 33980 16726 34008 17167
rect 33968 16720 34020 16726
rect 33968 16662 34020 16668
rect 33876 16448 33928 16454
rect 33876 16390 33928 16396
rect 33508 15428 33560 15434
rect 33508 15370 33560 15376
rect 33324 15088 33376 15094
rect 33324 15030 33376 15036
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 33336 14074 33364 15030
rect 33324 14068 33376 14074
rect 33324 14010 33376 14016
rect 33416 14000 33468 14006
rect 33416 13942 33468 13948
rect 32864 13932 32916 13938
rect 32864 13874 32916 13880
rect 32864 13796 32916 13802
rect 32864 13738 32916 13744
rect 32876 13394 32904 13738
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32864 13388 32916 13394
rect 32864 13330 32916 13336
rect 33428 13326 33456 13942
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 32772 12980 32824 12986
rect 32772 12922 32824 12928
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 33520 12442 33548 15370
rect 33692 15360 33744 15366
rect 33692 15302 33744 15308
rect 33704 15178 33732 15302
rect 33612 15150 33732 15178
rect 33508 12436 33560 12442
rect 33508 12378 33560 12384
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32772 11212 32824 11218
rect 32772 11154 32824 11160
rect 32784 10606 32812 11154
rect 32772 10600 32824 10606
rect 32772 10542 32824 10548
rect 33416 10600 33468 10606
rect 33416 10542 33468 10548
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32784 10130 32812 10542
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33324 10260 33376 10266
rect 33324 10202 33376 10208
rect 32772 10124 32824 10130
rect 32772 10066 32824 10072
rect 33336 9926 33364 10202
rect 33232 9920 33284 9926
rect 33232 9862 33284 9868
rect 33324 9920 33376 9926
rect 33324 9862 33376 9868
rect 33244 9722 33272 9862
rect 32588 9716 32640 9722
rect 32588 9658 32640 9664
rect 33232 9716 33284 9722
rect 33232 9658 33284 9664
rect 32600 9058 32628 9658
rect 33230 9616 33286 9625
rect 33230 9551 33286 9560
rect 33244 9518 33272 9551
rect 33232 9512 33284 9518
rect 33232 9454 33284 9460
rect 32772 9376 32824 9382
rect 32772 9318 32824 9324
rect 32600 9042 32720 9058
rect 32784 9042 32812 9318
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32588 9036 32720 9042
rect 32640 9030 32720 9036
rect 32588 8978 32640 8984
rect 32586 8936 32642 8945
rect 32586 8871 32642 8880
rect 32600 8838 32628 8871
rect 32588 8832 32640 8838
rect 32588 8774 32640 8780
rect 32692 8498 32720 9030
rect 32772 9036 32824 9042
rect 32772 8978 32824 8984
rect 33336 8922 33364 9862
rect 33244 8894 33364 8922
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 33152 8344 33180 8774
rect 33244 8650 33272 8894
rect 33428 8838 33456 10542
rect 33520 9081 33548 11630
rect 33506 9072 33562 9081
rect 33506 9007 33562 9016
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33244 8622 33548 8650
rect 33152 8316 33364 8344
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32588 7948 32640 7954
rect 32588 7890 32640 7896
rect 32496 7472 32548 7478
rect 32496 7414 32548 7420
rect 32600 6662 32628 7890
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32588 6656 32640 6662
rect 32588 6598 32640 6604
rect 32600 6390 32628 6598
rect 32588 6384 32640 6390
rect 32588 6326 32640 6332
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32404 5704 32456 5710
rect 32404 5646 32456 5652
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 32128 3732 32180 3738
rect 32128 3674 32180 3680
rect 33336 3670 33364 8316
rect 33416 7744 33468 7750
rect 33416 7686 33468 7692
rect 33428 5914 33456 7686
rect 33416 5908 33468 5914
rect 33416 5850 33468 5856
rect 33324 3664 33376 3670
rect 33324 3606 33376 3612
rect 33520 3194 33548 8622
rect 33508 3188 33560 3194
rect 33508 3130 33560 3136
rect 31668 2984 31720 2990
rect 31668 2926 31720 2932
rect 31576 1828 31628 1834
rect 31576 1770 31628 1776
rect 31680 800 31708 2926
rect 32404 2916 32456 2922
rect 32404 2858 32456 2864
rect 32416 800 32444 2858
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33612 2582 33640 15150
rect 33784 13184 33836 13190
rect 33784 13126 33836 13132
rect 33692 12640 33744 12646
rect 33692 12582 33744 12588
rect 33704 12170 33732 12582
rect 33692 12164 33744 12170
rect 33692 12106 33744 12112
rect 33600 2576 33652 2582
rect 33600 2518 33652 2524
rect 33796 2446 33824 13126
rect 33888 12714 33916 16390
rect 34072 14958 34100 17546
rect 34060 14952 34112 14958
rect 34060 14894 34112 14900
rect 34072 12850 34100 14894
rect 34060 12844 34112 12850
rect 34060 12786 34112 12792
rect 33968 12776 34020 12782
rect 34164 12764 34192 17750
rect 34256 15502 34284 22066
rect 34348 19446 34376 28902
rect 34624 28200 34652 29582
rect 34532 28172 34652 28200
rect 34532 26994 34560 28172
rect 34612 28076 34664 28082
rect 34612 28018 34664 28024
rect 34624 27674 34652 28018
rect 34716 27878 34744 29990
rect 34808 29238 34836 31726
rect 34992 31278 35020 43590
rect 35164 31340 35216 31346
rect 35164 31282 35216 31288
rect 34980 31272 35032 31278
rect 34980 31214 35032 31220
rect 35176 30054 35204 31282
rect 35624 31272 35676 31278
rect 35624 31214 35676 31220
rect 35440 30660 35492 30666
rect 35440 30602 35492 30608
rect 35164 30048 35216 30054
rect 35164 29990 35216 29996
rect 35072 29776 35124 29782
rect 35072 29718 35124 29724
rect 34796 29232 34848 29238
rect 34796 29174 34848 29180
rect 34888 29232 34940 29238
rect 34888 29174 34940 29180
rect 34900 28506 34928 29174
rect 34808 28478 34928 28506
rect 34704 27872 34756 27878
rect 34704 27814 34756 27820
rect 34612 27668 34664 27674
rect 34612 27610 34664 27616
rect 34520 26988 34572 26994
rect 34520 26930 34572 26936
rect 34624 26024 34652 27610
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 34532 25996 34652 26024
rect 34428 25968 34480 25974
rect 34532 25956 34560 25996
rect 34480 25928 34560 25956
rect 34428 25910 34480 25916
rect 34440 24886 34468 25910
rect 34520 25356 34572 25362
rect 34520 25298 34572 25304
rect 34428 24880 34480 24886
rect 34428 24822 34480 24828
rect 34440 24206 34468 24822
rect 34428 24200 34480 24206
rect 34428 24142 34480 24148
rect 34440 23798 34468 24142
rect 34428 23792 34480 23798
rect 34428 23734 34480 23740
rect 34440 21622 34468 23734
rect 34532 22234 34560 25298
rect 34612 24948 34664 24954
rect 34612 24890 34664 24896
rect 34520 22228 34572 22234
rect 34520 22170 34572 22176
rect 34624 22094 34652 24890
rect 34716 23798 34744 26930
rect 34704 23792 34756 23798
rect 34704 23734 34756 23740
rect 34808 23730 34836 28478
rect 34888 28416 34940 28422
rect 34888 28358 34940 28364
rect 34900 27334 34928 28358
rect 34980 27872 35032 27878
rect 34980 27814 35032 27820
rect 34992 27538 35020 27814
rect 34980 27532 35032 27538
rect 34980 27474 35032 27480
rect 34888 27328 34940 27334
rect 34888 27270 34940 27276
rect 34992 25838 35020 27474
rect 35084 26450 35112 29718
rect 35256 29300 35308 29306
rect 35256 29242 35308 29248
rect 35164 29164 35216 29170
rect 35164 29106 35216 29112
rect 35176 26926 35204 29106
rect 35268 27130 35296 29242
rect 35348 28416 35400 28422
rect 35348 28358 35400 28364
rect 35360 27946 35388 28358
rect 35452 28150 35480 30602
rect 35636 30190 35664 31214
rect 35624 30184 35676 30190
rect 35624 30126 35676 30132
rect 35636 29850 35664 30126
rect 35624 29844 35676 29850
rect 35624 29786 35676 29792
rect 35532 29708 35584 29714
rect 35532 29650 35584 29656
rect 35544 28626 35572 29650
rect 35728 29073 35756 50662
rect 37950 50076 38258 50085
rect 37950 50074 37956 50076
rect 38012 50074 38036 50076
rect 38092 50074 38116 50076
rect 38172 50074 38196 50076
rect 38252 50074 38258 50076
rect 38012 50022 38014 50074
rect 38194 50022 38196 50074
rect 37950 50020 37956 50022
rect 38012 50020 38036 50022
rect 38092 50020 38116 50022
rect 38172 50020 38196 50022
rect 38252 50020 38258 50022
rect 37950 50011 38258 50020
rect 37950 48988 38258 48997
rect 37950 48986 37956 48988
rect 38012 48986 38036 48988
rect 38092 48986 38116 48988
rect 38172 48986 38196 48988
rect 38252 48986 38258 48988
rect 38012 48934 38014 48986
rect 38194 48934 38196 48986
rect 37950 48932 37956 48934
rect 38012 48932 38036 48934
rect 38092 48932 38116 48934
rect 38172 48932 38196 48934
rect 38252 48932 38258 48934
rect 37950 48923 38258 48932
rect 37950 47900 38258 47909
rect 37950 47898 37956 47900
rect 38012 47898 38036 47900
rect 38092 47898 38116 47900
rect 38172 47898 38196 47900
rect 38252 47898 38258 47900
rect 38012 47846 38014 47898
rect 38194 47846 38196 47898
rect 37950 47844 37956 47846
rect 38012 47844 38036 47846
rect 38092 47844 38116 47846
rect 38172 47844 38196 47846
rect 38252 47844 38258 47846
rect 37950 47835 38258 47844
rect 37950 46812 38258 46821
rect 37950 46810 37956 46812
rect 38012 46810 38036 46812
rect 38092 46810 38116 46812
rect 38172 46810 38196 46812
rect 38252 46810 38258 46812
rect 38012 46758 38014 46810
rect 38194 46758 38196 46810
rect 37950 46756 37956 46758
rect 38012 46756 38036 46758
rect 38092 46756 38116 46758
rect 38172 46756 38196 46758
rect 38252 46756 38258 46758
rect 37950 46747 38258 46756
rect 37950 45724 38258 45733
rect 37950 45722 37956 45724
rect 38012 45722 38036 45724
rect 38092 45722 38116 45724
rect 38172 45722 38196 45724
rect 38252 45722 38258 45724
rect 38012 45670 38014 45722
rect 38194 45670 38196 45722
rect 37950 45668 37956 45670
rect 38012 45668 38036 45670
rect 38092 45668 38116 45670
rect 38172 45668 38196 45670
rect 38252 45668 38258 45670
rect 37950 45659 38258 45668
rect 37950 44636 38258 44645
rect 37950 44634 37956 44636
rect 38012 44634 38036 44636
rect 38092 44634 38116 44636
rect 38172 44634 38196 44636
rect 38252 44634 38258 44636
rect 38012 44582 38014 44634
rect 38194 44582 38196 44634
rect 37950 44580 37956 44582
rect 38012 44580 38036 44582
rect 38092 44580 38116 44582
rect 38172 44580 38196 44582
rect 38252 44580 38258 44582
rect 37950 44571 38258 44580
rect 37950 43548 38258 43557
rect 37950 43546 37956 43548
rect 38012 43546 38036 43548
rect 38092 43546 38116 43548
rect 38172 43546 38196 43548
rect 38252 43546 38258 43548
rect 38012 43494 38014 43546
rect 38194 43494 38196 43546
rect 37950 43492 37956 43494
rect 38012 43492 38036 43494
rect 38092 43492 38116 43494
rect 38172 43492 38196 43494
rect 38252 43492 38258 43494
rect 37950 43483 38258 43492
rect 37950 42460 38258 42469
rect 37950 42458 37956 42460
rect 38012 42458 38036 42460
rect 38092 42458 38116 42460
rect 38172 42458 38196 42460
rect 38252 42458 38258 42460
rect 38012 42406 38014 42458
rect 38194 42406 38196 42458
rect 37950 42404 37956 42406
rect 38012 42404 38036 42406
rect 38092 42404 38116 42406
rect 38172 42404 38196 42406
rect 38252 42404 38258 42406
rect 37950 42395 38258 42404
rect 36820 41472 36872 41478
rect 36820 41414 36872 41420
rect 35900 30320 35952 30326
rect 35900 30262 35952 30268
rect 35808 30048 35860 30054
rect 35808 29990 35860 29996
rect 35820 29238 35848 29990
rect 35912 29714 35940 30262
rect 35992 30252 36044 30258
rect 35992 30194 36044 30200
rect 35900 29708 35952 29714
rect 35900 29650 35952 29656
rect 35808 29232 35860 29238
rect 35808 29174 35860 29180
rect 35714 29064 35770 29073
rect 35714 28999 35770 29008
rect 35808 29028 35860 29034
rect 35808 28970 35860 28976
rect 35716 28960 35768 28966
rect 35716 28902 35768 28908
rect 35532 28620 35584 28626
rect 35532 28562 35584 28568
rect 35440 28144 35492 28150
rect 35440 28086 35492 28092
rect 35348 27940 35400 27946
rect 35348 27882 35400 27888
rect 35624 27940 35676 27946
rect 35624 27882 35676 27888
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 35256 27124 35308 27130
rect 35308 27084 35388 27112
rect 35256 27066 35308 27072
rect 35164 26920 35216 26926
rect 35164 26862 35216 26868
rect 35072 26444 35124 26450
rect 35072 26386 35124 26392
rect 34980 25832 35032 25838
rect 34980 25774 35032 25780
rect 35084 25158 35112 26386
rect 35072 25152 35124 25158
rect 35072 25094 35124 25100
rect 34888 24676 34940 24682
rect 34888 24618 34940 24624
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 34796 23588 34848 23594
rect 34796 23530 34848 23536
rect 34532 22066 34652 22094
rect 34428 21616 34480 21622
rect 34428 21558 34480 21564
rect 34532 21570 34560 22066
rect 34532 21542 34652 21570
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 34428 20800 34480 20806
rect 34428 20742 34480 20748
rect 34336 19440 34388 19446
rect 34336 19382 34388 19388
rect 34440 19378 34468 20742
rect 34532 20534 34560 21422
rect 34520 20528 34572 20534
rect 34520 20470 34572 20476
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34428 18760 34480 18766
rect 34428 18702 34480 18708
rect 34336 18624 34388 18630
rect 34336 18566 34388 18572
rect 34348 18222 34376 18566
rect 34336 18216 34388 18222
rect 34336 18158 34388 18164
rect 34348 16658 34376 18158
rect 34336 16652 34388 16658
rect 34336 16594 34388 16600
rect 34244 15496 34296 15502
rect 34244 15438 34296 15444
rect 34164 12736 34284 12764
rect 33968 12718 34020 12724
rect 33876 12708 33928 12714
rect 33876 12650 33928 12656
rect 33876 12164 33928 12170
rect 33876 12106 33928 12112
rect 33888 11898 33916 12106
rect 33876 11892 33928 11898
rect 33876 11834 33928 11840
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 33152 800 33180 2246
rect 33888 800 33916 4014
rect 33980 3058 34008 12718
rect 34060 11076 34112 11082
rect 34060 11018 34112 11024
rect 34072 8498 34100 11018
rect 34256 10985 34284 12736
rect 34242 10976 34298 10985
rect 34242 10911 34298 10920
rect 34152 10600 34204 10606
rect 34152 10542 34204 10548
rect 34164 10266 34192 10542
rect 34152 10260 34204 10266
rect 34152 10202 34204 10208
rect 34060 8492 34112 8498
rect 34060 8434 34112 8440
rect 34072 6866 34100 8434
rect 34152 7336 34204 7342
rect 34152 7278 34204 7284
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 34164 6458 34192 7278
rect 34256 6798 34284 10911
rect 34440 8974 34468 18702
rect 34532 17746 34560 20470
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34532 16250 34560 17682
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34532 15570 34560 16186
rect 34520 15564 34572 15570
rect 34520 15506 34572 15512
rect 34532 15162 34560 15506
rect 34520 15156 34572 15162
rect 34520 15098 34572 15104
rect 34520 14000 34572 14006
rect 34520 13942 34572 13948
rect 34532 11286 34560 13942
rect 34520 11280 34572 11286
rect 34520 11222 34572 11228
rect 34624 9994 34652 21542
rect 34704 20392 34756 20398
rect 34704 20334 34756 20340
rect 34716 19718 34744 20334
rect 34808 20058 34836 23530
rect 34900 21468 34928 24618
rect 34980 23792 35032 23798
rect 34980 23734 35032 23740
rect 34992 23322 35020 23734
rect 34980 23316 35032 23322
rect 34980 23258 35032 23264
rect 34992 21962 35020 23258
rect 34980 21956 35032 21962
rect 34980 21898 35032 21904
rect 35072 21480 35124 21486
rect 34900 21440 35072 21468
rect 35072 21422 35124 21428
rect 34796 20052 34848 20058
rect 34796 19994 34848 20000
rect 34704 19712 34756 19718
rect 34704 19654 34756 19660
rect 34808 16250 34836 19994
rect 35072 19848 35124 19854
rect 35072 19790 35124 19796
rect 35084 18970 35112 19790
rect 35176 19514 35204 26862
rect 35256 26376 35308 26382
rect 35254 26344 35256 26353
rect 35308 26344 35310 26353
rect 35254 26279 35310 26288
rect 35360 26228 35388 27084
rect 35440 26920 35492 26926
rect 35440 26862 35492 26868
rect 35452 26450 35480 26862
rect 35440 26444 35492 26450
rect 35440 26386 35492 26392
rect 35268 26200 35388 26228
rect 35268 24206 35296 26200
rect 35348 25696 35400 25702
rect 35348 25638 35400 25644
rect 35256 24200 35308 24206
rect 35256 24142 35308 24148
rect 35268 23798 35296 24142
rect 35256 23792 35308 23798
rect 35256 23734 35308 23740
rect 35256 23520 35308 23526
rect 35256 23462 35308 23468
rect 35164 19508 35216 19514
rect 35164 19450 35216 19456
rect 35072 18964 35124 18970
rect 35072 18906 35124 18912
rect 34888 17536 34940 17542
rect 34888 17478 34940 17484
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 34808 16130 34836 16186
rect 34716 16102 34836 16130
rect 34716 14346 34744 16102
rect 34796 16040 34848 16046
rect 34796 15982 34848 15988
rect 34808 14482 34836 15982
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 34704 14340 34756 14346
rect 34704 14282 34756 14288
rect 34808 14074 34836 14418
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34900 13258 34928 17478
rect 35072 16584 35124 16590
rect 35072 16526 35124 16532
rect 35084 16182 35112 16526
rect 35072 16176 35124 16182
rect 35072 16118 35124 16124
rect 34980 15088 35032 15094
rect 34980 15030 35032 15036
rect 34992 13954 35020 15030
rect 35072 14544 35124 14550
rect 35072 14486 35124 14492
rect 35084 14074 35112 14486
rect 35072 14068 35124 14074
rect 35072 14010 35124 14016
rect 34992 13926 35112 13954
rect 34888 13252 34940 13258
rect 34888 13194 34940 13200
rect 34704 12708 34756 12714
rect 34704 12650 34756 12656
rect 34980 12708 35032 12714
rect 34980 12650 35032 12656
rect 34716 11830 34744 12650
rect 34796 12640 34848 12646
rect 34796 12582 34848 12588
rect 34808 11898 34836 12582
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 34704 11824 34756 11830
rect 34704 11766 34756 11772
rect 34704 10532 34756 10538
rect 34704 10474 34756 10480
rect 34612 9988 34664 9994
rect 34612 9930 34664 9936
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34428 8968 34480 8974
rect 34428 8910 34480 8916
rect 34532 8634 34560 9454
rect 34428 8628 34480 8634
rect 34428 8570 34480 8576
rect 34520 8628 34572 8634
rect 34520 8570 34572 8576
rect 34440 8537 34468 8570
rect 34426 8528 34482 8537
rect 34426 8463 34482 8472
rect 34532 7562 34560 8570
rect 34624 8022 34652 9930
rect 34716 9178 34744 10474
rect 34796 10464 34848 10470
rect 34848 10412 34928 10418
rect 34796 10406 34928 10412
rect 34808 10390 34928 10406
rect 34900 10062 34928 10390
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 34796 9648 34848 9654
rect 34796 9590 34848 9596
rect 34808 9353 34836 9590
rect 34794 9344 34850 9353
rect 34794 9279 34850 9288
rect 34704 9172 34756 9178
rect 34704 9114 34756 9120
rect 34900 8974 34928 9998
rect 34888 8968 34940 8974
rect 34888 8910 34940 8916
rect 34612 8016 34664 8022
rect 34612 7958 34664 7964
rect 34532 7534 34652 7562
rect 34900 7546 34928 8910
rect 34624 7342 34652 7534
rect 34888 7540 34940 7546
rect 34888 7482 34940 7488
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 34612 7336 34664 7342
rect 34612 7278 34664 7284
rect 34428 7200 34480 7206
rect 34428 7142 34480 7148
rect 34244 6792 34296 6798
rect 34244 6734 34296 6740
rect 34152 6452 34204 6458
rect 34152 6394 34204 6400
rect 34440 3534 34468 7142
rect 34716 6730 34744 7414
rect 34704 6724 34756 6730
rect 34704 6666 34756 6672
rect 34716 6390 34744 6666
rect 34704 6384 34756 6390
rect 34704 6326 34756 6332
rect 34612 3596 34664 3602
rect 34612 3538 34664 3544
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 33968 3052 34020 3058
rect 33968 2994 34020 3000
rect 34624 800 34652 3538
rect 34992 3058 35020 12650
rect 35084 10538 35112 13926
rect 35176 13326 35204 19450
rect 35268 18834 35296 23462
rect 35360 22778 35388 25638
rect 35452 24614 35480 26386
rect 35544 26042 35572 27270
rect 35532 26036 35584 26042
rect 35532 25978 35584 25984
rect 35636 24721 35664 27882
rect 35728 27538 35756 28902
rect 35716 27532 35768 27538
rect 35716 27474 35768 27480
rect 35820 26042 35848 28970
rect 35912 27470 35940 29650
rect 36004 29617 36032 30194
rect 35990 29608 36046 29617
rect 35990 29543 36046 29552
rect 35900 27464 35952 27470
rect 35900 27406 35952 27412
rect 35808 26036 35860 26042
rect 35808 25978 35860 25984
rect 35912 25226 35940 27406
rect 36004 27334 36032 29543
rect 36176 28552 36228 28558
rect 36176 28494 36228 28500
rect 36188 28014 36216 28494
rect 36176 28008 36228 28014
rect 36176 27950 36228 27956
rect 35992 27328 36044 27334
rect 35990 27296 35992 27305
rect 36044 27296 36046 27305
rect 35990 27231 36046 27240
rect 36188 26926 36216 27950
rect 36176 26920 36228 26926
rect 36176 26862 36228 26868
rect 36188 25770 36216 26862
rect 36268 26512 36320 26518
rect 36268 26454 36320 26460
rect 36176 25764 36228 25770
rect 36176 25706 36228 25712
rect 35900 25220 35952 25226
rect 35900 25162 35952 25168
rect 35912 24954 35940 25162
rect 35900 24948 35952 24954
rect 35900 24890 35952 24896
rect 35622 24712 35678 24721
rect 35622 24647 35678 24656
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 35636 24342 35664 24647
rect 35624 24336 35676 24342
rect 35624 24278 35676 24284
rect 35636 23662 35664 24278
rect 35440 23656 35492 23662
rect 35440 23598 35492 23604
rect 35624 23656 35676 23662
rect 35624 23598 35676 23604
rect 35452 23254 35480 23598
rect 35532 23520 35584 23526
rect 35532 23462 35584 23468
rect 35440 23248 35492 23254
rect 35440 23190 35492 23196
rect 35348 22772 35400 22778
rect 35348 22714 35400 22720
rect 35452 22098 35480 23190
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 35348 21616 35400 21622
rect 35348 21558 35400 21564
rect 35360 20874 35388 21558
rect 35440 21480 35492 21486
rect 35440 21422 35492 21428
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 35360 20466 35388 20810
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 35360 19786 35388 20402
rect 35452 20262 35480 21422
rect 35440 20256 35492 20262
rect 35440 20198 35492 20204
rect 35348 19780 35400 19786
rect 35348 19722 35400 19728
rect 35348 19304 35400 19310
rect 35348 19246 35400 19252
rect 35256 18828 35308 18834
rect 35256 18770 35308 18776
rect 35256 18624 35308 18630
rect 35256 18566 35308 18572
rect 35268 18426 35296 18566
rect 35256 18420 35308 18426
rect 35256 18362 35308 18368
rect 35360 15094 35388 19246
rect 35452 16522 35480 20198
rect 35544 18426 35572 23462
rect 35900 22160 35952 22166
rect 35900 22102 35952 22108
rect 35624 19712 35676 19718
rect 35624 19654 35676 19660
rect 35636 18970 35664 19654
rect 35624 18964 35676 18970
rect 35624 18906 35676 18912
rect 35716 18624 35768 18630
rect 35716 18566 35768 18572
rect 35532 18420 35584 18426
rect 35532 18362 35584 18368
rect 35440 16516 35492 16522
rect 35440 16458 35492 16464
rect 35532 16448 35584 16454
rect 35532 16390 35584 16396
rect 35348 15088 35400 15094
rect 35348 15030 35400 15036
rect 35348 14612 35400 14618
rect 35348 14554 35400 14560
rect 35256 14000 35308 14006
rect 35256 13942 35308 13948
rect 35268 13870 35296 13942
rect 35256 13864 35308 13870
rect 35256 13806 35308 13812
rect 35164 13320 35216 13326
rect 35164 13262 35216 13268
rect 35176 12306 35204 13262
rect 35360 12918 35388 14554
rect 35348 12912 35400 12918
rect 35348 12854 35400 12860
rect 35164 12300 35216 12306
rect 35164 12242 35216 12248
rect 35256 11620 35308 11626
rect 35256 11562 35308 11568
rect 35164 11212 35216 11218
rect 35164 11154 35216 11160
rect 35072 10532 35124 10538
rect 35072 10474 35124 10480
rect 35072 9988 35124 9994
rect 35072 9930 35124 9936
rect 35084 9586 35112 9930
rect 35072 9580 35124 9586
rect 35072 9522 35124 9528
rect 35176 8906 35204 11154
rect 35268 11082 35296 11562
rect 35346 11112 35402 11121
rect 35256 11076 35308 11082
rect 35346 11047 35348 11056
rect 35256 11018 35308 11024
rect 35400 11047 35402 11056
rect 35348 11018 35400 11024
rect 35360 10282 35388 11018
rect 35268 10254 35388 10282
rect 35268 9625 35296 10254
rect 35348 10192 35400 10198
rect 35544 10146 35572 16390
rect 35624 15564 35676 15570
rect 35624 15506 35676 15512
rect 35636 15094 35664 15506
rect 35624 15088 35676 15094
rect 35624 15030 35676 15036
rect 35624 14272 35676 14278
rect 35624 14214 35676 14220
rect 35636 13462 35664 14214
rect 35624 13456 35676 13462
rect 35624 13398 35676 13404
rect 35728 10742 35756 18566
rect 35808 16788 35860 16794
rect 35808 16730 35860 16736
rect 35820 13326 35848 16730
rect 35912 15570 35940 22102
rect 35992 20460 36044 20466
rect 35992 20402 36044 20408
rect 36004 15978 36032 20402
rect 36176 19780 36228 19786
rect 36176 19722 36228 19728
rect 36188 17610 36216 19722
rect 36280 18290 36308 26454
rect 36636 25152 36688 25158
rect 36636 25094 36688 25100
rect 36728 25152 36780 25158
rect 36728 25094 36780 25100
rect 36544 24948 36596 24954
rect 36544 24890 36596 24896
rect 36556 22778 36584 24890
rect 36648 24818 36676 25094
rect 36740 24954 36768 25094
rect 36728 24948 36780 24954
rect 36728 24890 36780 24896
rect 36636 24812 36688 24818
rect 36688 24772 36768 24800
rect 36636 24754 36688 24760
rect 36636 24608 36688 24614
rect 36636 24550 36688 24556
rect 36544 22772 36596 22778
rect 36544 22714 36596 22720
rect 36452 21344 36504 21350
rect 36452 21286 36504 21292
rect 36544 21344 36596 21350
rect 36544 21286 36596 21292
rect 36464 21078 36492 21286
rect 36452 21072 36504 21078
rect 36452 21014 36504 21020
rect 36556 21010 36584 21286
rect 36544 21004 36596 21010
rect 36544 20946 36596 20952
rect 36556 20482 36584 20946
rect 36648 20602 36676 24550
rect 36740 22710 36768 24772
rect 36728 22704 36780 22710
rect 36728 22646 36780 22652
rect 36636 20596 36688 20602
rect 36636 20538 36688 20544
rect 36556 20454 36676 20482
rect 36648 20398 36676 20454
rect 36636 20392 36688 20398
rect 36636 20334 36688 20340
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 36268 18284 36320 18290
rect 36268 18226 36320 18232
rect 36176 17604 36228 17610
rect 36176 17546 36228 17552
rect 36188 16182 36216 17546
rect 36176 16176 36228 16182
rect 36176 16118 36228 16124
rect 35992 15972 36044 15978
rect 35992 15914 36044 15920
rect 36188 15688 36216 16118
rect 36188 15660 36308 15688
rect 35900 15564 35952 15570
rect 35952 15524 36216 15552
rect 35900 15506 35952 15512
rect 35900 14340 35952 14346
rect 35900 14282 35952 14288
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35912 11150 35940 14282
rect 35992 13252 36044 13258
rect 35992 13194 36044 13200
rect 35900 11144 35952 11150
rect 35900 11086 35952 11092
rect 35716 10736 35768 10742
rect 35716 10678 35768 10684
rect 35400 10140 35572 10146
rect 35348 10134 35572 10140
rect 35360 10118 35572 10134
rect 35254 9616 35310 9625
rect 35254 9551 35310 9560
rect 35164 8900 35216 8906
rect 35164 8842 35216 8848
rect 35176 8090 35204 8842
rect 35544 8786 35572 10118
rect 35716 9988 35768 9994
rect 35716 9930 35768 9936
rect 35728 9178 35756 9930
rect 35716 9172 35768 9178
rect 35716 9114 35768 9120
rect 35544 8758 35664 8786
rect 35256 8628 35308 8634
rect 35256 8570 35308 8576
rect 35164 8084 35216 8090
rect 35164 8026 35216 8032
rect 35268 7478 35296 8570
rect 35348 8356 35400 8362
rect 35348 8298 35400 8304
rect 35256 7472 35308 7478
rect 35256 7414 35308 7420
rect 35360 4146 35388 8298
rect 35532 7812 35584 7818
rect 35532 7754 35584 7760
rect 35544 7410 35572 7754
rect 35532 7404 35584 7410
rect 35532 7346 35584 7352
rect 35636 6730 35664 8758
rect 35728 8634 35756 9114
rect 35716 8628 35768 8634
rect 35716 8570 35768 8576
rect 35808 8424 35860 8430
rect 35808 8366 35860 8372
rect 35820 7886 35848 8366
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35808 7880 35860 7886
rect 35808 7822 35860 7828
rect 35728 7478 35756 7822
rect 35820 7546 35848 7822
rect 35808 7540 35860 7546
rect 35808 7482 35860 7488
rect 35716 7472 35768 7478
rect 35716 7414 35768 7420
rect 35820 6866 35848 7482
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 35624 6724 35676 6730
rect 35624 6666 35676 6672
rect 35348 4140 35400 4146
rect 35348 4082 35400 4088
rect 36004 3398 36032 13194
rect 36188 12442 36216 15524
rect 36280 15450 36308 15660
rect 36280 15434 36400 15450
rect 36280 15428 36412 15434
rect 36280 15422 36360 15428
rect 36360 15370 36412 15376
rect 36556 15094 36584 19654
rect 36728 16652 36780 16658
rect 36728 16594 36780 16600
rect 36544 15088 36596 15094
rect 36544 15030 36596 15036
rect 36268 15020 36320 15026
rect 36268 14962 36320 14968
rect 36280 14346 36308 14962
rect 36452 14816 36504 14822
rect 36452 14758 36504 14764
rect 36268 14340 36320 14346
rect 36268 14282 36320 14288
rect 36268 13388 36320 13394
rect 36268 13330 36320 13336
rect 36176 12436 36228 12442
rect 36176 12378 36228 12384
rect 36280 12306 36308 13330
rect 36268 12300 36320 12306
rect 36268 12242 36320 12248
rect 36266 11792 36322 11801
rect 36266 11727 36268 11736
rect 36320 11727 36322 11736
rect 36268 11698 36320 11704
rect 36084 10736 36136 10742
rect 36082 10704 36084 10713
rect 36136 10704 36138 10713
rect 36082 10639 36138 10648
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 36268 9376 36320 9382
rect 36268 9318 36320 9324
rect 36176 8968 36228 8974
rect 36176 8910 36228 8916
rect 36188 8566 36216 8910
rect 36176 8560 36228 8566
rect 36176 8502 36228 8508
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 34980 3052 35032 3058
rect 34980 2994 35032 3000
rect 35348 2508 35400 2514
rect 35348 2450 35400 2456
rect 35360 800 35388 2450
rect 36096 800 36124 3538
rect 36280 2446 36308 9318
rect 36372 8498 36400 10406
rect 36464 9602 36492 14758
rect 36740 12434 36768 16594
rect 36832 14385 36860 41414
rect 37950 41372 38258 41381
rect 37950 41370 37956 41372
rect 38012 41370 38036 41372
rect 38092 41370 38116 41372
rect 38172 41370 38196 41372
rect 38252 41370 38258 41372
rect 38012 41318 38014 41370
rect 38194 41318 38196 41370
rect 37950 41316 37956 41318
rect 38012 41316 38036 41318
rect 38092 41316 38116 41318
rect 38172 41316 38196 41318
rect 38252 41316 38258 41318
rect 37950 41307 38258 41316
rect 37950 40284 38258 40293
rect 37950 40282 37956 40284
rect 38012 40282 38036 40284
rect 38092 40282 38116 40284
rect 38172 40282 38196 40284
rect 38252 40282 38258 40284
rect 38012 40230 38014 40282
rect 38194 40230 38196 40282
rect 37950 40228 37956 40230
rect 38012 40228 38036 40230
rect 38092 40228 38116 40230
rect 38172 40228 38196 40230
rect 38252 40228 38258 40230
rect 37950 40219 38258 40228
rect 37950 39196 38258 39205
rect 37950 39194 37956 39196
rect 38012 39194 38036 39196
rect 38092 39194 38116 39196
rect 38172 39194 38196 39196
rect 38252 39194 38258 39196
rect 38012 39142 38014 39194
rect 38194 39142 38196 39194
rect 37950 39140 37956 39142
rect 38012 39140 38036 39142
rect 38092 39140 38116 39142
rect 38172 39140 38196 39142
rect 38252 39140 38258 39142
rect 37950 39131 38258 39140
rect 37950 38108 38258 38117
rect 37950 38106 37956 38108
rect 38012 38106 38036 38108
rect 38092 38106 38116 38108
rect 38172 38106 38196 38108
rect 38252 38106 38258 38108
rect 38012 38054 38014 38106
rect 38194 38054 38196 38106
rect 37950 38052 37956 38054
rect 38012 38052 38036 38054
rect 38092 38052 38116 38054
rect 38172 38052 38196 38054
rect 38252 38052 38258 38054
rect 37950 38043 38258 38052
rect 37950 37020 38258 37029
rect 37950 37018 37956 37020
rect 38012 37018 38036 37020
rect 38092 37018 38116 37020
rect 38172 37018 38196 37020
rect 38252 37018 38258 37020
rect 38012 36966 38014 37018
rect 38194 36966 38196 37018
rect 37950 36964 37956 36966
rect 38012 36964 38036 36966
rect 38092 36964 38116 36966
rect 38172 36964 38196 36966
rect 38252 36964 38258 36966
rect 37950 36955 38258 36964
rect 37950 35932 38258 35941
rect 37950 35930 37956 35932
rect 38012 35930 38036 35932
rect 38092 35930 38116 35932
rect 38172 35930 38196 35932
rect 38252 35930 38258 35932
rect 38012 35878 38014 35930
rect 38194 35878 38196 35930
rect 37950 35876 37956 35878
rect 38012 35876 38036 35878
rect 38092 35876 38116 35878
rect 38172 35876 38196 35878
rect 38252 35876 38258 35878
rect 37950 35867 38258 35876
rect 37950 34844 38258 34853
rect 37950 34842 37956 34844
rect 38012 34842 38036 34844
rect 38092 34842 38116 34844
rect 38172 34842 38196 34844
rect 38252 34842 38258 34844
rect 38012 34790 38014 34842
rect 38194 34790 38196 34842
rect 37950 34788 37956 34790
rect 38012 34788 38036 34790
rect 38092 34788 38116 34790
rect 38172 34788 38196 34790
rect 38252 34788 38258 34790
rect 37950 34779 38258 34788
rect 38384 34128 38436 34134
rect 38384 34070 38436 34076
rect 37950 33756 38258 33765
rect 37950 33754 37956 33756
rect 38012 33754 38036 33756
rect 38092 33754 38116 33756
rect 38172 33754 38196 33756
rect 38252 33754 38258 33756
rect 38012 33702 38014 33754
rect 38194 33702 38196 33754
rect 37950 33700 37956 33702
rect 38012 33700 38036 33702
rect 38092 33700 38116 33702
rect 38172 33700 38196 33702
rect 38252 33700 38258 33702
rect 37950 33691 38258 33700
rect 37950 32668 38258 32677
rect 37950 32666 37956 32668
rect 38012 32666 38036 32668
rect 38092 32666 38116 32668
rect 38172 32666 38196 32668
rect 38252 32666 38258 32668
rect 38012 32614 38014 32666
rect 38194 32614 38196 32666
rect 37950 32612 37956 32614
rect 38012 32612 38036 32614
rect 38092 32612 38116 32614
rect 38172 32612 38196 32614
rect 38252 32612 38258 32614
rect 37950 32603 38258 32612
rect 38292 32224 38344 32230
rect 38292 32166 38344 32172
rect 37950 31580 38258 31589
rect 37950 31578 37956 31580
rect 38012 31578 38036 31580
rect 38092 31578 38116 31580
rect 38172 31578 38196 31580
rect 38252 31578 38258 31580
rect 38012 31526 38014 31578
rect 38194 31526 38196 31578
rect 37950 31524 37956 31526
rect 38012 31524 38036 31526
rect 38092 31524 38116 31526
rect 38172 31524 38196 31526
rect 38252 31524 38258 31526
rect 37950 31515 38258 31524
rect 38304 31278 38332 32166
rect 38292 31272 38344 31278
rect 38292 31214 38344 31220
rect 37464 30660 37516 30666
rect 37464 30602 37516 30608
rect 37476 30258 37504 30602
rect 38292 30592 38344 30598
rect 38292 30534 38344 30540
rect 37950 30492 38258 30501
rect 37950 30490 37956 30492
rect 38012 30490 38036 30492
rect 38092 30490 38116 30492
rect 38172 30490 38196 30492
rect 38252 30490 38258 30492
rect 38012 30438 38014 30490
rect 38194 30438 38196 30490
rect 37950 30436 37956 30438
rect 38012 30436 38036 30438
rect 38092 30436 38116 30438
rect 38172 30436 38196 30438
rect 38252 30436 38258 30438
rect 37950 30427 38258 30436
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 37476 29170 37504 30194
rect 37950 29404 38258 29413
rect 37950 29402 37956 29404
rect 38012 29402 38036 29404
rect 38092 29402 38116 29404
rect 38172 29402 38196 29404
rect 38252 29402 38258 29404
rect 38012 29350 38014 29402
rect 38194 29350 38196 29402
rect 37950 29348 37956 29350
rect 38012 29348 38036 29350
rect 38092 29348 38116 29350
rect 38172 29348 38196 29350
rect 38252 29348 38258 29350
rect 37950 29339 38258 29348
rect 37464 29164 37516 29170
rect 37464 29106 37516 29112
rect 37950 28316 38258 28325
rect 37950 28314 37956 28316
rect 38012 28314 38036 28316
rect 38092 28314 38116 28316
rect 38172 28314 38196 28316
rect 38252 28314 38258 28316
rect 38012 28262 38014 28314
rect 38194 28262 38196 28314
rect 37950 28260 37956 28262
rect 38012 28260 38036 28262
rect 38092 28260 38116 28262
rect 38172 28260 38196 28262
rect 38252 28260 38258 28262
rect 37950 28251 38258 28260
rect 37648 27872 37700 27878
rect 37648 27814 37700 27820
rect 37372 25152 37424 25158
rect 37372 25094 37424 25100
rect 37004 23656 37056 23662
rect 37004 23598 37056 23604
rect 36912 23588 36964 23594
rect 36912 23530 36964 23536
rect 36924 16522 36952 23530
rect 37016 21146 37044 23598
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 37188 21888 37240 21894
rect 37188 21830 37240 21836
rect 37004 21140 37056 21146
rect 37004 21082 37056 21088
rect 37016 19174 37044 21082
rect 37096 20868 37148 20874
rect 37096 20810 37148 20816
rect 37004 19168 37056 19174
rect 37004 19110 37056 19116
rect 37108 17882 37136 20810
rect 37096 17876 37148 17882
rect 37096 17818 37148 17824
rect 37004 17672 37056 17678
rect 37004 17614 37056 17620
rect 37016 17270 37044 17614
rect 37004 17264 37056 17270
rect 37004 17206 37056 17212
rect 37200 16590 37228 21830
rect 37188 16584 37240 16590
rect 37188 16526 37240 16532
rect 36912 16516 36964 16522
rect 36912 16458 36964 16464
rect 37292 15502 37320 21898
rect 37384 17746 37412 25094
rect 37556 23656 37608 23662
rect 37556 23598 37608 23604
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 37372 17740 37424 17746
rect 37372 17682 37424 17688
rect 37476 17338 37504 18158
rect 37464 17332 37516 17338
rect 37464 17274 37516 17280
rect 37372 16516 37424 16522
rect 37372 16458 37424 16464
rect 37280 15496 37332 15502
rect 37280 15438 37332 15444
rect 37280 15020 37332 15026
rect 37280 14962 37332 14968
rect 36818 14376 36874 14385
rect 36818 14311 36874 14320
rect 36832 12918 36860 14311
rect 37292 13682 37320 14962
rect 37384 14006 37412 16458
rect 37568 16114 37596 23598
rect 37660 18834 37688 27814
rect 37950 27228 38258 27237
rect 37950 27226 37956 27228
rect 38012 27226 38036 27228
rect 38092 27226 38116 27228
rect 38172 27226 38196 27228
rect 38252 27226 38258 27228
rect 38012 27174 38014 27226
rect 38194 27174 38196 27226
rect 37950 27172 37956 27174
rect 38012 27172 38036 27174
rect 38092 27172 38116 27174
rect 38172 27172 38196 27174
rect 38252 27172 38258 27174
rect 37950 27163 38258 27172
rect 38304 26450 38332 30534
rect 38396 28082 38424 34070
rect 38476 32360 38528 32366
rect 38476 32302 38528 32308
rect 38488 31414 38516 32302
rect 38476 31408 38528 31414
rect 38476 31350 38528 31356
rect 38488 30326 38516 31350
rect 38568 31272 38620 31278
rect 38568 31214 38620 31220
rect 38476 30320 38528 30326
rect 38476 30262 38528 30268
rect 38476 28960 38528 28966
rect 38476 28902 38528 28908
rect 38488 28626 38516 28902
rect 38476 28620 38528 28626
rect 38476 28562 38528 28568
rect 38384 28076 38436 28082
rect 38384 28018 38436 28024
rect 38384 27872 38436 27878
rect 38384 27814 38436 27820
rect 38292 26444 38344 26450
rect 38292 26386 38344 26392
rect 37950 26140 38258 26149
rect 37950 26138 37956 26140
rect 38012 26138 38036 26140
rect 38092 26138 38116 26140
rect 38172 26138 38196 26140
rect 38252 26138 38258 26140
rect 38012 26086 38014 26138
rect 38194 26086 38196 26138
rect 37950 26084 37956 26086
rect 38012 26084 38036 26086
rect 38092 26084 38116 26086
rect 38172 26084 38196 26086
rect 38252 26084 38258 26086
rect 37950 26075 38258 26084
rect 37740 25696 37792 25702
rect 37740 25638 37792 25644
rect 37752 25294 37780 25638
rect 37740 25288 37792 25294
rect 37740 25230 37792 25236
rect 37950 25052 38258 25061
rect 37950 25050 37956 25052
rect 38012 25050 38036 25052
rect 38092 25050 38116 25052
rect 38172 25050 38196 25052
rect 38252 25050 38258 25052
rect 38012 24998 38014 25050
rect 38194 24998 38196 25050
rect 37950 24996 37956 24998
rect 38012 24996 38036 24998
rect 38092 24996 38116 24998
rect 38172 24996 38196 24998
rect 38252 24996 38258 24998
rect 37950 24987 38258 24996
rect 37740 24812 37792 24818
rect 37740 24754 37792 24760
rect 37752 24138 37780 24754
rect 38396 24698 38424 27814
rect 38488 25362 38516 28562
rect 38580 28014 38608 31214
rect 39040 30054 39068 53926
rect 41236 46368 41288 46374
rect 41236 46310 41288 46316
rect 41248 34066 41276 46310
rect 41420 43784 41472 43790
rect 41420 43726 41472 43732
rect 41236 34060 41288 34066
rect 41236 34002 41288 34008
rect 39672 33992 39724 33998
rect 39672 33934 39724 33940
rect 39684 31142 39712 33934
rect 40960 33856 41012 33862
rect 40960 33798 41012 33804
rect 41236 33856 41288 33862
rect 41236 33798 41288 33804
rect 40590 33416 40646 33425
rect 40590 33351 40646 33360
rect 40224 33312 40276 33318
rect 40224 33254 40276 33260
rect 40132 32496 40184 32502
rect 40132 32438 40184 32444
rect 40040 31816 40092 31822
rect 40040 31758 40092 31764
rect 40052 31346 40080 31758
rect 40144 31414 40172 32438
rect 40132 31408 40184 31414
rect 40132 31350 40184 31356
rect 40040 31340 40092 31346
rect 40040 31282 40092 31288
rect 39672 31136 39724 31142
rect 39672 31078 39724 31084
rect 39120 30388 39172 30394
rect 39120 30330 39172 30336
rect 39028 30048 39080 30054
rect 39028 29990 39080 29996
rect 39132 29238 39160 30330
rect 39684 30190 39712 31078
rect 39948 30796 40000 30802
rect 39948 30738 40000 30744
rect 39672 30184 39724 30190
rect 39672 30126 39724 30132
rect 39488 30116 39540 30122
rect 39488 30058 39540 30064
rect 39120 29232 39172 29238
rect 39120 29174 39172 29180
rect 39132 28994 39160 29174
rect 39040 28966 39160 28994
rect 39040 28558 39068 28966
rect 39028 28552 39080 28558
rect 39028 28494 39080 28500
rect 39396 28552 39448 28558
rect 39396 28494 39448 28500
rect 38844 28484 38896 28490
rect 38844 28426 38896 28432
rect 38568 28008 38620 28014
rect 38568 27950 38620 27956
rect 38856 26450 38884 28426
rect 39040 28150 39068 28494
rect 39408 28218 39436 28494
rect 39500 28422 39528 30058
rect 39764 30048 39816 30054
rect 39764 29990 39816 29996
rect 39488 28416 39540 28422
rect 39488 28358 39540 28364
rect 39396 28212 39448 28218
rect 39396 28154 39448 28160
rect 39028 28144 39080 28150
rect 39028 28086 39080 28092
rect 39040 27062 39068 28086
rect 39500 27130 39528 28358
rect 39776 27538 39804 29990
rect 39960 29102 39988 30738
rect 40144 30326 40172 31350
rect 40132 30320 40184 30326
rect 40132 30262 40184 30268
rect 40040 29232 40092 29238
rect 40040 29174 40092 29180
rect 39948 29096 40000 29102
rect 39948 29038 40000 29044
rect 39948 28960 40000 28966
rect 39948 28902 40000 28908
rect 39960 28490 39988 28902
rect 40052 28558 40080 29174
rect 40040 28552 40092 28558
rect 40040 28494 40092 28500
rect 39948 28484 40000 28490
rect 39948 28426 40000 28432
rect 40052 28064 40080 28494
rect 40236 28218 40264 33254
rect 40316 31884 40368 31890
rect 40316 31826 40368 31832
rect 40328 31142 40356 31826
rect 40316 31136 40368 31142
rect 40316 31078 40368 31084
rect 40224 28212 40276 28218
rect 40224 28154 40276 28160
rect 40052 28036 40172 28064
rect 39856 27872 39908 27878
rect 39856 27814 39908 27820
rect 39764 27532 39816 27538
rect 39764 27474 39816 27480
rect 39488 27124 39540 27130
rect 39488 27066 39540 27072
rect 39028 27056 39080 27062
rect 39028 26998 39080 27004
rect 38844 26444 38896 26450
rect 38844 26386 38896 26392
rect 39040 26246 39068 26998
rect 39776 26314 39804 27474
rect 39764 26308 39816 26314
rect 39764 26250 39816 26256
rect 39028 26240 39080 26246
rect 39028 26182 39080 26188
rect 38568 25424 38620 25430
rect 38568 25366 38620 25372
rect 38476 25356 38528 25362
rect 38476 25298 38528 25304
rect 38580 24818 38608 25366
rect 38568 24812 38620 24818
rect 38568 24754 38620 24760
rect 38304 24670 38424 24698
rect 37832 24608 37884 24614
rect 37832 24550 37884 24556
rect 37740 24132 37792 24138
rect 37740 24074 37792 24080
rect 37740 23724 37792 23730
rect 37740 23666 37792 23672
rect 37752 23118 37780 23666
rect 37844 23633 37872 24550
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 37830 23624 37886 23633
rect 37830 23559 37886 23568
rect 37740 23112 37792 23118
rect 37740 23054 37792 23060
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37740 22500 37792 22506
rect 37740 22442 37792 22448
rect 37648 18828 37700 18834
rect 37648 18770 37700 18776
rect 37752 18442 37780 22442
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37832 21548 37884 21554
rect 37832 21490 37884 21496
rect 37844 21146 37872 21490
rect 37832 21140 37884 21146
rect 37832 21082 37884 21088
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 38304 18766 38332 24670
rect 38384 24608 38436 24614
rect 38384 24550 38436 24556
rect 39212 24608 39264 24614
rect 39212 24550 39264 24556
rect 38396 24342 38424 24550
rect 38384 24336 38436 24342
rect 38384 24278 38436 24284
rect 38660 24200 38712 24206
rect 38660 24142 38712 24148
rect 38672 23798 38700 24142
rect 38660 23792 38712 23798
rect 38660 23734 38712 23740
rect 39028 23724 39080 23730
rect 39028 23666 39080 23672
rect 38844 23520 38896 23526
rect 38844 23462 38896 23468
rect 38384 23180 38436 23186
rect 38384 23122 38436 23128
rect 38396 21690 38424 23122
rect 38476 22432 38528 22438
rect 38476 22374 38528 22380
rect 38384 21684 38436 21690
rect 38384 21626 38436 21632
rect 38292 18760 38344 18766
rect 38292 18702 38344 18708
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37660 18414 37780 18442
rect 38384 18420 38436 18426
rect 37660 18358 37688 18414
rect 38384 18362 38436 18368
rect 37648 18352 37700 18358
rect 37648 18294 37700 18300
rect 37660 17218 37688 18294
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37660 17190 37872 17218
rect 37556 16108 37608 16114
rect 37556 16050 37608 16056
rect 37556 15904 37608 15910
rect 37556 15846 37608 15852
rect 37464 15428 37516 15434
rect 37464 15370 37516 15376
rect 37372 14000 37424 14006
rect 37372 13942 37424 13948
rect 37108 13654 37320 13682
rect 37108 13530 37136 13654
rect 37096 13524 37148 13530
rect 37096 13466 37148 13472
rect 37188 13524 37240 13530
rect 37188 13466 37240 13472
rect 36820 12912 36872 12918
rect 36820 12854 36872 12860
rect 37200 12442 37228 13466
rect 37280 13252 37332 13258
rect 37280 13194 37332 13200
rect 37188 12436 37240 12442
rect 36740 12406 36860 12434
rect 36636 12164 36688 12170
rect 36636 12106 36688 12112
rect 36648 10266 36676 12106
rect 36832 11830 36860 12406
rect 37188 12378 37240 12384
rect 37292 12170 37320 13194
rect 37476 12434 37504 15370
rect 37384 12406 37504 12434
rect 37280 12164 37332 12170
rect 37280 12106 37332 12112
rect 36820 11824 36872 11830
rect 36820 11766 36872 11772
rect 36636 10260 36688 10266
rect 36636 10202 36688 10208
rect 36464 9574 36676 9602
rect 36452 9512 36504 9518
rect 36556 9489 36584 9574
rect 36452 9454 36504 9460
rect 36542 9480 36598 9489
rect 36464 8634 36492 9454
rect 36542 9415 36598 9424
rect 36452 8628 36504 8634
rect 36452 8570 36504 8576
rect 36360 8492 36412 8498
rect 36360 8434 36412 8440
rect 36464 7002 36492 8570
rect 36452 6996 36504 7002
rect 36452 6938 36504 6944
rect 36360 6792 36412 6798
rect 36360 6734 36412 6740
rect 36372 2446 36400 6734
rect 36648 5302 36676 9574
rect 36728 9512 36780 9518
rect 36728 9454 36780 9460
rect 36740 8566 36768 9454
rect 36728 8560 36780 8566
rect 36728 8502 36780 8508
rect 36832 5642 36860 11766
rect 37004 11076 37056 11082
rect 37004 11018 37056 11024
rect 37016 10606 37044 11018
rect 37004 10600 37056 10606
rect 37004 10542 37056 10548
rect 37016 10130 37044 10542
rect 37292 10146 37320 12106
rect 37004 10124 37056 10130
rect 37004 10066 37056 10072
rect 37200 10118 37320 10146
rect 37016 9586 37044 10066
rect 37200 10062 37228 10118
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 37004 9580 37056 9586
rect 37004 9522 37056 9528
rect 37004 8968 37056 8974
rect 37200 8922 37228 9998
rect 37384 9353 37412 12406
rect 37568 11014 37596 15846
rect 37660 13734 37688 17190
rect 37844 17134 37872 17190
rect 37740 17128 37792 17134
rect 37740 17070 37792 17076
rect 37832 17128 37884 17134
rect 37832 17070 37884 17076
rect 37752 15706 37780 17070
rect 37832 16720 37884 16726
rect 37832 16662 37884 16668
rect 37740 15700 37792 15706
rect 37740 15642 37792 15648
rect 37844 14056 37872 16662
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 38292 15904 38344 15910
rect 38292 15846 38344 15852
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 37924 14068 37976 14074
rect 37844 14028 37924 14056
rect 37924 14010 37976 14016
rect 37648 13728 37700 13734
rect 37648 13670 37700 13676
rect 37740 13184 37792 13190
rect 37740 13126 37792 13132
rect 37648 12640 37700 12646
rect 37648 12582 37700 12588
rect 37556 11008 37608 11014
rect 37556 10950 37608 10956
rect 37464 9376 37516 9382
rect 37370 9344 37426 9353
rect 37464 9318 37516 9324
rect 37370 9279 37426 9288
rect 37280 9104 37332 9110
rect 37280 9046 37332 9052
rect 37056 8916 37228 8922
rect 37004 8910 37228 8916
rect 37016 8894 37228 8910
rect 37200 8566 37228 8894
rect 37292 8838 37320 9046
rect 37280 8832 37332 8838
rect 37280 8774 37332 8780
rect 37188 8560 37240 8566
rect 37188 8502 37240 8508
rect 37200 7886 37228 8502
rect 37188 7880 37240 7886
rect 37188 7822 37240 7828
rect 37200 6730 37228 7822
rect 37188 6724 37240 6730
rect 37188 6666 37240 6672
rect 37200 6322 37228 6666
rect 37188 6316 37240 6322
rect 37188 6258 37240 6264
rect 37384 5710 37412 9279
rect 37476 8906 37504 9318
rect 37464 8900 37516 8906
rect 37464 8842 37516 8848
rect 37568 6390 37596 10950
rect 37556 6384 37608 6390
rect 37556 6326 37608 6332
rect 37372 5704 37424 5710
rect 37372 5646 37424 5652
rect 36820 5636 36872 5642
rect 36820 5578 36872 5584
rect 36636 5296 36688 5302
rect 36636 5238 36688 5244
rect 37660 5030 37688 12582
rect 37752 12442 37780 13126
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37740 12436 37792 12442
rect 37740 12378 37792 12384
rect 37752 11762 37780 12378
rect 38304 12209 38332 15846
rect 38290 12200 38346 12209
rect 37832 12164 37884 12170
rect 38290 12135 38346 12144
rect 37832 12106 37884 12112
rect 37844 11898 37872 12106
rect 38292 12096 38344 12102
rect 38292 12038 38344 12044
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 37832 11892 37884 11898
rect 37832 11834 37884 11840
rect 38304 11830 38332 12038
rect 38292 11824 38344 11830
rect 38292 11766 38344 11772
rect 37740 11756 37792 11762
rect 37740 11698 37792 11704
rect 37924 11688 37976 11694
rect 37924 11630 37976 11636
rect 38290 11656 38346 11665
rect 37936 11286 37964 11630
rect 38290 11591 38346 11600
rect 37924 11280 37976 11286
rect 38304 11257 38332 11591
rect 37924 11222 37976 11228
rect 38290 11248 38346 11257
rect 38290 11183 38346 11192
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 37844 10470 37872 11086
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 37832 10464 37884 10470
rect 37832 10406 37884 10412
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 37740 7948 37792 7954
rect 37740 7890 37792 7896
rect 37752 6866 37780 7890
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 37740 6860 37792 6866
rect 37740 6802 37792 6808
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 38304 6390 38332 11183
rect 38396 9654 38424 18362
rect 38488 16658 38516 22374
rect 38856 21622 38884 23462
rect 39040 21690 39068 23666
rect 39120 23248 39172 23254
rect 39120 23190 39172 23196
rect 39132 22030 39160 23190
rect 39224 22098 39252 24550
rect 39868 23798 39896 27814
rect 39948 26920 40000 26926
rect 39948 26862 40000 26868
rect 39960 25770 39988 26862
rect 40144 26382 40172 28036
rect 40328 28014 40356 31078
rect 40604 30734 40632 33351
rect 40592 30728 40644 30734
rect 40592 30670 40644 30676
rect 40592 30048 40644 30054
rect 40592 29990 40644 29996
rect 40408 28076 40460 28082
rect 40408 28018 40460 28024
rect 40316 28008 40368 28014
rect 40316 27950 40368 27956
rect 40420 27674 40448 28018
rect 40408 27668 40460 27674
rect 40408 27610 40460 27616
rect 40500 27328 40552 27334
rect 40500 27270 40552 27276
rect 40132 26376 40184 26382
rect 40132 26318 40184 26324
rect 40144 26042 40172 26318
rect 40132 26036 40184 26042
rect 40132 25978 40184 25984
rect 39948 25764 40000 25770
rect 39948 25706 40000 25712
rect 39856 23792 39908 23798
rect 39856 23734 39908 23740
rect 39960 23662 39988 25706
rect 40408 25696 40460 25702
rect 40408 25638 40460 25644
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 39948 23656 40000 23662
rect 39948 23598 40000 23604
rect 40052 23594 40080 25230
rect 40316 24200 40368 24206
rect 40316 24142 40368 24148
rect 40328 23798 40356 24142
rect 40316 23792 40368 23798
rect 40316 23734 40368 23740
rect 40420 23610 40448 25638
rect 40512 23798 40540 27270
rect 40604 25226 40632 29990
rect 40972 27402 41000 33798
rect 41248 33425 41276 33798
rect 41234 33416 41290 33425
rect 41234 33351 41290 33360
rect 41432 31482 41460 43726
rect 41512 32496 41564 32502
rect 41512 32438 41564 32444
rect 41524 31890 41552 32438
rect 41512 31884 41564 31890
rect 41512 31826 41564 31832
rect 41524 31482 41552 31826
rect 41708 31754 41736 53926
rect 42950 53884 43258 53893
rect 42950 53882 42956 53884
rect 43012 53882 43036 53884
rect 43092 53882 43116 53884
rect 43172 53882 43196 53884
rect 43252 53882 43258 53884
rect 43012 53830 43014 53882
rect 43194 53830 43196 53882
rect 42950 53828 42956 53830
rect 43012 53828 43036 53830
rect 43092 53828 43116 53830
rect 43172 53828 43196 53830
rect 43252 53828 43258 53830
rect 42950 53819 43258 53828
rect 43444 53440 43496 53446
rect 43444 53382 43496 53388
rect 42950 52796 43258 52805
rect 42950 52794 42956 52796
rect 43012 52794 43036 52796
rect 43092 52794 43116 52796
rect 43172 52794 43196 52796
rect 43252 52794 43258 52796
rect 43012 52742 43014 52794
rect 43194 52742 43196 52794
rect 42950 52740 42956 52742
rect 43012 52740 43036 52742
rect 43092 52740 43116 52742
rect 43172 52740 43196 52742
rect 43252 52740 43258 52742
rect 42950 52731 43258 52740
rect 42950 51708 43258 51717
rect 42950 51706 42956 51708
rect 43012 51706 43036 51708
rect 43092 51706 43116 51708
rect 43172 51706 43196 51708
rect 43252 51706 43258 51708
rect 43012 51654 43014 51706
rect 43194 51654 43196 51706
rect 42950 51652 42956 51654
rect 43012 51652 43036 51654
rect 43092 51652 43116 51654
rect 43172 51652 43196 51654
rect 43252 51652 43258 51654
rect 42950 51643 43258 51652
rect 42950 50620 43258 50629
rect 42950 50618 42956 50620
rect 43012 50618 43036 50620
rect 43092 50618 43116 50620
rect 43172 50618 43196 50620
rect 43252 50618 43258 50620
rect 43012 50566 43014 50618
rect 43194 50566 43196 50618
rect 42950 50564 42956 50566
rect 43012 50564 43036 50566
rect 43092 50564 43116 50566
rect 43172 50564 43196 50566
rect 43252 50564 43258 50566
rect 42950 50555 43258 50564
rect 42950 49532 43258 49541
rect 42950 49530 42956 49532
rect 43012 49530 43036 49532
rect 43092 49530 43116 49532
rect 43172 49530 43196 49532
rect 43252 49530 43258 49532
rect 43012 49478 43014 49530
rect 43194 49478 43196 49530
rect 42950 49476 42956 49478
rect 43012 49476 43036 49478
rect 43092 49476 43116 49478
rect 43172 49476 43196 49478
rect 43252 49476 43258 49478
rect 42950 49467 43258 49476
rect 42950 48444 43258 48453
rect 42950 48442 42956 48444
rect 43012 48442 43036 48444
rect 43092 48442 43116 48444
rect 43172 48442 43196 48444
rect 43252 48442 43258 48444
rect 43012 48390 43014 48442
rect 43194 48390 43196 48442
rect 42950 48388 42956 48390
rect 43012 48388 43036 48390
rect 43092 48388 43116 48390
rect 43172 48388 43196 48390
rect 43252 48388 43258 48390
rect 42950 48379 43258 48388
rect 42950 47356 43258 47365
rect 42950 47354 42956 47356
rect 43012 47354 43036 47356
rect 43092 47354 43116 47356
rect 43172 47354 43196 47356
rect 43252 47354 43258 47356
rect 43012 47302 43014 47354
rect 43194 47302 43196 47354
rect 42950 47300 42956 47302
rect 43012 47300 43036 47302
rect 43092 47300 43116 47302
rect 43172 47300 43196 47302
rect 43252 47300 43258 47302
rect 42950 47291 43258 47300
rect 42950 46268 43258 46277
rect 42950 46266 42956 46268
rect 43012 46266 43036 46268
rect 43092 46266 43116 46268
rect 43172 46266 43196 46268
rect 43252 46266 43258 46268
rect 43012 46214 43014 46266
rect 43194 46214 43196 46266
rect 42950 46212 42956 46214
rect 43012 46212 43036 46214
rect 43092 46212 43116 46214
rect 43172 46212 43196 46214
rect 43252 46212 43258 46214
rect 42950 46203 43258 46212
rect 42950 45180 43258 45189
rect 42950 45178 42956 45180
rect 43012 45178 43036 45180
rect 43092 45178 43116 45180
rect 43172 45178 43196 45180
rect 43252 45178 43258 45180
rect 43012 45126 43014 45178
rect 43194 45126 43196 45178
rect 42950 45124 42956 45126
rect 43012 45124 43036 45126
rect 43092 45124 43116 45126
rect 43172 45124 43196 45126
rect 43252 45124 43258 45126
rect 42950 45115 43258 45124
rect 42950 44092 43258 44101
rect 42950 44090 42956 44092
rect 43012 44090 43036 44092
rect 43092 44090 43116 44092
rect 43172 44090 43196 44092
rect 43252 44090 43258 44092
rect 43012 44038 43014 44090
rect 43194 44038 43196 44090
rect 42950 44036 42956 44038
rect 43012 44036 43036 44038
rect 43092 44036 43116 44038
rect 43172 44036 43196 44038
rect 43252 44036 43258 44038
rect 42950 44027 43258 44036
rect 43456 43858 43484 53382
rect 43444 43852 43496 43858
rect 43444 43794 43496 43800
rect 42800 43716 42852 43722
rect 42800 43658 42852 43664
rect 42708 34060 42760 34066
rect 42708 34002 42760 34008
rect 41788 32360 41840 32366
rect 41788 32302 41840 32308
rect 41800 31958 41828 32302
rect 41788 31952 41840 31958
rect 41788 31894 41840 31900
rect 41880 31952 41932 31958
rect 41880 31894 41932 31900
rect 41616 31726 41736 31754
rect 41420 31476 41472 31482
rect 41420 31418 41472 31424
rect 41512 31476 41564 31482
rect 41512 31418 41564 31424
rect 41432 30802 41460 31418
rect 41420 30796 41472 30802
rect 41420 30738 41472 30744
rect 41432 30258 41460 30738
rect 41420 30252 41472 30258
rect 41420 30194 41472 30200
rect 41512 30048 41564 30054
rect 41512 29990 41564 29996
rect 41524 29850 41552 29990
rect 41512 29844 41564 29850
rect 41512 29786 41564 29792
rect 41616 29782 41644 31726
rect 41696 30660 41748 30666
rect 41696 30602 41748 30608
rect 41708 30054 41736 30602
rect 41696 30048 41748 30054
rect 41696 29990 41748 29996
rect 41604 29776 41656 29782
rect 41604 29718 41656 29724
rect 41512 29708 41564 29714
rect 41512 29650 41564 29656
rect 41524 29510 41552 29650
rect 41512 29504 41564 29510
rect 41512 29446 41564 29452
rect 41420 29232 41472 29238
rect 41708 29186 41736 29990
rect 41420 29174 41472 29180
rect 41432 28558 41460 29174
rect 41616 29158 41736 29186
rect 41420 28552 41472 28558
rect 41420 28494 41472 28500
rect 41512 28076 41564 28082
rect 41512 28018 41564 28024
rect 40960 27396 41012 27402
rect 40960 27338 41012 27344
rect 41144 26784 41196 26790
rect 41144 26726 41196 26732
rect 40684 25356 40736 25362
rect 40684 25298 40736 25304
rect 40592 25220 40644 25226
rect 40592 25162 40644 25168
rect 40500 23792 40552 23798
rect 40500 23734 40552 23740
rect 40696 23662 40724 25298
rect 40040 23588 40092 23594
rect 40040 23530 40092 23536
rect 40328 23582 40448 23610
rect 40684 23656 40736 23662
rect 40684 23598 40736 23604
rect 40052 23186 40080 23530
rect 39304 23180 39356 23186
rect 39304 23122 39356 23128
rect 40040 23180 40092 23186
rect 40040 23122 40092 23128
rect 39316 22574 39344 23122
rect 40052 22778 40080 23122
rect 40132 23112 40184 23118
rect 40132 23054 40184 23060
rect 40144 22778 40172 23054
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 40132 22772 40184 22778
rect 40132 22714 40184 22720
rect 39304 22568 39356 22574
rect 39304 22510 39356 22516
rect 39396 22568 39448 22574
rect 39396 22510 39448 22516
rect 39316 22166 39344 22510
rect 39304 22160 39356 22166
rect 39304 22102 39356 22108
rect 39408 22098 39436 22510
rect 39672 22432 39724 22438
rect 39672 22374 39724 22380
rect 39488 22228 39540 22234
rect 39488 22170 39540 22176
rect 39212 22092 39264 22098
rect 39212 22034 39264 22040
rect 39396 22092 39448 22098
rect 39396 22034 39448 22040
rect 39120 22024 39172 22030
rect 39120 21966 39172 21972
rect 39028 21684 39080 21690
rect 39028 21626 39080 21632
rect 38844 21616 38896 21622
rect 38844 21558 38896 21564
rect 38752 21480 38804 21486
rect 38752 21422 38804 21428
rect 39028 21480 39080 21486
rect 39028 21422 39080 21428
rect 38764 20874 38792 21422
rect 38844 21412 38896 21418
rect 38844 21354 38896 21360
rect 38752 20868 38804 20874
rect 38752 20810 38804 20816
rect 38660 20528 38712 20534
rect 38660 20470 38712 20476
rect 38672 17746 38700 20470
rect 38764 20398 38792 20810
rect 38752 20392 38804 20398
rect 38752 20334 38804 20340
rect 38856 19854 38884 21354
rect 38844 19848 38896 19854
rect 38844 19790 38896 19796
rect 38844 18284 38896 18290
rect 38844 18226 38896 18232
rect 38660 17740 38712 17746
rect 38660 17682 38712 17688
rect 38568 17332 38620 17338
rect 38568 17274 38620 17280
rect 38476 16652 38528 16658
rect 38476 16594 38528 16600
rect 38580 15026 38608 17274
rect 38856 17202 38884 18226
rect 38844 17196 38896 17202
rect 38844 17138 38896 17144
rect 39040 17066 39068 21422
rect 39212 21344 39264 21350
rect 39212 21286 39264 21292
rect 39028 17060 39080 17066
rect 39028 17002 39080 17008
rect 38660 15428 38712 15434
rect 38660 15370 38712 15376
rect 38672 15162 38700 15370
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 39040 15094 39068 17002
rect 39028 15088 39080 15094
rect 38948 15036 39028 15042
rect 38948 15030 39080 15036
rect 38568 15020 38620 15026
rect 38568 14962 38620 14968
rect 38948 15014 39068 15030
rect 38580 14482 38608 14962
rect 38568 14476 38620 14482
rect 38568 14418 38620 14424
rect 38580 13938 38608 14418
rect 38752 14272 38804 14278
rect 38752 14214 38804 14220
rect 38844 14272 38896 14278
rect 38844 14214 38896 14220
rect 38764 14074 38792 14214
rect 38752 14068 38804 14074
rect 38752 14010 38804 14016
rect 38568 13932 38620 13938
rect 38568 13874 38620 13880
rect 38660 13524 38712 13530
rect 38660 13466 38712 13472
rect 38672 12850 38700 13466
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 38476 12096 38528 12102
rect 38476 12038 38528 12044
rect 38488 11830 38516 12038
rect 38476 11824 38528 11830
rect 38476 11766 38528 11772
rect 38568 11756 38620 11762
rect 38568 11698 38620 11704
rect 38384 9648 38436 9654
rect 38384 9590 38436 9596
rect 38476 8900 38528 8906
rect 38476 8842 38528 8848
rect 38488 8566 38516 8842
rect 38476 8560 38528 8566
rect 38476 8502 38528 8508
rect 38292 6384 38344 6390
rect 38292 6326 38344 6332
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 37648 5024 37700 5030
rect 37648 4966 37700 4972
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 38580 3534 38608 11698
rect 38672 11150 38700 12786
rect 38856 11286 38884 14214
rect 38948 11558 38976 15014
rect 39224 14482 39252 21286
rect 39500 19122 39528 22170
rect 39684 19854 39712 22374
rect 40040 20936 40092 20942
rect 40040 20878 40092 20884
rect 39948 20460 40000 20466
rect 39948 20402 40000 20408
rect 39960 20058 39988 20402
rect 40052 20262 40080 20878
rect 40040 20256 40092 20262
rect 40040 20198 40092 20204
rect 40132 20256 40184 20262
rect 40132 20198 40184 20204
rect 39948 20052 40000 20058
rect 39948 19994 40000 20000
rect 40052 19922 40080 20198
rect 40144 20058 40172 20198
rect 40132 20052 40184 20058
rect 40132 19994 40184 20000
rect 40040 19916 40092 19922
rect 40040 19858 40092 19864
rect 39672 19848 39724 19854
rect 39672 19790 39724 19796
rect 39408 19094 39528 19122
rect 39408 16114 39436 19094
rect 39488 18624 39540 18630
rect 39488 18566 39540 18572
rect 39396 16108 39448 16114
rect 39396 16050 39448 16056
rect 39396 14816 39448 14822
rect 39396 14758 39448 14764
rect 39408 14482 39436 14758
rect 39212 14476 39264 14482
rect 39212 14418 39264 14424
rect 39396 14476 39448 14482
rect 39396 14418 39448 14424
rect 39120 14408 39172 14414
rect 39120 14350 39172 14356
rect 39028 13932 39080 13938
rect 39028 13874 39080 13880
rect 39040 13394 39068 13874
rect 39028 13388 39080 13394
rect 39028 13330 39080 13336
rect 39040 12850 39068 13330
rect 39028 12844 39080 12850
rect 39028 12786 39080 12792
rect 39132 11762 39160 14350
rect 39408 14006 39436 14418
rect 39396 14000 39448 14006
rect 39396 13942 39448 13948
rect 39500 13326 39528 18566
rect 39948 18148 40000 18154
rect 39948 18090 40000 18096
rect 39672 17332 39724 17338
rect 39672 17274 39724 17280
rect 39684 17202 39712 17274
rect 39672 17196 39724 17202
rect 39672 17138 39724 17144
rect 39960 17134 39988 18090
rect 39948 17128 40000 17134
rect 39948 17070 40000 17076
rect 39960 16658 39988 17070
rect 39948 16652 40000 16658
rect 39948 16594 40000 16600
rect 40328 16590 40356 23582
rect 40868 23316 40920 23322
rect 40868 23258 40920 23264
rect 40776 23044 40828 23050
rect 40776 22986 40828 22992
rect 40592 22704 40644 22710
rect 40592 22646 40644 22652
rect 40408 22432 40460 22438
rect 40408 22374 40460 22380
rect 40420 22234 40448 22374
rect 40408 22228 40460 22234
rect 40408 22170 40460 22176
rect 40604 21554 40632 22646
rect 40788 22574 40816 22986
rect 40776 22568 40828 22574
rect 40776 22510 40828 22516
rect 40592 21548 40644 21554
rect 40592 21490 40644 21496
rect 40500 20868 40552 20874
rect 40500 20810 40552 20816
rect 40512 19718 40540 20810
rect 40592 19780 40644 19786
rect 40592 19722 40644 19728
rect 40500 19712 40552 19718
rect 40500 19654 40552 19660
rect 40604 19553 40632 19722
rect 40590 19544 40646 19553
rect 40590 19479 40646 19488
rect 40880 18834 40908 23258
rect 41052 19712 41104 19718
rect 41052 19654 41104 19660
rect 41064 18834 41092 19654
rect 40868 18828 40920 18834
rect 40868 18770 40920 18776
rect 41052 18828 41104 18834
rect 41052 18770 41104 18776
rect 40408 18692 40460 18698
rect 40408 18634 40460 18640
rect 40420 17678 40448 18634
rect 40868 18624 40920 18630
rect 40868 18566 40920 18572
rect 40880 18222 40908 18566
rect 41156 18290 41184 26726
rect 41420 26240 41472 26246
rect 41420 26182 41472 26188
rect 41432 25974 41460 26182
rect 41420 25968 41472 25974
rect 41420 25910 41472 25916
rect 41524 25786 41552 28018
rect 41616 26926 41644 29158
rect 41788 27872 41840 27878
rect 41788 27814 41840 27820
rect 41696 27464 41748 27470
rect 41696 27406 41748 27412
rect 41708 27130 41736 27406
rect 41696 27124 41748 27130
rect 41696 27066 41748 27072
rect 41604 26920 41656 26926
rect 41604 26862 41656 26868
rect 41432 25758 41552 25786
rect 41696 25832 41748 25838
rect 41800 25786 41828 27814
rect 41892 27130 41920 31894
rect 42720 31890 42748 34002
rect 42708 31884 42760 31890
rect 42708 31826 42760 31832
rect 42812 31414 42840 43658
rect 42950 43004 43258 43013
rect 42950 43002 42956 43004
rect 43012 43002 43036 43004
rect 43092 43002 43116 43004
rect 43172 43002 43196 43004
rect 43252 43002 43258 43004
rect 43012 42950 43014 43002
rect 43194 42950 43196 43002
rect 42950 42948 42956 42950
rect 43012 42948 43036 42950
rect 43092 42948 43116 42950
rect 43172 42948 43196 42950
rect 43252 42948 43258 42950
rect 42950 42939 43258 42948
rect 42950 41916 43258 41925
rect 42950 41914 42956 41916
rect 43012 41914 43036 41916
rect 43092 41914 43116 41916
rect 43172 41914 43196 41916
rect 43252 41914 43258 41916
rect 43012 41862 43014 41914
rect 43194 41862 43196 41914
rect 42950 41860 42956 41862
rect 43012 41860 43036 41862
rect 43092 41860 43116 41862
rect 43172 41860 43196 41862
rect 43252 41860 43258 41862
rect 42950 41851 43258 41860
rect 42950 40828 43258 40837
rect 42950 40826 42956 40828
rect 43012 40826 43036 40828
rect 43092 40826 43116 40828
rect 43172 40826 43196 40828
rect 43252 40826 43258 40828
rect 43012 40774 43014 40826
rect 43194 40774 43196 40826
rect 42950 40772 42956 40774
rect 43012 40772 43036 40774
rect 43092 40772 43116 40774
rect 43172 40772 43196 40774
rect 43252 40772 43258 40774
rect 42950 40763 43258 40772
rect 42950 39740 43258 39749
rect 42950 39738 42956 39740
rect 43012 39738 43036 39740
rect 43092 39738 43116 39740
rect 43172 39738 43196 39740
rect 43252 39738 43258 39740
rect 43012 39686 43014 39738
rect 43194 39686 43196 39738
rect 42950 39684 42956 39686
rect 43012 39684 43036 39686
rect 43092 39684 43116 39686
rect 43172 39684 43196 39686
rect 43252 39684 43258 39686
rect 42950 39675 43258 39684
rect 42950 38652 43258 38661
rect 42950 38650 42956 38652
rect 43012 38650 43036 38652
rect 43092 38650 43116 38652
rect 43172 38650 43196 38652
rect 43252 38650 43258 38652
rect 43012 38598 43014 38650
rect 43194 38598 43196 38650
rect 42950 38596 42956 38598
rect 43012 38596 43036 38598
rect 43092 38596 43116 38598
rect 43172 38596 43196 38598
rect 43252 38596 43258 38598
rect 42950 38587 43258 38596
rect 42950 37564 43258 37573
rect 42950 37562 42956 37564
rect 43012 37562 43036 37564
rect 43092 37562 43116 37564
rect 43172 37562 43196 37564
rect 43252 37562 43258 37564
rect 43012 37510 43014 37562
rect 43194 37510 43196 37562
rect 42950 37508 42956 37510
rect 43012 37508 43036 37510
rect 43092 37508 43116 37510
rect 43172 37508 43196 37510
rect 43252 37508 43258 37510
rect 42950 37499 43258 37508
rect 42950 36476 43258 36485
rect 42950 36474 42956 36476
rect 43012 36474 43036 36476
rect 43092 36474 43116 36476
rect 43172 36474 43196 36476
rect 43252 36474 43258 36476
rect 43012 36422 43014 36474
rect 43194 36422 43196 36474
rect 42950 36420 42956 36422
rect 43012 36420 43036 36422
rect 43092 36420 43116 36422
rect 43172 36420 43196 36422
rect 43252 36420 43258 36422
rect 42950 36411 43258 36420
rect 42950 35388 43258 35397
rect 42950 35386 42956 35388
rect 43012 35386 43036 35388
rect 43092 35386 43116 35388
rect 43172 35386 43196 35388
rect 43252 35386 43258 35388
rect 43012 35334 43014 35386
rect 43194 35334 43196 35386
rect 42950 35332 42956 35334
rect 43012 35332 43036 35334
rect 43092 35332 43116 35334
rect 43172 35332 43196 35334
rect 43252 35332 43258 35334
rect 42950 35323 43258 35332
rect 44180 34740 44232 34746
rect 44180 34682 44232 34688
rect 42950 34300 43258 34309
rect 42950 34298 42956 34300
rect 43012 34298 43036 34300
rect 43092 34298 43116 34300
rect 43172 34298 43196 34300
rect 43252 34298 43258 34300
rect 43012 34246 43014 34298
rect 43194 34246 43196 34298
rect 42950 34244 42956 34246
rect 43012 34244 43036 34246
rect 43092 34244 43116 34246
rect 43172 34244 43196 34246
rect 43252 34244 43258 34246
rect 42950 34235 43258 34244
rect 43720 34128 43772 34134
rect 43720 34070 43772 34076
rect 42892 34060 42944 34066
rect 42892 34002 42944 34008
rect 42904 33862 42932 34002
rect 42892 33856 42944 33862
rect 42892 33798 42944 33804
rect 43628 33516 43680 33522
rect 43628 33458 43680 33464
rect 43536 33448 43588 33454
rect 43536 33390 43588 33396
rect 42950 33212 43258 33221
rect 42950 33210 42956 33212
rect 43012 33210 43036 33212
rect 43092 33210 43116 33212
rect 43172 33210 43196 33212
rect 43252 33210 43258 33212
rect 43012 33158 43014 33210
rect 43194 33158 43196 33210
rect 42950 33156 42956 33158
rect 43012 33156 43036 33158
rect 43092 33156 43116 33158
rect 43172 33156 43196 33158
rect 43252 33156 43258 33158
rect 42950 33147 43258 33156
rect 42950 32124 43258 32133
rect 42950 32122 42956 32124
rect 43012 32122 43036 32124
rect 43092 32122 43116 32124
rect 43172 32122 43196 32124
rect 43252 32122 43258 32124
rect 43012 32070 43014 32122
rect 43194 32070 43196 32122
rect 42950 32068 42956 32070
rect 43012 32068 43036 32070
rect 43092 32068 43116 32070
rect 43172 32068 43196 32070
rect 43252 32068 43258 32070
rect 42950 32059 43258 32068
rect 42892 32020 42944 32026
rect 42892 31962 42944 31968
rect 42904 31822 42932 31962
rect 43352 31884 43404 31890
rect 43352 31826 43404 31832
rect 42892 31816 42944 31822
rect 42892 31758 42944 31764
rect 42904 31414 42932 31758
rect 42800 31408 42852 31414
rect 42800 31350 42852 31356
rect 42892 31408 42944 31414
rect 42892 31350 42944 31356
rect 42524 31204 42576 31210
rect 42524 31146 42576 31152
rect 41972 29572 42024 29578
rect 41972 29514 42024 29520
rect 41984 27470 42012 29514
rect 42432 28960 42484 28966
rect 42432 28902 42484 28908
rect 42064 28756 42116 28762
rect 42064 28698 42116 28704
rect 42076 27946 42104 28698
rect 42444 28422 42472 28902
rect 42536 28490 42564 31146
rect 42812 30734 42840 31350
rect 42950 31036 43258 31045
rect 42950 31034 42956 31036
rect 43012 31034 43036 31036
rect 43092 31034 43116 31036
rect 43172 31034 43196 31036
rect 43252 31034 43258 31036
rect 43012 30982 43014 31034
rect 43194 30982 43196 31034
rect 42950 30980 42956 30982
rect 43012 30980 43036 30982
rect 43092 30980 43116 30982
rect 43172 30980 43196 30982
rect 43252 30980 43258 30982
rect 42950 30971 43258 30980
rect 42800 30728 42852 30734
rect 42800 30670 42852 30676
rect 43364 30546 43392 31826
rect 43548 31278 43576 33390
rect 43640 33318 43668 33458
rect 43628 33312 43680 33318
rect 43628 33254 43680 33260
rect 43536 31272 43588 31278
rect 43536 31214 43588 31220
rect 43444 31136 43496 31142
rect 43444 31078 43496 31084
rect 42996 30518 43392 30546
rect 42616 30252 42668 30258
rect 42616 30194 42668 30200
rect 42628 29714 42656 30194
rect 42996 30190 43024 30518
rect 43260 30388 43312 30394
rect 43260 30330 43312 30336
rect 42984 30184 43036 30190
rect 42984 30126 43036 30132
rect 43272 30138 43300 30330
rect 43272 30110 43392 30138
rect 42950 29948 43258 29957
rect 42950 29946 42956 29948
rect 43012 29946 43036 29948
rect 43092 29946 43116 29948
rect 43172 29946 43196 29948
rect 43252 29946 43258 29948
rect 43012 29894 43014 29946
rect 43194 29894 43196 29946
rect 42950 29892 42956 29894
rect 43012 29892 43036 29894
rect 43092 29892 43116 29894
rect 43172 29892 43196 29894
rect 43252 29892 43258 29894
rect 42950 29883 43258 29892
rect 42616 29708 42668 29714
rect 42616 29650 42668 29656
rect 42628 29170 42656 29650
rect 42616 29164 42668 29170
rect 42616 29106 42668 29112
rect 42628 28626 42656 29106
rect 42950 28860 43258 28869
rect 42950 28858 42956 28860
rect 43012 28858 43036 28860
rect 43092 28858 43116 28860
rect 43172 28858 43196 28860
rect 43252 28858 43258 28860
rect 43012 28806 43014 28858
rect 43194 28806 43196 28858
rect 42950 28804 42956 28806
rect 43012 28804 43036 28806
rect 43092 28804 43116 28806
rect 43172 28804 43196 28806
rect 43252 28804 43258 28806
rect 42950 28795 43258 28804
rect 42616 28620 42668 28626
rect 42616 28562 42668 28568
rect 42524 28484 42576 28490
rect 42524 28426 42576 28432
rect 42432 28416 42484 28422
rect 42432 28358 42484 28364
rect 42064 27940 42116 27946
rect 42064 27882 42116 27888
rect 41972 27464 42024 27470
rect 41972 27406 42024 27412
rect 41880 27124 41932 27130
rect 41880 27066 41932 27072
rect 41880 25968 41932 25974
rect 41880 25910 41932 25916
rect 41748 25780 41828 25786
rect 41696 25774 41828 25780
rect 41708 25758 41828 25774
rect 41328 23588 41380 23594
rect 41328 23530 41380 23536
rect 41340 22030 41368 23530
rect 41432 22778 41460 25758
rect 41800 25430 41828 25758
rect 41788 25424 41840 25430
rect 41788 25366 41840 25372
rect 41892 25226 41920 25910
rect 41880 25220 41932 25226
rect 41880 25162 41932 25168
rect 41892 24886 41920 25162
rect 41880 24880 41932 24886
rect 41880 24822 41932 24828
rect 41696 24812 41748 24818
rect 41696 24754 41748 24760
rect 41512 23180 41564 23186
rect 41512 23122 41564 23128
rect 41420 22772 41472 22778
rect 41420 22714 41472 22720
rect 41524 22642 41552 23122
rect 41708 22778 41736 24754
rect 41892 23118 41920 24822
rect 41984 23798 42012 27406
rect 42444 25838 42472 28358
rect 42616 27872 42668 27878
rect 42616 27814 42668 27820
rect 42524 26376 42576 26382
rect 42524 26318 42576 26324
rect 42536 26042 42564 26318
rect 42524 26036 42576 26042
rect 42524 25978 42576 25984
rect 42432 25832 42484 25838
rect 42432 25774 42484 25780
rect 42064 24676 42116 24682
rect 42064 24618 42116 24624
rect 41972 23792 42024 23798
rect 41972 23734 42024 23740
rect 41880 23112 41932 23118
rect 41880 23054 41932 23060
rect 41696 22772 41748 22778
rect 41696 22714 41748 22720
rect 41512 22636 41564 22642
rect 41512 22578 41564 22584
rect 41328 22024 41380 22030
rect 41328 21966 41380 21972
rect 41524 21978 41552 22578
rect 41340 19922 41368 21966
rect 41524 21962 41644 21978
rect 41524 21956 41656 21962
rect 41524 21950 41604 21956
rect 41604 21898 41656 21904
rect 41616 20942 41644 21898
rect 41604 20936 41656 20942
rect 41604 20878 41656 20884
rect 41616 20534 41644 20878
rect 41604 20528 41656 20534
rect 41604 20470 41656 20476
rect 41328 19916 41380 19922
rect 41328 19858 41380 19864
rect 41340 19802 41368 19858
rect 41616 19854 41644 20470
rect 41604 19848 41656 19854
rect 41340 19774 41414 19802
rect 41604 19790 41656 19796
rect 41386 19700 41414 19774
rect 41386 19672 41460 19700
rect 41432 18834 41460 19672
rect 41420 18828 41472 18834
rect 41420 18770 41472 18776
rect 41432 18290 41460 18770
rect 41144 18284 41196 18290
rect 41144 18226 41196 18232
rect 41420 18284 41472 18290
rect 41420 18226 41472 18232
rect 40776 18216 40828 18222
rect 40776 18158 40828 18164
rect 40868 18216 40920 18222
rect 40868 18158 40920 18164
rect 40408 17672 40460 17678
rect 40408 17614 40460 17620
rect 40408 17264 40460 17270
rect 40408 17206 40460 17212
rect 40420 17134 40448 17206
rect 40408 17128 40460 17134
rect 40408 17070 40460 17076
rect 40316 16584 40368 16590
rect 40316 16526 40368 16532
rect 40040 16448 40092 16454
rect 40040 16390 40092 16396
rect 40224 16448 40276 16454
rect 40224 16390 40276 16396
rect 39488 13320 39540 13326
rect 39488 13262 39540 13268
rect 39212 13184 39264 13190
rect 39212 13126 39264 13132
rect 39120 11756 39172 11762
rect 39120 11698 39172 11704
rect 38936 11552 38988 11558
rect 38936 11494 38988 11500
rect 38844 11280 38896 11286
rect 38844 11222 38896 11228
rect 38660 11144 38712 11150
rect 38660 11086 38712 11092
rect 38936 11144 38988 11150
rect 38936 11086 38988 11092
rect 38844 11076 38896 11082
rect 38844 11018 38896 11024
rect 38752 10532 38804 10538
rect 38752 10474 38804 10480
rect 38660 10056 38712 10062
rect 38660 9998 38712 10004
rect 38672 8974 38700 9998
rect 38764 9654 38792 10474
rect 38752 9648 38804 9654
rect 38752 9590 38804 9596
rect 38660 8968 38712 8974
rect 38660 8910 38712 8916
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 38856 3058 38884 11018
rect 38948 8974 38976 11086
rect 39120 9716 39172 9722
rect 39224 9704 39252 13126
rect 39304 12232 39356 12238
rect 39304 12174 39356 12180
rect 39316 11898 39344 12174
rect 39304 11892 39356 11898
rect 39304 11834 39356 11840
rect 39488 11212 39540 11218
rect 39488 11154 39540 11160
rect 39172 9676 39252 9704
rect 39120 9658 39172 9664
rect 39028 9648 39080 9654
rect 39028 9590 39080 9596
rect 38936 8968 38988 8974
rect 38936 8910 38988 8916
rect 39040 8906 39068 9590
rect 39120 9376 39172 9382
rect 39120 9318 39172 9324
rect 39028 8900 39080 8906
rect 39028 8842 39080 8848
rect 39028 7200 39080 7206
rect 39028 7142 39080 7148
rect 39040 6798 39068 7142
rect 39132 6798 39160 9318
rect 39028 6792 39080 6798
rect 39028 6734 39080 6740
rect 39120 6792 39172 6798
rect 39120 6734 39172 6740
rect 38936 6724 38988 6730
rect 38936 6666 38988 6672
rect 38948 4146 38976 6666
rect 39224 5710 39252 9676
rect 39500 6390 39528 11154
rect 40052 9518 40080 16390
rect 40236 12646 40264 16390
rect 40420 15094 40448 17070
rect 40500 16516 40552 16522
rect 40500 16458 40552 16464
rect 40408 15088 40460 15094
rect 40408 15030 40460 15036
rect 40420 13938 40448 15030
rect 40408 13932 40460 13938
rect 40408 13874 40460 13880
rect 40224 12640 40276 12646
rect 40224 12582 40276 12588
rect 40420 12434 40448 13874
rect 40512 13326 40540 16458
rect 40788 16114 40816 18158
rect 41328 17740 41380 17746
rect 41328 17682 41380 17688
rect 41052 17060 41104 17066
rect 41052 17002 41104 17008
rect 40776 16108 40828 16114
rect 40776 16050 40828 16056
rect 40868 15632 40920 15638
rect 40868 15574 40920 15580
rect 40592 13932 40644 13938
rect 40592 13874 40644 13880
rect 40500 13320 40552 13326
rect 40500 13262 40552 13268
rect 40500 13184 40552 13190
rect 40500 13126 40552 13132
rect 40328 12406 40448 12434
rect 40132 10804 40184 10810
rect 40132 10746 40184 10752
rect 40040 9512 40092 9518
rect 40040 9454 40092 9460
rect 40040 9104 40092 9110
rect 40040 9046 40092 9052
rect 40052 6798 40080 9046
rect 40144 8566 40172 10746
rect 40328 10674 40356 12406
rect 40316 10668 40368 10674
rect 40316 10610 40368 10616
rect 40408 9920 40460 9926
rect 40408 9862 40460 9868
rect 40224 9376 40276 9382
rect 40224 9318 40276 9324
rect 40132 8560 40184 8566
rect 40132 8502 40184 8508
rect 40236 8498 40264 9318
rect 40316 8968 40368 8974
rect 40316 8910 40368 8916
rect 40328 8634 40356 8910
rect 40316 8628 40368 8634
rect 40316 8570 40368 8576
rect 40224 8492 40276 8498
rect 40224 8434 40276 8440
rect 40224 7880 40276 7886
rect 40224 7822 40276 7828
rect 40236 7274 40264 7822
rect 40224 7268 40276 7274
rect 40224 7210 40276 7216
rect 40040 6792 40092 6798
rect 40040 6734 40092 6740
rect 39488 6384 39540 6390
rect 39488 6326 39540 6332
rect 40040 6248 40092 6254
rect 40040 6190 40092 6196
rect 39488 6180 39540 6186
rect 39488 6122 39540 6128
rect 39212 5704 39264 5710
rect 39212 5646 39264 5652
rect 38936 4140 38988 4146
rect 38936 4082 38988 4088
rect 39028 4072 39080 4078
rect 39028 4014 39080 4020
rect 38844 3052 38896 3058
rect 38844 2994 38896 3000
rect 36820 2984 36872 2990
rect 36820 2926 36872 2932
rect 36268 2440 36320 2446
rect 36268 2382 36320 2388
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 36832 800 36860 2926
rect 37556 2916 37608 2922
rect 37556 2858 37608 2864
rect 37568 800 37596 2858
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38304 800 38332 2246
rect 39040 800 39068 4014
rect 39500 2378 39528 6122
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39488 2372 39540 2378
rect 39488 2314 39540 2320
rect 39776 800 39804 3538
rect 40052 3534 40080 6190
rect 40224 5908 40276 5914
rect 40224 5850 40276 5856
rect 40132 5772 40184 5778
rect 40132 5714 40184 5720
rect 40144 3534 40172 5714
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 40236 2582 40264 5850
rect 40420 5778 40448 9862
rect 40512 8945 40540 13126
rect 40604 12850 40632 13874
rect 40684 13864 40736 13870
rect 40684 13806 40736 13812
rect 40592 12844 40644 12850
rect 40592 12786 40644 12792
rect 40696 12730 40724 13806
rect 40776 13728 40828 13734
rect 40776 13670 40828 13676
rect 40788 12782 40816 13670
rect 40880 12850 40908 15574
rect 40960 14272 41012 14278
rect 40960 14214 41012 14220
rect 40868 12844 40920 12850
rect 40868 12786 40920 12792
rect 40604 12702 40724 12730
rect 40776 12776 40828 12782
rect 40776 12718 40828 12724
rect 40604 11898 40632 12702
rect 40684 12640 40736 12646
rect 40684 12582 40736 12588
rect 40592 11892 40644 11898
rect 40592 11834 40644 11840
rect 40696 11694 40724 12582
rect 40868 12096 40920 12102
rect 40868 12038 40920 12044
rect 40684 11688 40736 11694
rect 40684 11630 40736 11636
rect 40696 10606 40724 11630
rect 40684 10600 40736 10606
rect 40684 10542 40736 10548
rect 40498 8936 40554 8945
rect 40498 8871 40554 8880
rect 40408 5772 40460 5778
rect 40408 5714 40460 5720
rect 40512 5574 40540 8871
rect 40880 8537 40908 12038
rect 40972 11218 41000 14214
rect 41064 12238 41092 17002
rect 41340 16794 41368 17682
rect 41328 16788 41380 16794
rect 41328 16730 41380 16736
rect 41156 14606 41368 14634
rect 41156 14482 41184 14606
rect 41236 14544 41288 14550
rect 41236 14486 41288 14492
rect 41144 14476 41196 14482
rect 41144 14418 41196 14424
rect 41248 14414 41276 14486
rect 41340 14482 41368 14606
rect 41328 14476 41380 14482
rect 41328 14418 41380 14424
rect 41236 14408 41288 14414
rect 41236 14350 41288 14356
rect 41052 12232 41104 12238
rect 41052 12174 41104 12180
rect 40960 11212 41012 11218
rect 40960 11154 41012 11160
rect 40866 8528 40922 8537
rect 40866 8463 40922 8472
rect 40592 6656 40644 6662
rect 40592 6598 40644 6604
rect 40604 5710 40632 6598
rect 40592 5704 40644 5710
rect 40592 5646 40644 5652
rect 40500 5568 40552 5574
rect 40500 5510 40552 5516
rect 40880 5302 40908 8463
rect 41236 8356 41288 8362
rect 41236 8298 41288 8304
rect 41248 7410 41276 8298
rect 41236 7404 41288 7410
rect 41236 7346 41288 7352
rect 40868 5296 40920 5302
rect 40868 5238 40920 5244
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 40224 2576 40276 2582
rect 40224 2518 40276 2524
rect 40592 2508 40644 2514
rect 40512 2468 40592 2496
rect 40512 800 40540 2468
rect 40592 2450 40644 2456
rect 41248 800 41276 3538
rect 41708 2774 41736 22714
rect 42076 22166 42104 24618
rect 42064 22160 42116 22166
rect 42064 22102 42116 22108
rect 41788 21412 41840 21418
rect 41788 21354 41840 21360
rect 41800 20058 41828 21354
rect 42076 21146 42104 22102
rect 42064 21140 42116 21146
rect 42064 21082 42116 21088
rect 42156 20256 42208 20262
rect 42156 20198 42208 20204
rect 41788 20052 41840 20058
rect 41788 19994 41840 20000
rect 41800 18970 41828 19994
rect 41788 18964 41840 18970
rect 41788 18906 41840 18912
rect 42168 14346 42196 20198
rect 42340 19168 42392 19174
rect 42340 19110 42392 19116
rect 42156 14340 42208 14346
rect 42156 14282 42208 14288
rect 42352 13394 42380 19110
rect 42524 17808 42576 17814
rect 42524 17750 42576 17756
rect 42536 15366 42564 17750
rect 42628 16658 42656 27814
rect 42950 27772 43258 27781
rect 42950 27770 42956 27772
rect 43012 27770 43036 27772
rect 43092 27770 43116 27772
rect 43172 27770 43196 27772
rect 43252 27770 43258 27772
rect 43012 27718 43014 27770
rect 43194 27718 43196 27770
rect 42950 27716 42956 27718
rect 43012 27716 43036 27718
rect 43092 27716 43116 27718
rect 43172 27716 43196 27718
rect 43252 27716 43258 27718
rect 42950 27707 43258 27716
rect 42708 27396 42760 27402
rect 42708 27338 42760 27344
rect 42720 26450 42748 27338
rect 42950 26684 43258 26693
rect 42950 26682 42956 26684
rect 43012 26682 43036 26684
rect 43092 26682 43116 26684
rect 43172 26682 43196 26684
rect 43252 26682 43258 26684
rect 43012 26630 43014 26682
rect 43194 26630 43196 26682
rect 42950 26628 42956 26630
rect 43012 26628 43036 26630
rect 43092 26628 43116 26630
rect 43172 26628 43196 26630
rect 43252 26628 43258 26630
rect 42950 26619 43258 26628
rect 43364 26450 43392 30110
rect 42708 26444 42760 26450
rect 42708 26386 42760 26392
rect 42892 26444 42944 26450
rect 42892 26386 42944 26392
rect 43352 26444 43404 26450
rect 43352 26386 43404 26392
rect 42720 26042 42748 26386
rect 42708 26036 42760 26042
rect 42708 25978 42760 25984
rect 42904 25684 42932 26386
rect 43352 26308 43404 26314
rect 43352 26250 43404 26256
rect 42885 25656 42932 25684
rect 42885 25480 42913 25656
rect 42950 25596 43258 25605
rect 42950 25594 42956 25596
rect 43012 25594 43036 25596
rect 43092 25594 43116 25596
rect 43172 25594 43196 25596
rect 43252 25594 43258 25596
rect 43012 25542 43014 25594
rect 43194 25542 43196 25594
rect 42950 25540 42956 25542
rect 43012 25540 43036 25542
rect 43092 25540 43116 25542
rect 43172 25540 43196 25542
rect 43252 25540 43258 25542
rect 42950 25531 43258 25540
rect 42885 25452 43024 25480
rect 42996 25129 43024 25452
rect 42982 25120 43038 25129
rect 42982 25055 43038 25064
rect 42996 24818 43024 25055
rect 42984 24812 43036 24818
rect 42984 24754 43036 24760
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 43168 24404 43220 24410
rect 43168 24346 43220 24352
rect 42800 24268 42852 24274
rect 42800 24210 42852 24216
rect 42812 23254 42840 24210
rect 43180 24138 43208 24346
rect 43260 24200 43312 24206
rect 43260 24142 43312 24148
rect 43168 24132 43220 24138
rect 43168 24074 43220 24080
rect 43272 23576 43300 24142
rect 43364 24070 43392 26250
rect 43456 25702 43484 31078
rect 43548 30938 43576 31214
rect 43536 30932 43588 30938
rect 43536 30874 43588 30880
rect 43640 30818 43668 33254
rect 43732 31482 43760 34070
rect 43812 33856 43864 33862
rect 43812 33798 43864 33804
rect 43720 31476 43772 31482
rect 43720 31418 43772 31424
rect 43548 30790 43668 30818
rect 43548 30394 43576 30790
rect 43628 30728 43680 30734
rect 43628 30670 43680 30676
rect 43536 30388 43588 30394
rect 43536 30330 43588 30336
rect 43640 30326 43668 30670
rect 43628 30320 43680 30326
rect 43628 30262 43680 30268
rect 43536 30184 43588 30190
rect 43536 30126 43588 30132
rect 43548 29306 43576 30126
rect 43536 29300 43588 29306
rect 43536 29242 43588 29248
rect 43640 29238 43668 30262
rect 43628 29232 43680 29238
rect 43628 29174 43680 29180
rect 43640 28762 43668 29174
rect 43628 28756 43680 28762
rect 43628 28698 43680 28704
rect 43640 28558 43668 28698
rect 43628 28552 43680 28558
rect 43628 28494 43680 28500
rect 43732 27470 43760 31418
rect 43720 27464 43772 27470
rect 43720 27406 43772 27412
rect 43628 26784 43680 26790
rect 43628 26726 43680 26732
rect 43536 25832 43588 25838
rect 43536 25774 43588 25780
rect 43444 25696 43496 25702
rect 43444 25638 43496 25644
rect 43444 24744 43496 24750
rect 43444 24686 43496 24692
rect 43352 24064 43404 24070
rect 43352 24006 43404 24012
rect 43272 23548 43392 23576
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 42800 23248 42852 23254
rect 42800 23190 42852 23196
rect 42812 22234 42840 23190
rect 42984 23112 43036 23118
rect 42984 23054 43036 23060
rect 42996 22778 43024 23054
rect 42984 22772 43036 22778
rect 42984 22714 43036 22720
rect 43364 22574 43392 23548
rect 43456 23526 43484 24686
rect 43548 24206 43576 25774
rect 43536 24200 43588 24206
rect 43536 24142 43588 24148
rect 43536 24064 43588 24070
rect 43536 24006 43588 24012
rect 43444 23520 43496 23526
rect 43444 23462 43496 23468
rect 43352 22568 43404 22574
rect 43352 22510 43404 22516
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42800 22228 42852 22234
rect 42800 22170 42852 22176
rect 42800 21344 42852 21350
rect 42800 21286 42852 21292
rect 42812 17762 42840 21286
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 43456 21010 43484 23462
rect 43444 21004 43496 21010
rect 43444 20946 43496 20952
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42984 19780 43036 19786
rect 42984 19722 43036 19728
rect 42996 19242 43024 19722
rect 43548 19394 43576 24006
rect 43640 22778 43668 26726
rect 43732 24138 43760 27406
rect 43824 27130 43852 33798
rect 43904 31408 43956 31414
rect 43904 31350 43956 31356
rect 43916 28218 43944 31350
rect 43904 28212 43956 28218
rect 43904 28154 43956 28160
rect 44192 28150 44220 34682
rect 44180 28144 44232 28150
rect 44180 28086 44232 28092
rect 44376 28082 44404 53926
rect 46204 47456 46256 47462
rect 46204 47398 46256 47404
rect 45652 31952 45704 31958
rect 45652 31894 45704 31900
rect 44364 28076 44416 28082
rect 44364 28018 44416 28024
rect 44088 28008 44140 28014
rect 44088 27950 44140 27956
rect 43904 27532 43956 27538
rect 43904 27474 43956 27480
rect 43812 27124 43864 27130
rect 43812 27066 43864 27072
rect 43824 24206 43852 27066
rect 43916 25786 43944 27474
rect 44100 26518 44128 27950
rect 45100 26920 45152 26926
rect 45100 26862 45152 26868
rect 44088 26512 44140 26518
rect 44088 26454 44140 26460
rect 44100 26330 44128 26454
rect 44100 26302 44220 26330
rect 43916 25758 44036 25786
rect 44008 25702 44036 25758
rect 43996 25696 44048 25702
rect 43996 25638 44048 25644
rect 43904 25424 43956 25430
rect 43904 25366 43956 25372
rect 43812 24200 43864 24206
rect 43812 24142 43864 24148
rect 43720 24132 43772 24138
rect 43720 24074 43772 24080
rect 43732 23050 43760 24074
rect 43720 23044 43772 23050
rect 43720 22986 43772 22992
rect 43628 22772 43680 22778
rect 43628 22714 43680 22720
rect 43824 22094 43852 24142
rect 43732 22066 43852 22094
rect 43916 22094 43944 25366
rect 44008 25158 44036 25638
rect 44192 25378 44220 26302
rect 45112 25974 45140 26862
rect 45468 26308 45520 26314
rect 45468 26250 45520 26256
rect 45100 25968 45152 25974
rect 45100 25910 45152 25916
rect 44364 25900 44416 25906
rect 44364 25842 44416 25848
rect 44088 25356 44140 25362
rect 44192 25350 44312 25378
rect 44088 25298 44140 25304
rect 43996 25152 44048 25158
rect 43996 25094 44048 25100
rect 43996 24948 44048 24954
rect 43996 24890 44048 24896
rect 44008 22710 44036 24890
rect 44100 24818 44128 25298
rect 44088 24812 44140 24818
rect 44088 24754 44140 24760
rect 44100 23798 44128 24754
rect 44088 23792 44140 23798
rect 44088 23734 44140 23740
rect 44180 23044 44232 23050
rect 44180 22986 44232 22992
rect 43996 22704 44048 22710
rect 43996 22646 44048 22652
rect 44192 22098 44220 22986
rect 43916 22066 44128 22094
rect 43732 21690 43760 22066
rect 43904 21888 43956 21894
rect 43824 21836 43904 21842
rect 43824 21830 43956 21836
rect 43824 21814 43944 21830
rect 43720 21684 43772 21690
rect 43720 21626 43772 21632
rect 43824 21622 43852 21814
rect 43996 21684 44048 21690
rect 43996 21626 44048 21632
rect 43812 21616 43864 21622
rect 43812 21558 43864 21564
rect 43628 21072 43680 21078
rect 43628 21014 43680 21020
rect 43364 19378 43576 19394
rect 43352 19372 43576 19378
rect 43404 19366 43576 19372
rect 43352 19314 43404 19320
rect 42984 19236 43036 19242
rect 42984 19178 43036 19184
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42892 18624 42944 18630
rect 42892 18566 42944 18572
rect 43352 18624 43404 18630
rect 43352 18566 43404 18572
rect 42904 18358 42932 18566
rect 42892 18352 42944 18358
rect 42892 18294 42944 18300
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 42812 17734 42932 17762
rect 42800 17672 42852 17678
rect 42800 17614 42852 17620
rect 42616 16652 42668 16658
rect 42616 16594 42668 16600
rect 42812 16522 42840 17614
rect 42904 17270 42932 17734
rect 42892 17264 42944 17270
rect 42892 17206 42944 17212
rect 43364 17134 43392 18566
rect 43444 18216 43496 18222
rect 43444 18158 43496 18164
rect 43456 17882 43484 18158
rect 43444 17876 43496 17882
rect 43444 17818 43496 17824
rect 43536 17536 43588 17542
rect 43536 17478 43588 17484
rect 43352 17128 43404 17134
rect 43352 17070 43404 17076
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 42800 16516 42852 16522
rect 42800 16458 42852 16464
rect 42708 15904 42760 15910
rect 42708 15846 42760 15852
rect 42524 15360 42576 15366
rect 42524 15302 42576 15308
rect 42432 14068 42484 14074
rect 42432 14010 42484 14016
rect 42340 13388 42392 13394
rect 42340 13330 42392 13336
rect 42444 11762 42472 14010
rect 42720 14006 42748 15846
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 43548 15026 43576 17478
rect 43640 15502 43668 21014
rect 43824 19310 43852 21558
rect 44008 21486 44036 21626
rect 43996 21480 44048 21486
rect 43996 21422 44048 21428
rect 43904 20800 43956 20806
rect 43904 20742 43956 20748
rect 43916 19854 43944 20742
rect 44008 19922 44036 21422
rect 44100 20874 44128 22066
rect 44180 22092 44232 22098
rect 44180 22034 44232 22040
rect 44088 20868 44140 20874
rect 44088 20810 44140 20816
rect 43996 19916 44048 19922
rect 43996 19858 44048 19864
rect 43904 19848 43956 19854
rect 43904 19790 43956 19796
rect 43902 19544 43958 19553
rect 43902 19479 43958 19488
rect 43916 19446 43944 19479
rect 43904 19440 43956 19446
rect 43904 19382 43956 19388
rect 43812 19304 43864 19310
rect 43812 19246 43864 19252
rect 43996 19236 44048 19242
rect 43996 19178 44048 19184
rect 44008 18698 44036 19178
rect 43996 18692 44048 18698
rect 43996 18634 44048 18640
rect 44008 18290 44036 18634
rect 43996 18284 44048 18290
rect 44048 18244 44128 18272
rect 43996 18226 44048 18232
rect 44100 17338 44128 18244
rect 44088 17332 44140 17338
rect 44088 17274 44140 17280
rect 43996 17060 44048 17066
rect 44100 17048 44128 17274
rect 44284 17270 44312 25350
rect 44376 25294 44404 25842
rect 44364 25288 44416 25294
rect 44364 25230 44416 25236
rect 44376 24886 44404 25230
rect 44364 24880 44416 24886
rect 44364 24822 44416 24828
rect 45112 24750 45140 25910
rect 45480 25294 45508 26250
rect 45664 25362 45692 31894
rect 46216 28218 46244 47398
rect 46848 33312 46900 33318
rect 46848 33254 46900 33260
rect 46204 28212 46256 28218
rect 46204 28154 46256 28160
rect 46860 27470 46888 33254
rect 46952 31686 46980 53926
rect 48424 53582 48452 56199
rect 49146 54632 49202 54641
rect 49146 54567 49202 54576
rect 49056 54188 49108 54194
rect 49056 54130 49108 54136
rect 48504 53984 48556 53990
rect 48504 53926 48556 53932
rect 48872 53984 48924 53990
rect 48872 53926 48924 53932
rect 48412 53576 48464 53582
rect 48412 53518 48464 53524
rect 48412 53440 48464 53446
rect 48412 53382 48464 53388
rect 47950 53340 48258 53349
rect 47950 53338 47956 53340
rect 48012 53338 48036 53340
rect 48092 53338 48116 53340
rect 48172 53338 48196 53340
rect 48252 53338 48258 53340
rect 48012 53286 48014 53338
rect 48194 53286 48196 53338
rect 47950 53284 47956 53286
rect 48012 53284 48036 53286
rect 48092 53284 48116 53286
rect 48172 53284 48196 53286
rect 48252 53284 48258 53286
rect 47950 53275 48258 53284
rect 47950 52252 48258 52261
rect 47950 52250 47956 52252
rect 48012 52250 48036 52252
rect 48092 52250 48116 52252
rect 48172 52250 48196 52252
rect 48252 52250 48258 52252
rect 48012 52198 48014 52250
rect 48194 52198 48196 52250
rect 47950 52196 47956 52198
rect 48012 52196 48036 52198
rect 48092 52196 48116 52198
rect 48172 52196 48196 52198
rect 48252 52196 48258 52198
rect 47950 52187 48258 52196
rect 47950 51164 48258 51173
rect 47950 51162 47956 51164
rect 48012 51162 48036 51164
rect 48092 51162 48116 51164
rect 48172 51162 48196 51164
rect 48252 51162 48258 51164
rect 48012 51110 48014 51162
rect 48194 51110 48196 51162
rect 47950 51108 47956 51110
rect 48012 51108 48036 51110
rect 48092 51108 48116 51110
rect 48172 51108 48196 51110
rect 48252 51108 48258 51110
rect 47950 51099 48258 51108
rect 47950 50076 48258 50085
rect 47950 50074 47956 50076
rect 48012 50074 48036 50076
rect 48092 50074 48116 50076
rect 48172 50074 48196 50076
rect 48252 50074 48258 50076
rect 48012 50022 48014 50074
rect 48194 50022 48196 50074
rect 47950 50020 47956 50022
rect 48012 50020 48036 50022
rect 48092 50020 48116 50022
rect 48172 50020 48196 50022
rect 48252 50020 48258 50022
rect 47950 50011 48258 50020
rect 47950 48988 48258 48997
rect 47950 48986 47956 48988
rect 48012 48986 48036 48988
rect 48092 48986 48116 48988
rect 48172 48986 48196 48988
rect 48252 48986 48258 48988
rect 48012 48934 48014 48986
rect 48194 48934 48196 48986
rect 47950 48932 47956 48934
rect 48012 48932 48036 48934
rect 48092 48932 48116 48934
rect 48172 48932 48196 48934
rect 48252 48932 48258 48934
rect 47950 48923 48258 48932
rect 47950 47900 48258 47909
rect 47950 47898 47956 47900
rect 48012 47898 48036 47900
rect 48092 47898 48116 47900
rect 48172 47898 48196 47900
rect 48252 47898 48258 47900
rect 48012 47846 48014 47898
rect 48194 47846 48196 47898
rect 47950 47844 47956 47846
rect 48012 47844 48036 47846
rect 48092 47844 48116 47846
rect 48172 47844 48196 47846
rect 48252 47844 48258 47846
rect 47950 47835 48258 47844
rect 47950 46812 48258 46821
rect 47950 46810 47956 46812
rect 48012 46810 48036 46812
rect 48092 46810 48116 46812
rect 48172 46810 48196 46812
rect 48252 46810 48258 46812
rect 48012 46758 48014 46810
rect 48194 46758 48196 46810
rect 47950 46756 47956 46758
rect 48012 46756 48036 46758
rect 48092 46756 48116 46758
rect 48172 46756 48196 46758
rect 48252 46756 48258 46758
rect 47950 46747 48258 46756
rect 47950 45724 48258 45733
rect 47950 45722 47956 45724
rect 48012 45722 48036 45724
rect 48092 45722 48116 45724
rect 48172 45722 48196 45724
rect 48252 45722 48258 45724
rect 48012 45670 48014 45722
rect 48194 45670 48196 45722
rect 47950 45668 47956 45670
rect 48012 45668 48036 45670
rect 48092 45668 48116 45670
rect 48172 45668 48196 45670
rect 48252 45668 48258 45670
rect 47950 45659 48258 45668
rect 47950 44636 48258 44645
rect 47950 44634 47956 44636
rect 48012 44634 48036 44636
rect 48092 44634 48116 44636
rect 48172 44634 48196 44636
rect 48252 44634 48258 44636
rect 48012 44582 48014 44634
rect 48194 44582 48196 44634
rect 47950 44580 47956 44582
rect 48012 44580 48036 44582
rect 48092 44580 48116 44582
rect 48172 44580 48196 44582
rect 48252 44580 48258 44582
rect 47950 44571 48258 44580
rect 47950 43548 48258 43557
rect 47950 43546 47956 43548
rect 48012 43546 48036 43548
rect 48092 43546 48116 43548
rect 48172 43546 48196 43548
rect 48252 43546 48258 43548
rect 48012 43494 48014 43546
rect 48194 43494 48196 43546
rect 47950 43492 47956 43494
rect 48012 43492 48036 43494
rect 48092 43492 48116 43494
rect 48172 43492 48196 43494
rect 48252 43492 48258 43494
rect 47950 43483 48258 43492
rect 47950 42460 48258 42469
rect 47950 42458 47956 42460
rect 48012 42458 48036 42460
rect 48092 42458 48116 42460
rect 48172 42458 48196 42460
rect 48252 42458 48258 42460
rect 48012 42406 48014 42458
rect 48194 42406 48196 42458
rect 47950 42404 47956 42406
rect 48012 42404 48036 42406
rect 48092 42404 48116 42406
rect 48172 42404 48196 42406
rect 48252 42404 48258 42406
rect 47950 42395 48258 42404
rect 47950 41372 48258 41381
rect 47950 41370 47956 41372
rect 48012 41370 48036 41372
rect 48092 41370 48116 41372
rect 48172 41370 48196 41372
rect 48252 41370 48258 41372
rect 48012 41318 48014 41370
rect 48194 41318 48196 41370
rect 47950 41316 47956 41318
rect 48012 41316 48036 41318
rect 48092 41316 48116 41318
rect 48172 41316 48196 41318
rect 48252 41316 48258 41318
rect 47950 41307 48258 41316
rect 48320 40928 48372 40934
rect 48320 40870 48372 40876
rect 47950 40284 48258 40293
rect 47950 40282 47956 40284
rect 48012 40282 48036 40284
rect 48092 40282 48116 40284
rect 48172 40282 48196 40284
rect 48252 40282 48258 40284
rect 48012 40230 48014 40282
rect 48194 40230 48196 40282
rect 47950 40228 47956 40230
rect 48012 40228 48036 40230
rect 48092 40228 48116 40230
rect 48172 40228 48196 40230
rect 48252 40228 48258 40230
rect 47950 40219 48258 40228
rect 47950 39196 48258 39205
rect 47950 39194 47956 39196
rect 48012 39194 48036 39196
rect 48092 39194 48116 39196
rect 48172 39194 48196 39196
rect 48252 39194 48258 39196
rect 48012 39142 48014 39194
rect 48194 39142 48196 39194
rect 47950 39140 47956 39142
rect 48012 39140 48036 39142
rect 48092 39140 48116 39142
rect 48172 39140 48196 39142
rect 48252 39140 48258 39142
rect 47950 39131 48258 39140
rect 47950 38108 48258 38117
rect 47950 38106 47956 38108
rect 48012 38106 48036 38108
rect 48092 38106 48116 38108
rect 48172 38106 48196 38108
rect 48252 38106 48258 38108
rect 48012 38054 48014 38106
rect 48194 38054 48196 38106
rect 47950 38052 47956 38054
rect 48012 38052 48036 38054
rect 48092 38052 48116 38054
rect 48172 38052 48196 38054
rect 48252 38052 48258 38054
rect 47950 38043 48258 38052
rect 47950 37020 48258 37029
rect 47950 37018 47956 37020
rect 48012 37018 48036 37020
rect 48092 37018 48116 37020
rect 48172 37018 48196 37020
rect 48252 37018 48258 37020
rect 48012 36966 48014 37018
rect 48194 36966 48196 37018
rect 47950 36964 47956 36966
rect 48012 36964 48036 36966
rect 48092 36964 48116 36966
rect 48172 36964 48196 36966
rect 48252 36964 48258 36966
rect 47950 36955 48258 36964
rect 47950 35932 48258 35941
rect 47950 35930 47956 35932
rect 48012 35930 48036 35932
rect 48092 35930 48116 35932
rect 48172 35930 48196 35932
rect 48252 35930 48258 35932
rect 48012 35878 48014 35930
rect 48194 35878 48196 35930
rect 47950 35876 47956 35878
rect 48012 35876 48036 35878
rect 48092 35876 48116 35878
rect 48172 35876 48196 35878
rect 48252 35876 48258 35878
rect 47950 35867 48258 35876
rect 47950 34844 48258 34853
rect 47950 34842 47956 34844
rect 48012 34842 48036 34844
rect 48092 34842 48116 34844
rect 48172 34842 48196 34844
rect 48252 34842 48258 34844
rect 48012 34790 48014 34842
rect 48194 34790 48196 34842
rect 47950 34788 47956 34790
rect 48012 34788 48036 34790
rect 48092 34788 48116 34790
rect 48172 34788 48196 34790
rect 48252 34788 48258 34790
rect 47950 34779 48258 34788
rect 47950 33756 48258 33765
rect 47950 33754 47956 33756
rect 48012 33754 48036 33756
rect 48092 33754 48116 33756
rect 48172 33754 48196 33756
rect 48252 33754 48258 33756
rect 48012 33702 48014 33754
rect 48194 33702 48196 33754
rect 47950 33700 47956 33702
rect 48012 33700 48036 33702
rect 48092 33700 48116 33702
rect 48172 33700 48196 33702
rect 48252 33700 48258 33702
rect 47950 33691 48258 33700
rect 47400 32768 47452 32774
rect 47400 32710 47452 32716
rect 46940 31680 46992 31686
rect 46940 31622 46992 31628
rect 46940 28416 46992 28422
rect 46940 28358 46992 28364
rect 46848 27464 46900 27470
rect 46848 27406 46900 27412
rect 46112 25968 46164 25974
rect 46032 25916 46112 25922
rect 46032 25910 46164 25916
rect 46032 25894 46152 25910
rect 45652 25356 45704 25362
rect 45652 25298 45704 25304
rect 45928 25356 45980 25362
rect 45928 25298 45980 25304
rect 45468 25288 45520 25294
rect 45468 25230 45520 25236
rect 45560 25152 45612 25158
rect 45558 25120 45560 25129
rect 45612 25120 45614 25129
rect 45558 25055 45614 25064
rect 45836 24812 45888 24818
rect 45836 24754 45888 24760
rect 45100 24744 45152 24750
rect 45100 24686 45152 24692
rect 45744 24268 45796 24274
rect 45744 24210 45796 24216
rect 45192 24064 45244 24070
rect 45192 24006 45244 24012
rect 44640 23724 44692 23730
rect 44640 23666 44692 23672
rect 44364 23180 44416 23186
rect 44364 23122 44416 23128
rect 44376 20058 44404 23122
rect 44652 22642 44680 23666
rect 44640 22636 44692 22642
rect 44640 22578 44692 22584
rect 44916 22636 44968 22642
rect 44916 22578 44968 22584
rect 44548 22568 44600 22574
rect 44548 22510 44600 22516
rect 44560 21894 44588 22510
rect 44928 22030 44956 22578
rect 44916 22024 44968 22030
rect 44916 21966 44968 21972
rect 44548 21888 44600 21894
rect 44548 21830 44600 21836
rect 44560 20398 44588 21830
rect 44928 21690 44956 21966
rect 44916 21684 44968 21690
rect 44916 21626 44968 21632
rect 45204 20602 45232 24006
rect 45560 22094 45612 22098
rect 45756 22094 45784 24210
rect 45848 22778 45876 24754
rect 45940 23662 45968 25298
rect 46032 24886 46060 25894
rect 46020 24880 46072 24886
rect 46020 24822 46072 24828
rect 46032 23730 46060 24822
rect 46572 24336 46624 24342
rect 46572 24278 46624 24284
rect 46584 24206 46612 24278
rect 46572 24200 46624 24206
rect 46572 24142 46624 24148
rect 46388 24064 46440 24070
rect 46388 24006 46440 24012
rect 46400 23730 46428 24006
rect 46020 23724 46072 23730
rect 46020 23666 46072 23672
rect 46388 23724 46440 23730
rect 46388 23666 46440 23672
rect 45928 23656 45980 23662
rect 45928 23598 45980 23604
rect 46032 23474 46060 23666
rect 46664 23656 46716 23662
rect 46664 23598 46716 23604
rect 45940 23446 46060 23474
rect 45836 22772 45888 22778
rect 45836 22714 45888 22720
rect 45940 22710 45968 23446
rect 46676 22778 46704 23598
rect 46952 23254 46980 28358
rect 47412 27130 47440 32710
rect 47950 32668 48258 32677
rect 47950 32666 47956 32668
rect 48012 32666 48036 32668
rect 48092 32666 48116 32668
rect 48172 32666 48196 32668
rect 48252 32666 48258 32668
rect 48012 32614 48014 32666
rect 48194 32614 48196 32666
rect 47950 32612 47956 32614
rect 48012 32612 48036 32614
rect 48092 32612 48116 32614
rect 48172 32612 48196 32614
rect 48252 32612 48258 32614
rect 47950 32603 48258 32612
rect 48332 31822 48360 40870
rect 48320 31816 48372 31822
rect 48320 31758 48372 31764
rect 47950 31580 48258 31589
rect 47950 31578 47956 31580
rect 48012 31578 48036 31580
rect 48092 31578 48116 31580
rect 48172 31578 48196 31580
rect 48252 31578 48258 31580
rect 48012 31526 48014 31578
rect 48194 31526 48196 31578
rect 47950 31524 47956 31526
rect 48012 31524 48036 31526
rect 48092 31524 48116 31526
rect 48172 31524 48196 31526
rect 48252 31524 48258 31526
rect 47950 31515 48258 31524
rect 48320 31136 48372 31142
rect 48320 31078 48372 31084
rect 47950 30492 48258 30501
rect 47950 30490 47956 30492
rect 48012 30490 48036 30492
rect 48092 30490 48116 30492
rect 48172 30490 48196 30492
rect 48252 30490 48258 30492
rect 48012 30438 48014 30490
rect 48194 30438 48196 30490
rect 47950 30436 47956 30438
rect 48012 30436 48036 30438
rect 48092 30436 48116 30438
rect 48172 30436 48196 30438
rect 48252 30436 48258 30438
rect 47950 30427 48258 30436
rect 47950 29404 48258 29413
rect 47950 29402 47956 29404
rect 48012 29402 48036 29404
rect 48092 29402 48116 29404
rect 48172 29402 48196 29404
rect 48252 29402 48258 29404
rect 48012 29350 48014 29402
rect 48194 29350 48196 29402
rect 47950 29348 47956 29350
rect 48012 29348 48036 29350
rect 48092 29348 48116 29350
rect 48172 29348 48196 29350
rect 48252 29348 48258 29350
rect 47950 29339 48258 29348
rect 47950 28316 48258 28325
rect 47950 28314 47956 28316
rect 48012 28314 48036 28316
rect 48092 28314 48116 28316
rect 48172 28314 48196 28316
rect 48252 28314 48258 28316
rect 48012 28262 48014 28314
rect 48194 28262 48196 28314
rect 47950 28260 47956 28262
rect 48012 28260 48036 28262
rect 48092 28260 48116 28262
rect 48172 28260 48196 28262
rect 48252 28260 48258 28262
rect 47950 28251 48258 28260
rect 47950 27228 48258 27237
rect 47950 27226 47956 27228
rect 48012 27226 48036 27228
rect 48092 27226 48116 27228
rect 48172 27226 48196 27228
rect 48252 27226 48258 27228
rect 48012 27174 48014 27226
rect 48194 27174 48196 27226
rect 47950 27172 47956 27174
rect 48012 27172 48036 27174
rect 48092 27172 48116 27174
rect 48172 27172 48196 27174
rect 48252 27172 48258 27174
rect 47950 27163 48258 27172
rect 47400 27124 47452 27130
rect 47400 27066 47452 27072
rect 47032 26784 47084 26790
rect 47032 26726 47084 26732
rect 46940 23248 46992 23254
rect 46940 23190 46992 23196
rect 46756 23044 46808 23050
rect 46756 22986 46808 22992
rect 46664 22772 46716 22778
rect 46664 22714 46716 22720
rect 45928 22704 45980 22710
rect 45928 22646 45980 22652
rect 45560 22092 45784 22094
rect 45612 22066 45784 22092
rect 45560 22034 45612 22040
rect 45572 22003 45600 22034
rect 45756 21690 45784 22066
rect 45940 21962 45968 22646
rect 46768 22030 46796 22986
rect 47044 22438 47072 26726
rect 47950 26140 48258 26149
rect 47950 26138 47956 26140
rect 48012 26138 48036 26140
rect 48092 26138 48116 26140
rect 48172 26138 48196 26140
rect 48252 26138 48258 26140
rect 48012 26086 48014 26138
rect 48194 26086 48196 26138
rect 47950 26084 47956 26086
rect 48012 26084 48036 26086
rect 48092 26084 48116 26086
rect 48172 26084 48196 26086
rect 48252 26084 48258 26086
rect 47950 26075 48258 26084
rect 47950 25052 48258 25061
rect 47950 25050 47956 25052
rect 48012 25050 48036 25052
rect 48092 25050 48116 25052
rect 48172 25050 48196 25052
rect 48252 25050 48258 25052
rect 48012 24998 48014 25050
rect 48194 24998 48196 25050
rect 47950 24996 47956 24998
rect 48012 24996 48036 24998
rect 48092 24996 48116 24998
rect 48172 24996 48196 24998
rect 48252 24996 48258 24998
rect 47950 24987 48258 24996
rect 48332 24138 48360 31078
rect 48424 29646 48452 53382
rect 48412 29640 48464 29646
rect 48412 29582 48464 29588
rect 48412 29504 48464 29510
rect 48412 29446 48464 29452
rect 48424 24614 48452 29446
rect 48516 29102 48544 53926
rect 48688 44736 48740 44742
rect 48688 44678 48740 44684
rect 48596 39296 48648 39302
rect 48596 39238 48648 39244
rect 48608 30598 48636 39238
rect 48700 33658 48728 44678
rect 48780 36576 48832 36582
rect 48780 36518 48832 36524
rect 48688 33652 48740 33658
rect 48688 33594 48740 33600
rect 48596 30592 48648 30598
rect 48596 30534 48648 30540
rect 48688 30048 48740 30054
rect 48688 29990 48740 29996
rect 48504 29096 48556 29102
rect 48504 29038 48556 29044
rect 48504 26376 48556 26382
rect 48504 26318 48556 26324
rect 48596 26376 48648 26382
rect 48596 26318 48648 26324
rect 48516 26081 48544 26318
rect 48502 26072 48558 26081
rect 48502 26007 48558 26016
rect 48412 24608 48464 24614
rect 48412 24550 48464 24556
rect 48320 24132 48372 24138
rect 48320 24074 48372 24080
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47032 22432 47084 22438
rect 47032 22374 47084 22380
rect 46756 22024 46808 22030
rect 46756 21966 46808 21972
rect 45928 21956 45980 21962
rect 45928 21898 45980 21904
rect 45744 21684 45796 21690
rect 45744 21626 45796 21632
rect 45940 21622 45968 21898
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 45928 21616 45980 21622
rect 45928 21558 45980 21564
rect 47032 21548 47084 21554
rect 47032 21490 47084 21496
rect 45192 20596 45244 20602
rect 45192 20538 45244 20544
rect 47044 20534 47072 21490
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47032 20528 47084 20534
rect 47032 20470 47084 20476
rect 46940 20460 46992 20466
rect 46940 20402 46992 20408
rect 44548 20392 44600 20398
rect 44548 20334 44600 20340
rect 44364 20052 44416 20058
rect 44364 19994 44416 20000
rect 44376 18426 44404 19994
rect 46952 19310 46980 20402
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47952 19508 48004 19514
rect 47952 19450 48004 19456
rect 46940 19304 46992 19310
rect 46940 19246 46992 19252
rect 47964 18766 47992 19450
rect 47952 18760 48004 18766
rect 47952 18702 48004 18708
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 44364 18420 44416 18426
rect 44364 18362 44416 18368
rect 44548 17604 44600 17610
rect 44548 17546 44600 17552
rect 45468 17604 45520 17610
rect 45468 17546 45520 17552
rect 44272 17264 44324 17270
rect 44272 17206 44324 17212
rect 44048 17020 44128 17048
rect 43996 17002 44048 17008
rect 44456 16584 44508 16590
rect 44456 16526 44508 16532
rect 43628 15496 43680 15502
rect 43628 15438 43680 15444
rect 43536 15020 43588 15026
rect 43536 14962 43588 14968
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 44468 14074 44496 16526
rect 44456 14068 44508 14074
rect 44456 14010 44508 14016
rect 42708 14000 42760 14006
rect 42708 13942 42760 13948
rect 43352 13932 43404 13938
rect 43352 13874 43404 13880
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 43364 12170 43392 13874
rect 44364 13320 44416 13326
rect 44364 13262 44416 13268
rect 44180 12640 44232 12646
rect 44180 12582 44232 12588
rect 43352 12164 43404 12170
rect 43352 12106 43404 12112
rect 42432 11756 42484 11762
rect 42432 11698 42484 11704
rect 43720 11688 43772 11694
rect 43720 11630 43772 11636
rect 42800 11620 42852 11626
rect 42800 11562 42852 11568
rect 42812 10674 42840 11562
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 42800 10668 42852 10674
rect 42800 10610 42852 10616
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 43732 9586 43760 11630
rect 44088 10464 44140 10470
rect 44088 10406 44140 10412
rect 44100 9586 44128 10406
rect 44192 9994 44220 12582
rect 44376 11354 44404 13262
rect 44364 11348 44416 11354
rect 44364 11290 44416 11296
rect 44180 9988 44232 9994
rect 44180 9930 44232 9936
rect 43720 9580 43772 9586
rect 43720 9522 43772 9528
rect 44088 9580 44140 9586
rect 44088 9522 44140 9528
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 44180 8968 44232 8974
rect 44180 8910 44232 8916
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 44192 8090 44220 8910
rect 44180 8084 44232 8090
rect 44180 8026 44232 8032
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 44088 6656 44140 6662
rect 44088 6598 44140 6604
rect 42616 6112 42668 6118
rect 42616 6054 42668 6060
rect 42628 3058 42656 6054
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 43352 5840 43404 5846
rect 43352 5782 43404 5788
rect 42800 5636 42852 5642
rect 42800 5578 42852 5584
rect 42708 5092 42760 5098
rect 42708 5034 42760 5040
rect 42720 3534 42748 5034
rect 42812 4146 42840 5578
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 42800 4140 42852 4146
rect 42800 4082 42852 4088
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43364 3058 43392 5782
rect 44100 5234 44128 6598
rect 44088 5228 44140 5234
rect 44088 5170 44140 5176
rect 44180 4072 44232 4078
rect 44180 4014 44232 4020
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 41972 2984 42024 2990
rect 41972 2926 42024 2932
rect 41616 2746 41736 2774
rect 41616 2038 41644 2746
rect 41604 2032 41656 2038
rect 41604 1974 41656 1980
rect 41984 800 42012 2926
rect 42708 2916 42760 2922
rect 42708 2858 42760 2864
rect 42720 800 42748 2858
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 43444 2508 43496 2514
rect 43444 2450 43496 2456
rect 43456 800 43484 2450
rect 44192 800 44220 4014
rect 44560 3126 44588 17546
rect 44732 15496 44784 15502
rect 44732 15438 44784 15444
rect 44640 13456 44692 13462
rect 44640 13398 44692 13404
rect 44652 10062 44680 13398
rect 44744 13394 44772 15438
rect 44732 13388 44784 13394
rect 44732 13330 44784 13336
rect 45480 12434 45508 17546
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 45560 17196 45612 17202
rect 45560 17138 45612 17144
rect 45572 15638 45600 17138
rect 46112 16992 46164 16998
rect 46112 16934 46164 16940
rect 46124 16658 46152 16934
rect 46112 16652 46164 16658
rect 46112 16594 46164 16600
rect 45560 15632 45612 15638
rect 45560 15574 45612 15580
rect 45928 13864 45980 13870
rect 45928 13806 45980 13812
rect 45388 12406 45508 12434
rect 45192 11552 45244 11558
rect 45192 11494 45244 11500
rect 44640 10056 44692 10062
rect 44640 9998 44692 10004
rect 45204 8566 45232 11494
rect 45284 8900 45336 8906
rect 45284 8842 45336 8848
rect 45192 8560 45244 8566
rect 45192 8502 45244 8508
rect 45296 8022 45324 8842
rect 45284 8016 45336 8022
rect 45284 7958 45336 7964
rect 45192 6316 45244 6322
rect 45192 6258 45244 6264
rect 45204 5914 45232 6258
rect 45192 5908 45244 5914
rect 45192 5850 45244 5856
rect 44916 3596 44968 3602
rect 44916 3538 44968 3544
rect 44548 3120 44600 3126
rect 44548 3062 44600 3068
rect 44928 800 44956 3538
rect 45388 2650 45416 12406
rect 45940 12238 45968 13806
rect 45928 12232 45980 12238
rect 45928 12174 45980 12180
rect 45560 10668 45612 10674
rect 45560 10610 45612 10616
rect 45468 9376 45520 9382
rect 45468 9318 45520 9324
rect 45480 7410 45508 9318
rect 45572 9178 45600 10610
rect 45560 9172 45612 9178
rect 45560 9114 45612 9120
rect 45468 7404 45520 7410
rect 45468 7346 45520 7352
rect 45468 7200 45520 7206
rect 45468 7142 45520 7148
rect 45480 5710 45508 7142
rect 45468 5704 45520 5710
rect 45468 5646 45520 5652
rect 45468 5568 45520 5574
rect 45468 5510 45520 5516
rect 45480 4146 45508 5510
rect 46124 4622 46152 16594
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47768 15428 47820 15434
rect 47768 15370 47820 15376
rect 47780 13938 47808 15370
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47952 15020 48004 15026
rect 47952 14962 48004 14968
rect 47860 14816 47912 14822
rect 47860 14758 47912 14764
rect 47768 13932 47820 13938
rect 47768 13874 47820 13880
rect 47872 13326 47900 14758
rect 47964 14618 47992 14962
rect 47952 14612 48004 14618
rect 47952 14554 48004 14560
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47860 13320 47912 13326
rect 47860 13262 47912 13268
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 48608 12986 48636 26318
rect 48700 24274 48728 29990
rect 48688 24268 48740 24274
rect 48688 24210 48740 24216
rect 48792 13530 48820 36518
rect 48884 29782 48912 53926
rect 49068 53825 49096 54130
rect 49054 53816 49110 53825
rect 49054 53751 49110 53760
rect 49160 53582 49188 54567
rect 49436 53650 49464 56200
rect 49424 53644 49476 53650
rect 49424 53586 49476 53592
rect 49148 53576 49200 53582
rect 49148 53518 49200 53524
rect 50160 53440 50212 53446
rect 50160 53382 50212 53388
rect 49056 53100 49108 53106
rect 49056 53042 49108 53048
rect 49068 53009 49096 53042
rect 49054 53000 49110 53009
rect 49054 52935 49110 52944
rect 49976 52488 50028 52494
rect 49976 52430 50028 52436
rect 48964 52420 49016 52426
rect 48964 52362 49016 52368
rect 48976 52193 49004 52362
rect 48962 52184 49018 52193
rect 48962 52119 49018 52128
rect 48962 51368 49018 51377
rect 48962 51303 48964 51312
rect 49016 51303 49018 51312
rect 49608 51332 49660 51338
rect 48964 51274 49016 51280
rect 49608 51274 49660 51280
rect 48964 50924 49016 50930
rect 48964 50866 49016 50872
rect 48976 50561 49004 50866
rect 48962 50552 49018 50561
rect 48962 50487 49018 50496
rect 49148 49836 49200 49842
rect 49148 49778 49200 49784
rect 49160 49745 49188 49778
rect 49516 49768 49568 49774
rect 49146 49736 49202 49745
rect 49516 49710 49568 49716
rect 49146 49671 49202 49680
rect 49148 49156 49200 49162
rect 49148 49098 49200 49104
rect 49160 48929 49188 49098
rect 49146 48920 49202 48929
rect 49146 48855 49202 48864
rect 49146 48104 49202 48113
rect 49146 48039 49148 48048
rect 49200 48039 49202 48048
rect 49148 48010 49200 48016
rect 49332 47660 49384 47666
rect 49332 47602 49384 47608
rect 49344 47297 49372 47602
rect 49330 47288 49386 47297
rect 49330 47223 49386 47232
rect 49332 46572 49384 46578
rect 49332 46514 49384 46520
rect 49344 46481 49372 46514
rect 49330 46472 49386 46481
rect 49330 46407 49386 46416
rect 49332 45960 49384 45966
rect 49332 45902 49384 45908
rect 49344 45665 49372 45902
rect 49330 45656 49386 45665
rect 49330 45591 49386 45600
rect 49332 44872 49384 44878
rect 49330 44840 49332 44849
rect 49384 44840 49386 44849
rect 49330 44775 49386 44784
rect 49148 44396 49200 44402
rect 49148 44338 49200 44344
rect 49160 44033 49188 44338
rect 49146 44024 49202 44033
rect 49146 43959 49202 43968
rect 49148 43308 49200 43314
rect 49148 43250 49200 43256
rect 49160 43217 49188 43250
rect 49146 43208 49202 43217
rect 49146 43143 49202 43152
rect 49148 42628 49200 42634
rect 49148 42570 49200 42576
rect 49160 42401 49188 42570
rect 49240 42560 49292 42566
rect 49240 42502 49292 42508
rect 49146 42392 49202 42401
rect 49146 42327 49202 42336
rect 49146 41576 49202 41585
rect 49146 41511 49148 41520
rect 49200 41511 49202 41520
rect 49148 41482 49200 41488
rect 49056 40180 49108 40186
rect 49056 40122 49108 40128
rect 48964 38208 49016 38214
rect 48964 38150 49016 38156
rect 48976 29850 49004 38150
rect 49068 31482 49096 40122
rect 49148 37868 49200 37874
rect 49148 37810 49200 37816
rect 49160 37505 49188 37810
rect 49146 37496 49202 37505
rect 49146 37431 49202 37440
rect 49148 36780 49200 36786
rect 49148 36722 49200 36728
rect 49160 36689 49188 36722
rect 49146 36680 49202 36689
rect 49146 36615 49202 36624
rect 49056 31476 49108 31482
rect 49056 31418 49108 31424
rect 48964 29844 49016 29850
rect 48964 29786 49016 29792
rect 48872 29776 48924 29782
rect 48872 29718 48924 29724
rect 48872 27872 48924 27878
rect 48872 27814 48924 27820
rect 48884 21486 48912 27814
rect 49148 25288 49200 25294
rect 49146 25256 49148 25265
rect 49200 25256 49202 25265
rect 49146 25191 49202 25200
rect 49148 24744 49200 24750
rect 49148 24686 49200 24692
rect 49160 24449 49188 24686
rect 49146 24440 49202 24449
rect 49146 24375 49202 24384
rect 49148 23656 49200 23662
rect 49146 23624 49148 23633
rect 49200 23624 49202 23633
rect 49146 23559 49202 23568
rect 49148 23044 49200 23050
rect 49148 22986 49200 22992
rect 49160 22817 49188 22986
rect 49146 22808 49202 22817
rect 49146 22743 49202 22752
rect 49148 22024 49200 22030
rect 49146 21992 49148 22001
rect 49200 21992 49202 22001
rect 49146 21927 49202 21936
rect 48872 21480 48924 21486
rect 48872 21422 48924 21428
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21185 49188 21422
rect 49146 21176 49202 21185
rect 49146 21111 49202 21120
rect 49148 20392 49200 20398
rect 49146 20360 49148 20369
rect 49200 20360 49202 20369
rect 49146 20295 49202 20304
rect 49148 19780 49200 19786
rect 49148 19722 49200 19728
rect 49160 19553 49188 19722
rect 49146 19544 49202 19553
rect 49146 19479 49202 19488
rect 49148 18760 49200 18766
rect 49146 18728 49148 18737
rect 49200 18728 49202 18737
rect 49146 18663 49202 18672
rect 49148 18216 49200 18222
rect 49148 18158 49200 18164
rect 49160 17921 49188 18158
rect 49146 17912 49202 17921
rect 49146 17847 49202 17856
rect 49148 17128 49200 17134
rect 49146 17096 49148 17105
rect 49200 17096 49202 17105
rect 49146 17031 49202 17040
rect 49148 16516 49200 16522
rect 49148 16458 49200 16464
rect 49160 16289 49188 16458
rect 49146 16280 49202 16289
rect 49146 16215 49202 16224
rect 49148 15496 49200 15502
rect 49146 15464 49148 15473
rect 49200 15464 49202 15473
rect 49146 15399 49202 15408
rect 49148 14952 49200 14958
rect 49148 14894 49200 14900
rect 49160 14657 49188 14894
rect 49146 14648 49202 14657
rect 49146 14583 49202 14592
rect 49252 14550 49280 42502
rect 49332 41132 49384 41138
rect 49332 41074 49384 41080
rect 49344 40769 49372 41074
rect 49330 40760 49386 40769
rect 49330 40695 49386 40704
rect 49332 40044 49384 40050
rect 49332 39986 49384 39992
rect 49344 39953 49372 39986
rect 49330 39944 49386 39953
rect 49330 39879 49386 39888
rect 49332 39432 49384 39438
rect 49332 39374 49384 39380
rect 49344 39137 49372 39374
rect 49330 39128 49386 39137
rect 49330 39063 49386 39072
rect 49332 38344 49384 38350
rect 49330 38312 49332 38321
rect 49384 38312 49386 38321
rect 49330 38247 49386 38256
rect 49424 36576 49476 36582
rect 49424 36518 49476 36524
rect 49332 36168 49384 36174
rect 49332 36110 49384 36116
rect 49344 35873 49372 36110
rect 49330 35864 49386 35873
rect 49330 35799 49386 35808
rect 49332 35080 49384 35086
rect 49330 35048 49332 35057
rect 49384 35048 49386 35057
rect 49330 34983 49386 34992
rect 49332 34604 49384 34610
rect 49332 34546 49384 34552
rect 49344 34241 49372 34546
rect 49330 34232 49386 34241
rect 49330 34167 49386 34176
rect 49332 33516 49384 33522
rect 49332 33458 49384 33464
rect 49344 33425 49372 33458
rect 49330 33416 49386 33425
rect 49330 33351 49386 33360
rect 49332 32904 49384 32910
rect 49332 32846 49384 32852
rect 49344 32609 49372 32846
rect 49330 32600 49386 32609
rect 49330 32535 49386 32544
rect 49332 31816 49384 31822
rect 49330 31784 49332 31793
rect 49384 31784 49386 31793
rect 49330 31719 49386 31728
rect 49332 31340 49384 31346
rect 49332 31282 49384 31288
rect 49344 30977 49372 31282
rect 49330 30968 49386 30977
rect 49330 30903 49386 30912
rect 49332 30252 49384 30258
rect 49332 30194 49384 30200
rect 49344 30161 49372 30194
rect 49330 30152 49386 30161
rect 49330 30087 49386 30096
rect 49332 29640 49384 29646
rect 49332 29582 49384 29588
rect 49344 29345 49372 29582
rect 49330 29336 49386 29345
rect 49330 29271 49386 29280
rect 49332 28552 49384 28558
rect 49330 28520 49332 28529
rect 49384 28520 49386 28529
rect 49330 28455 49386 28464
rect 49332 28076 49384 28082
rect 49332 28018 49384 28024
rect 49344 27713 49372 28018
rect 49330 27704 49386 27713
rect 49330 27639 49386 27648
rect 49332 26988 49384 26994
rect 49332 26930 49384 26936
rect 49344 26897 49372 26930
rect 49330 26888 49386 26897
rect 49330 26823 49386 26832
rect 49436 17542 49464 36518
rect 49528 24410 49556 49710
rect 49620 27946 49648 51274
rect 49884 45824 49936 45830
rect 49884 45766 49936 45772
rect 49700 44260 49752 44266
rect 49700 44202 49752 44208
rect 49712 36582 49740 44202
rect 49792 43172 49844 43178
rect 49792 43114 49844 43120
rect 49700 36576 49752 36582
rect 49700 36518 49752 36524
rect 49700 36032 49752 36038
rect 49700 35974 49752 35980
rect 49608 27940 49660 27946
rect 49608 27882 49660 27888
rect 49516 24404 49568 24410
rect 49516 24346 49568 24352
rect 49712 17746 49740 35974
rect 49804 17814 49832 43114
rect 49896 34066 49924 45766
rect 49884 34060 49936 34066
rect 49884 34002 49936 34008
rect 49988 29617 50016 52430
rect 50068 34944 50120 34950
rect 50068 34886 50120 34892
rect 49974 29608 50030 29617
rect 49974 29543 50030 29552
rect 49792 17808 49844 17814
rect 49792 17750 49844 17756
rect 49700 17740 49752 17746
rect 49700 17682 49752 17688
rect 50080 17678 50108 34886
rect 50172 29578 50200 53382
rect 50436 49156 50488 49162
rect 50436 49098 50488 49104
rect 50160 29572 50212 29578
rect 50160 29514 50212 29520
rect 50448 25809 50476 49098
rect 50528 37732 50580 37738
rect 50528 37674 50580 37680
rect 50434 25800 50490 25809
rect 50434 25735 50490 25744
rect 50068 17672 50120 17678
rect 50068 17614 50120 17620
rect 49424 17536 49476 17542
rect 49424 17478 49476 17484
rect 49240 14544 49292 14550
rect 49240 14486 49292 14492
rect 50540 14482 50568 37674
rect 50528 14476 50580 14482
rect 50528 14418 50580 14424
rect 49148 13864 49200 13870
rect 49146 13832 49148 13841
rect 49200 13832 49202 13841
rect 49146 13767 49202 13776
rect 48780 13524 48832 13530
rect 48780 13466 48832 13472
rect 49148 13252 49200 13258
rect 49148 13194 49200 13200
rect 49160 13025 49188 13194
rect 49146 13016 49202 13025
rect 48596 12980 48648 12986
rect 49146 12951 49202 12960
rect 48596 12922 48648 12928
rect 49148 12232 49200 12238
rect 49146 12200 49148 12209
rect 49200 12200 49202 12209
rect 49146 12135 49202 12144
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 49148 11688 49200 11694
rect 49148 11630 49200 11636
rect 49160 11393 49188 11630
rect 49146 11384 49202 11393
rect 49146 11319 49202 11328
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 49148 10600 49200 10606
rect 49146 10568 49148 10577
rect 49200 10568 49202 10577
rect 49146 10503 49202 10512
rect 46940 10056 46992 10062
rect 46940 9998 46992 10004
rect 46296 9988 46348 9994
rect 46296 9930 46348 9936
rect 46308 7478 46336 9930
rect 46952 9178 46980 9998
rect 47032 9988 47084 9994
rect 47032 9930 47084 9936
rect 49148 9988 49200 9994
rect 49148 9930 49200 9936
rect 46940 9172 46992 9178
rect 46940 9114 46992 9120
rect 46848 8356 46900 8362
rect 46848 8298 46900 8304
rect 46296 7472 46348 7478
rect 46296 7414 46348 7420
rect 46860 5846 46888 8298
rect 46940 7200 46992 7206
rect 46940 7142 46992 7148
rect 46848 5840 46900 5846
rect 46848 5782 46900 5788
rect 46952 5234 46980 7142
rect 47044 6798 47072 9930
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 49160 9761 49188 9930
rect 49146 9752 49202 9761
rect 49146 9687 49202 9696
rect 47860 9376 47912 9382
rect 47860 9318 47912 9324
rect 47872 8498 47900 9318
rect 49146 8936 49202 8945
rect 49146 8871 49148 8880
rect 49200 8871 49202 8880
rect 49148 8842 49200 8848
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 47860 8492 47912 8498
rect 47860 8434 47912 8440
rect 49148 8424 49200 8430
rect 49148 8366 49200 8372
rect 49160 8129 49188 8366
rect 49146 8120 49202 8129
rect 49146 8055 49202 8064
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 49148 7336 49200 7342
rect 49146 7304 49148 7313
rect 49200 7304 49202 7313
rect 49146 7239 49202 7248
rect 47032 6792 47084 6798
rect 47032 6734 47084 6740
rect 49148 6724 49200 6730
rect 49148 6666 49200 6672
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 49160 6497 49188 6666
rect 49146 6488 49202 6497
rect 49146 6423 49202 6432
rect 48504 6248 48556 6254
rect 48504 6190 48556 6196
rect 49240 6248 49292 6254
rect 49240 6190 49292 6196
rect 47032 5636 47084 5642
rect 47032 5578 47084 5584
rect 46940 5228 46992 5234
rect 46940 5170 46992 5176
rect 46388 4820 46440 4826
rect 46388 4762 46440 4768
rect 46112 4616 46164 4622
rect 46112 4558 46164 4564
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3058 46336 3878
rect 46296 3052 46348 3058
rect 46296 2994 46348 3000
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 45376 2644 45428 2650
rect 45376 2586 45428 2592
rect 45664 800 45692 2790
rect 46400 800 46428 4762
rect 47044 4146 47072 5578
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 47768 5160 47820 5166
rect 47768 5102 47820 5108
rect 47032 4140 47084 4146
rect 47032 4082 47084 4088
rect 47124 3460 47176 3466
rect 47124 3402 47176 3408
rect 47136 800 47164 3402
rect 47780 2446 47808 5102
rect 47952 5024 48004 5030
rect 47952 4966 48004 4972
rect 47860 4684 47912 4690
rect 47860 4626 47912 4632
rect 47768 2440 47820 2446
rect 47872 2417 47900 4626
rect 47964 4622 47992 4966
rect 47952 4616 48004 4622
rect 47952 4558 48004 4564
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 48516 3738 48544 6190
rect 49146 5672 49202 5681
rect 49146 5607 49148 5616
rect 49200 5607 49202 5616
rect 49148 5578 49200 5584
rect 49148 5160 49200 5166
rect 49148 5102 49200 5108
rect 49160 4865 49188 5102
rect 49146 4856 49202 4865
rect 49146 4791 49202 4800
rect 48688 4548 48740 4554
rect 48688 4490 48740 4496
rect 48504 3732 48556 3738
rect 48504 3674 48556 3680
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48320 2848 48372 2854
rect 48320 2790 48372 2796
rect 48332 2514 48360 2790
rect 48320 2508 48372 2514
rect 48320 2450 48372 2456
rect 47768 2382 47820 2388
rect 47858 2408 47914 2417
rect 47858 2343 47914 2352
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 28092 734 28396 762
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 30930 0 30986 800
rect 31666 0 31722 800
rect 32402 0 32458 800
rect 33138 0 33194 800
rect 33874 0 33930 800
rect 34610 0 34666 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37554 0 37610 800
rect 38290 0 38346 800
rect 39026 0 39082 800
rect 39762 0 39818 800
rect 40498 0 40554 800
rect 41234 0 41290 800
rect 41970 0 42026 800
rect 42706 0 42762 800
rect 43442 0 43498 800
rect 44178 0 44234 800
rect 44914 0 44970 800
rect 45650 0 45706 800
rect 46386 0 46442 800
rect 47122 0 47178 800
rect 47858 0 47914 800
rect 48594 0 48650 800
rect 48700 785 48728 4490
rect 49148 4072 49200 4078
rect 49146 4040 49148 4049
rect 49200 4040 49202 4049
rect 49146 3975 49202 3984
rect 49146 3224 49202 3233
rect 49146 3159 49202 3168
rect 49160 3126 49188 3159
rect 49148 3120 49200 3126
rect 49148 3062 49200 3068
rect 49252 1601 49280 6190
rect 49238 1592 49294 1601
rect 49238 1527 49294 1536
rect 48686 776 48742 785
rect 48686 711 48742 720
<< via2 >>
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 27956 54426 28012 54428
rect 28036 54426 28092 54428
rect 28116 54426 28172 54428
rect 28196 54426 28252 54428
rect 27956 54374 28002 54426
rect 28002 54374 28012 54426
rect 28036 54374 28066 54426
rect 28066 54374 28078 54426
rect 28078 54374 28092 54426
rect 28116 54374 28130 54426
rect 28130 54374 28142 54426
rect 28142 54374 28172 54426
rect 28196 54374 28206 54426
rect 28206 54374 28252 54426
rect 27956 54372 28012 54374
rect 28036 54372 28092 54374
rect 28116 54372 28172 54374
rect 28196 54372 28252 54374
rect 48410 56208 48466 56264
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 27956 53338 28012 53340
rect 28036 53338 28092 53340
rect 28116 53338 28172 53340
rect 28196 53338 28252 53340
rect 27956 53286 28002 53338
rect 28002 53286 28012 53338
rect 28036 53286 28066 53338
rect 28066 53286 28078 53338
rect 28078 53286 28092 53338
rect 28116 53286 28130 53338
rect 28130 53286 28142 53338
rect 28142 53286 28172 53338
rect 28196 53286 28206 53338
rect 28206 53286 28252 53338
rect 27956 53284 28012 53286
rect 28036 53284 28092 53286
rect 28116 53284 28172 53286
rect 28196 53284 28252 53286
rect 27956 52250 28012 52252
rect 28036 52250 28092 52252
rect 28116 52250 28172 52252
rect 28196 52250 28252 52252
rect 27956 52198 28002 52250
rect 28002 52198 28012 52250
rect 28036 52198 28066 52250
rect 28066 52198 28078 52250
rect 28078 52198 28092 52250
rect 28116 52198 28130 52250
rect 28130 52198 28142 52250
rect 28142 52198 28172 52250
rect 28196 52198 28206 52250
rect 28206 52198 28252 52250
rect 27956 52196 28012 52198
rect 28036 52196 28092 52198
rect 28116 52196 28172 52198
rect 28196 52196 28252 52198
rect 27956 51162 28012 51164
rect 28036 51162 28092 51164
rect 28116 51162 28172 51164
rect 28196 51162 28252 51164
rect 27956 51110 28002 51162
rect 28002 51110 28012 51162
rect 28036 51110 28066 51162
rect 28066 51110 28078 51162
rect 28078 51110 28092 51162
rect 28116 51110 28130 51162
rect 28130 51110 28142 51162
rect 28142 51110 28172 51162
rect 28196 51110 28206 51162
rect 28206 51110 28252 51162
rect 27956 51108 28012 51110
rect 28036 51108 28092 51110
rect 28116 51108 28172 51110
rect 28196 51108 28252 51110
rect 27956 50074 28012 50076
rect 28036 50074 28092 50076
rect 28116 50074 28172 50076
rect 28196 50074 28252 50076
rect 27956 50022 28002 50074
rect 28002 50022 28012 50074
rect 28036 50022 28066 50074
rect 28066 50022 28078 50074
rect 28078 50022 28092 50074
rect 28116 50022 28130 50074
rect 28130 50022 28142 50074
rect 28142 50022 28172 50074
rect 28196 50022 28206 50074
rect 28206 50022 28252 50074
rect 27956 50020 28012 50022
rect 28036 50020 28092 50022
rect 28116 50020 28172 50022
rect 28196 50020 28252 50022
rect 27956 48986 28012 48988
rect 28036 48986 28092 48988
rect 28116 48986 28172 48988
rect 28196 48986 28252 48988
rect 27956 48934 28002 48986
rect 28002 48934 28012 48986
rect 28036 48934 28066 48986
rect 28066 48934 28078 48986
rect 28078 48934 28092 48986
rect 28116 48934 28130 48986
rect 28130 48934 28142 48986
rect 28142 48934 28172 48986
rect 28196 48934 28206 48986
rect 28206 48934 28252 48986
rect 27956 48932 28012 48934
rect 28036 48932 28092 48934
rect 28116 48932 28172 48934
rect 28196 48932 28252 48934
rect 27956 47898 28012 47900
rect 28036 47898 28092 47900
rect 28116 47898 28172 47900
rect 28196 47898 28252 47900
rect 27956 47846 28002 47898
rect 28002 47846 28012 47898
rect 28036 47846 28066 47898
rect 28066 47846 28078 47898
rect 28078 47846 28092 47898
rect 28116 47846 28130 47898
rect 28130 47846 28142 47898
rect 28142 47846 28172 47898
rect 28196 47846 28206 47898
rect 28206 47846 28252 47898
rect 27956 47844 28012 47846
rect 28036 47844 28092 47846
rect 28116 47844 28172 47846
rect 28196 47844 28252 47846
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 27956 46810 28012 46812
rect 28036 46810 28092 46812
rect 28116 46810 28172 46812
rect 28196 46810 28252 46812
rect 27956 46758 28002 46810
rect 28002 46758 28012 46810
rect 28036 46758 28066 46810
rect 28066 46758 28078 46810
rect 28078 46758 28092 46810
rect 28116 46758 28130 46810
rect 28130 46758 28142 46810
rect 28142 46758 28172 46810
rect 28196 46758 28206 46810
rect 28206 46758 28252 46810
rect 27956 46756 28012 46758
rect 28036 46756 28092 46758
rect 28116 46756 28172 46758
rect 28196 46756 28252 46758
rect 27956 45722 28012 45724
rect 28036 45722 28092 45724
rect 28116 45722 28172 45724
rect 28196 45722 28252 45724
rect 27956 45670 28002 45722
rect 28002 45670 28012 45722
rect 28036 45670 28066 45722
rect 28066 45670 28078 45722
rect 28078 45670 28092 45722
rect 28116 45670 28130 45722
rect 28130 45670 28142 45722
rect 28142 45670 28172 45722
rect 28196 45670 28206 45722
rect 28206 45670 28252 45722
rect 27956 45668 28012 45670
rect 28036 45668 28092 45670
rect 28116 45668 28172 45670
rect 28196 45668 28252 45670
rect 27956 44634 28012 44636
rect 28036 44634 28092 44636
rect 28116 44634 28172 44636
rect 28196 44634 28252 44636
rect 27956 44582 28002 44634
rect 28002 44582 28012 44634
rect 28036 44582 28066 44634
rect 28066 44582 28078 44634
rect 28078 44582 28092 44634
rect 28116 44582 28130 44634
rect 28130 44582 28142 44634
rect 28142 44582 28172 44634
rect 28196 44582 28206 44634
rect 28206 44582 28252 44634
rect 27956 44580 28012 44582
rect 28036 44580 28092 44582
rect 28116 44580 28172 44582
rect 28196 44580 28252 44582
rect 27956 43546 28012 43548
rect 28036 43546 28092 43548
rect 28116 43546 28172 43548
rect 28196 43546 28252 43548
rect 27956 43494 28002 43546
rect 28002 43494 28012 43546
rect 28036 43494 28066 43546
rect 28066 43494 28078 43546
rect 28078 43494 28092 43546
rect 28116 43494 28130 43546
rect 28130 43494 28142 43546
rect 28142 43494 28172 43546
rect 28196 43494 28206 43546
rect 28206 43494 28252 43546
rect 27956 43492 28012 43494
rect 28036 43492 28092 43494
rect 28116 43492 28172 43494
rect 28196 43492 28252 43494
rect 27956 42458 28012 42460
rect 28036 42458 28092 42460
rect 28116 42458 28172 42460
rect 28196 42458 28252 42460
rect 27956 42406 28002 42458
rect 28002 42406 28012 42458
rect 28036 42406 28066 42458
rect 28066 42406 28078 42458
rect 28078 42406 28092 42458
rect 28116 42406 28130 42458
rect 28130 42406 28142 42458
rect 28142 42406 28172 42458
rect 28196 42406 28206 42458
rect 28206 42406 28252 42458
rect 27956 42404 28012 42406
rect 28036 42404 28092 42406
rect 28116 42404 28172 42406
rect 28196 42404 28252 42406
rect 27956 41370 28012 41372
rect 28036 41370 28092 41372
rect 28116 41370 28172 41372
rect 28196 41370 28252 41372
rect 27956 41318 28002 41370
rect 28002 41318 28012 41370
rect 28036 41318 28066 41370
rect 28066 41318 28078 41370
rect 28078 41318 28092 41370
rect 28116 41318 28130 41370
rect 28130 41318 28142 41370
rect 28142 41318 28172 41370
rect 28196 41318 28206 41370
rect 28206 41318 28252 41370
rect 27956 41316 28012 41318
rect 28036 41316 28092 41318
rect 28116 41316 28172 41318
rect 28196 41316 28252 41318
rect 27956 40282 28012 40284
rect 28036 40282 28092 40284
rect 28116 40282 28172 40284
rect 28196 40282 28252 40284
rect 27956 40230 28002 40282
rect 28002 40230 28012 40282
rect 28036 40230 28066 40282
rect 28066 40230 28078 40282
rect 28078 40230 28092 40282
rect 28116 40230 28130 40282
rect 28130 40230 28142 40282
rect 28142 40230 28172 40282
rect 28196 40230 28206 40282
rect 28206 40230 28252 40282
rect 27956 40228 28012 40230
rect 28036 40228 28092 40230
rect 28116 40228 28172 40230
rect 28196 40228 28252 40230
rect 27956 39194 28012 39196
rect 28036 39194 28092 39196
rect 28116 39194 28172 39196
rect 28196 39194 28252 39196
rect 27956 39142 28002 39194
rect 28002 39142 28012 39194
rect 28036 39142 28066 39194
rect 28066 39142 28078 39194
rect 28078 39142 28092 39194
rect 28116 39142 28130 39194
rect 28130 39142 28142 39194
rect 28142 39142 28172 39194
rect 28196 39142 28206 39194
rect 28206 39142 28252 39194
rect 27956 39140 28012 39142
rect 28036 39140 28092 39142
rect 28116 39140 28172 39142
rect 28196 39140 28252 39142
rect 27956 38106 28012 38108
rect 28036 38106 28092 38108
rect 28116 38106 28172 38108
rect 28196 38106 28252 38108
rect 27956 38054 28002 38106
rect 28002 38054 28012 38106
rect 28036 38054 28066 38106
rect 28066 38054 28078 38106
rect 28078 38054 28092 38106
rect 28116 38054 28130 38106
rect 28130 38054 28142 38106
rect 28142 38054 28172 38106
rect 28196 38054 28206 38106
rect 28206 38054 28252 38106
rect 27956 38052 28012 38054
rect 28036 38052 28092 38054
rect 28116 38052 28172 38054
rect 28196 38052 28252 38054
rect 27956 37018 28012 37020
rect 28036 37018 28092 37020
rect 28116 37018 28172 37020
rect 28196 37018 28252 37020
rect 27956 36966 28002 37018
rect 28002 36966 28012 37018
rect 28036 36966 28066 37018
rect 28066 36966 28078 37018
rect 28078 36966 28092 37018
rect 28116 36966 28130 37018
rect 28130 36966 28142 37018
rect 28142 36966 28172 37018
rect 28196 36966 28206 37018
rect 28206 36966 28252 37018
rect 27956 36964 28012 36966
rect 28036 36964 28092 36966
rect 28116 36964 28172 36966
rect 28196 36964 28252 36966
rect 27956 35930 28012 35932
rect 28036 35930 28092 35932
rect 28116 35930 28172 35932
rect 28196 35930 28252 35932
rect 27956 35878 28002 35930
rect 28002 35878 28012 35930
rect 28036 35878 28066 35930
rect 28066 35878 28078 35930
rect 28078 35878 28092 35930
rect 28116 35878 28130 35930
rect 28130 35878 28142 35930
rect 28142 35878 28172 35930
rect 28196 35878 28206 35930
rect 28206 35878 28252 35930
rect 27956 35876 28012 35878
rect 28036 35876 28092 35878
rect 28116 35876 28172 35878
rect 28196 35876 28252 35878
rect 27956 34842 28012 34844
rect 28036 34842 28092 34844
rect 28116 34842 28172 34844
rect 28196 34842 28252 34844
rect 27956 34790 28002 34842
rect 28002 34790 28012 34842
rect 28036 34790 28066 34842
rect 28066 34790 28078 34842
rect 28078 34790 28092 34842
rect 28116 34790 28130 34842
rect 28130 34790 28142 34842
rect 28142 34790 28172 34842
rect 28196 34790 28206 34842
rect 28206 34790 28252 34842
rect 27956 34788 28012 34790
rect 28036 34788 28092 34790
rect 28116 34788 28172 34790
rect 28196 34788 28252 34790
rect 27956 33754 28012 33756
rect 28036 33754 28092 33756
rect 28116 33754 28172 33756
rect 28196 33754 28252 33756
rect 27956 33702 28002 33754
rect 28002 33702 28012 33754
rect 28036 33702 28066 33754
rect 28066 33702 28078 33754
rect 28078 33702 28092 33754
rect 28116 33702 28130 33754
rect 28130 33702 28142 33754
rect 28142 33702 28172 33754
rect 28196 33702 28206 33754
rect 28206 33702 28252 33754
rect 27956 33700 28012 33702
rect 28036 33700 28092 33702
rect 28116 33700 28172 33702
rect 28196 33700 28252 33702
rect 27526 33632 27582 33688
rect 37956 54426 38012 54428
rect 38036 54426 38092 54428
rect 38116 54426 38172 54428
rect 38196 54426 38252 54428
rect 37956 54374 38002 54426
rect 38002 54374 38012 54426
rect 38036 54374 38066 54426
rect 38066 54374 38078 54426
rect 38078 54374 38092 54426
rect 38116 54374 38130 54426
rect 38130 54374 38142 54426
rect 38142 54374 38172 54426
rect 38196 54374 38206 54426
rect 38206 54374 38252 54426
rect 37956 54372 38012 54374
rect 38036 54372 38092 54374
rect 38116 54372 38172 54374
rect 38196 54372 38252 54374
rect 48226 55392 48282 55448
rect 47956 54426 48012 54428
rect 48036 54426 48092 54428
rect 48116 54426 48172 54428
rect 48196 54426 48252 54428
rect 47956 54374 48002 54426
rect 48002 54374 48012 54426
rect 48036 54374 48066 54426
rect 48066 54374 48078 54426
rect 48078 54374 48092 54426
rect 48116 54374 48130 54426
rect 48130 54374 48142 54426
rect 48142 54374 48172 54426
rect 48196 54374 48206 54426
rect 48206 54374 48252 54426
rect 47956 54372 48012 54374
rect 48036 54372 48092 54374
rect 48116 54372 48172 54374
rect 48196 54372 48252 54374
rect 32956 53882 33012 53884
rect 33036 53882 33092 53884
rect 33116 53882 33172 53884
rect 33196 53882 33252 53884
rect 32956 53830 33002 53882
rect 33002 53830 33012 53882
rect 33036 53830 33066 53882
rect 33066 53830 33078 53882
rect 33078 53830 33092 53882
rect 33116 53830 33130 53882
rect 33130 53830 33142 53882
rect 33142 53830 33172 53882
rect 33196 53830 33206 53882
rect 33206 53830 33252 53882
rect 32956 53828 33012 53830
rect 33036 53828 33092 53830
rect 33116 53828 33172 53830
rect 33196 53828 33252 53830
rect 37956 53338 38012 53340
rect 38036 53338 38092 53340
rect 38116 53338 38172 53340
rect 38196 53338 38252 53340
rect 37956 53286 38002 53338
rect 38002 53286 38012 53338
rect 38036 53286 38066 53338
rect 38066 53286 38078 53338
rect 38078 53286 38092 53338
rect 38116 53286 38130 53338
rect 38130 53286 38142 53338
rect 38142 53286 38172 53338
rect 38196 53286 38206 53338
rect 38206 53286 38252 53338
rect 37956 53284 38012 53286
rect 38036 53284 38092 53286
rect 38116 53284 38172 53286
rect 38196 53284 38252 53286
rect 32956 52794 33012 52796
rect 33036 52794 33092 52796
rect 33116 52794 33172 52796
rect 33196 52794 33252 52796
rect 32956 52742 33002 52794
rect 33002 52742 33012 52794
rect 33036 52742 33066 52794
rect 33066 52742 33078 52794
rect 33078 52742 33092 52794
rect 33116 52742 33130 52794
rect 33130 52742 33142 52794
rect 33142 52742 33172 52794
rect 33196 52742 33206 52794
rect 33206 52742 33252 52794
rect 32956 52740 33012 52742
rect 33036 52740 33092 52742
rect 33116 52740 33172 52742
rect 33196 52740 33252 52742
rect 32956 51706 33012 51708
rect 33036 51706 33092 51708
rect 33116 51706 33172 51708
rect 33196 51706 33252 51708
rect 32956 51654 33002 51706
rect 33002 51654 33012 51706
rect 33036 51654 33066 51706
rect 33066 51654 33078 51706
rect 33078 51654 33092 51706
rect 33116 51654 33130 51706
rect 33130 51654 33142 51706
rect 33142 51654 33172 51706
rect 33196 51654 33206 51706
rect 33206 51654 33252 51706
rect 32956 51652 33012 51654
rect 33036 51652 33092 51654
rect 33116 51652 33172 51654
rect 33196 51652 33252 51654
rect 32956 50618 33012 50620
rect 33036 50618 33092 50620
rect 33116 50618 33172 50620
rect 33196 50618 33252 50620
rect 32956 50566 33002 50618
rect 33002 50566 33012 50618
rect 33036 50566 33066 50618
rect 33066 50566 33078 50618
rect 33078 50566 33092 50618
rect 33116 50566 33130 50618
rect 33130 50566 33142 50618
rect 33142 50566 33172 50618
rect 33196 50566 33206 50618
rect 33206 50566 33252 50618
rect 32956 50564 33012 50566
rect 33036 50564 33092 50566
rect 33116 50564 33172 50566
rect 33196 50564 33252 50566
rect 32956 49530 33012 49532
rect 33036 49530 33092 49532
rect 33116 49530 33172 49532
rect 33196 49530 33252 49532
rect 32956 49478 33002 49530
rect 33002 49478 33012 49530
rect 33036 49478 33066 49530
rect 33066 49478 33078 49530
rect 33078 49478 33092 49530
rect 33116 49478 33130 49530
rect 33130 49478 33142 49530
rect 33142 49478 33172 49530
rect 33196 49478 33206 49530
rect 33206 49478 33252 49530
rect 32956 49476 33012 49478
rect 33036 49476 33092 49478
rect 33116 49476 33172 49478
rect 33196 49476 33252 49478
rect 32956 48442 33012 48444
rect 33036 48442 33092 48444
rect 33116 48442 33172 48444
rect 33196 48442 33252 48444
rect 32956 48390 33002 48442
rect 33002 48390 33012 48442
rect 33036 48390 33066 48442
rect 33066 48390 33078 48442
rect 33078 48390 33092 48442
rect 33116 48390 33130 48442
rect 33130 48390 33142 48442
rect 33142 48390 33172 48442
rect 33196 48390 33206 48442
rect 33206 48390 33252 48442
rect 32956 48388 33012 48390
rect 33036 48388 33092 48390
rect 33116 48388 33172 48390
rect 33196 48388 33252 48390
rect 32956 47354 33012 47356
rect 33036 47354 33092 47356
rect 33116 47354 33172 47356
rect 33196 47354 33252 47356
rect 32956 47302 33002 47354
rect 33002 47302 33012 47354
rect 33036 47302 33066 47354
rect 33066 47302 33078 47354
rect 33078 47302 33092 47354
rect 33116 47302 33130 47354
rect 33130 47302 33142 47354
rect 33142 47302 33172 47354
rect 33196 47302 33206 47354
rect 33206 47302 33252 47354
rect 32956 47300 33012 47302
rect 33036 47300 33092 47302
rect 33116 47300 33172 47302
rect 33196 47300 33252 47302
rect 32956 46266 33012 46268
rect 33036 46266 33092 46268
rect 33116 46266 33172 46268
rect 33196 46266 33252 46268
rect 32956 46214 33002 46266
rect 33002 46214 33012 46266
rect 33036 46214 33066 46266
rect 33066 46214 33078 46266
rect 33078 46214 33092 46266
rect 33116 46214 33130 46266
rect 33130 46214 33142 46266
rect 33142 46214 33172 46266
rect 33196 46214 33206 46266
rect 33206 46214 33252 46266
rect 32956 46212 33012 46214
rect 33036 46212 33092 46214
rect 33116 46212 33172 46214
rect 33196 46212 33252 46214
rect 32956 45178 33012 45180
rect 33036 45178 33092 45180
rect 33116 45178 33172 45180
rect 33196 45178 33252 45180
rect 32956 45126 33002 45178
rect 33002 45126 33012 45178
rect 33036 45126 33066 45178
rect 33066 45126 33078 45178
rect 33078 45126 33092 45178
rect 33116 45126 33130 45178
rect 33130 45126 33142 45178
rect 33142 45126 33172 45178
rect 33196 45126 33206 45178
rect 33206 45126 33252 45178
rect 32956 45124 33012 45126
rect 33036 45124 33092 45126
rect 33116 45124 33172 45126
rect 33196 45124 33252 45126
rect 32956 44090 33012 44092
rect 33036 44090 33092 44092
rect 33116 44090 33172 44092
rect 33196 44090 33252 44092
rect 32956 44038 33002 44090
rect 33002 44038 33012 44090
rect 33036 44038 33066 44090
rect 33066 44038 33078 44090
rect 33078 44038 33092 44090
rect 33116 44038 33130 44090
rect 33130 44038 33142 44090
rect 33142 44038 33172 44090
rect 33196 44038 33206 44090
rect 33206 44038 33252 44090
rect 32956 44036 33012 44038
rect 33036 44036 33092 44038
rect 33116 44036 33172 44038
rect 33196 44036 33252 44038
rect 32956 43002 33012 43004
rect 33036 43002 33092 43004
rect 33116 43002 33172 43004
rect 33196 43002 33252 43004
rect 32956 42950 33002 43002
rect 33002 42950 33012 43002
rect 33036 42950 33066 43002
rect 33066 42950 33078 43002
rect 33078 42950 33092 43002
rect 33116 42950 33130 43002
rect 33130 42950 33142 43002
rect 33142 42950 33172 43002
rect 33196 42950 33206 43002
rect 33206 42950 33252 43002
rect 32956 42948 33012 42950
rect 33036 42948 33092 42950
rect 33116 42948 33172 42950
rect 33196 42948 33252 42950
rect 32956 41914 33012 41916
rect 33036 41914 33092 41916
rect 33116 41914 33172 41916
rect 33196 41914 33252 41916
rect 32956 41862 33002 41914
rect 33002 41862 33012 41914
rect 33036 41862 33066 41914
rect 33066 41862 33078 41914
rect 33078 41862 33092 41914
rect 33116 41862 33130 41914
rect 33130 41862 33142 41914
rect 33142 41862 33172 41914
rect 33196 41862 33206 41914
rect 33206 41862 33252 41914
rect 32956 41860 33012 41862
rect 33036 41860 33092 41862
rect 33116 41860 33172 41862
rect 33196 41860 33252 41862
rect 32956 40826 33012 40828
rect 33036 40826 33092 40828
rect 33116 40826 33172 40828
rect 33196 40826 33252 40828
rect 32956 40774 33002 40826
rect 33002 40774 33012 40826
rect 33036 40774 33066 40826
rect 33066 40774 33078 40826
rect 33078 40774 33092 40826
rect 33116 40774 33130 40826
rect 33130 40774 33142 40826
rect 33142 40774 33172 40826
rect 33196 40774 33206 40826
rect 33206 40774 33252 40826
rect 32956 40772 33012 40774
rect 33036 40772 33092 40774
rect 33116 40772 33172 40774
rect 33196 40772 33252 40774
rect 32956 39738 33012 39740
rect 33036 39738 33092 39740
rect 33116 39738 33172 39740
rect 33196 39738 33252 39740
rect 32956 39686 33002 39738
rect 33002 39686 33012 39738
rect 33036 39686 33066 39738
rect 33066 39686 33078 39738
rect 33078 39686 33092 39738
rect 33116 39686 33130 39738
rect 33130 39686 33142 39738
rect 33142 39686 33172 39738
rect 33196 39686 33206 39738
rect 33206 39686 33252 39738
rect 32956 39684 33012 39686
rect 33036 39684 33092 39686
rect 33116 39684 33172 39686
rect 33196 39684 33252 39686
rect 32956 38650 33012 38652
rect 33036 38650 33092 38652
rect 33116 38650 33172 38652
rect 33196 38650 33252 38652
rect 32956 38598 33002 38650
rect 33002 38598 33012 38650
rect 33036 38598 33066 38650
rect 33066 38598 33078 38650
rect 33078 38598 33092 38650
rect 33116 38598 33130 38650
rect 33130 38598 33142 38650
rect 33142 38598 33172 38650
rect 33196 38598 33206 38650
rect 33206 38598 33252 38650
rect 32956 38596 33012 38598
rect 33036 38596 33092 38598
rect 33116 38596 33172 38598
rect 33196 38596 33252 38598
rect 32956 37562 33012 37564
rect 33036 37562 33092 37564
rect 33116 37562 33172 37564
rect 33196 37562 33252 37564
rect 32956 37510 33002 37562
rect 33002 37510 33012 37562
rect 33036 37510 33066 37562
rect 33066 37510 33078 37562
rect 33078 37510 33092 37562
rect 33116 37510 33130 37562
rect 33130 37510 33142 37562
rect 33142 37510 33172 37562
rect 33196 37510 33206 37562
rect 33206 37510 33252 37562
rect 32956 37508 33012 37510
rect 33036 37508 33092 37510
rect 33116 37508 33172 37510
rect 33196 37508 33252 37510
rect 32956 36474 33012 36476
rect 33036 36474 33092 36476
rect 33116 36474 33172 36476
rect 33196 36474 33252 36476
rect 32956 36422 33002 36474
rect 33002 36422 33012 36474
rect 33036 36422 33066 36474
rect 33066 36422 33078 36474
rect 33078 36422 33092 36474
rect 33116 36422 33130 36474
rect 33130 36422 33142 36474
rect 33142 36422 33172 36474
rect 33196 36422 33206 36474
rect 33206 36422 33252 36474
rect 32956 36420 33012 36422
rect 33036 36420 33092 36422
rect 33116 36420 33172 36422
rect 33196 36420 33252 36422
rect 32956 35386 33012 35388
rect 33036 35386 33092 35388
rect 33116 35386 33172 35388
rect 33196 35386 33252 35388
rect 32956 35334 33002 35386
rect 33002 35334 33012 35386
rect 33036 35334 33066 35386
rect 33066 35334 33078 35386
rect 33078 35334 33092 35386
rect 33116 35334 33130 35386
rect 33130 35334 33142 35386
rect 33142 35334 33172 35386
rect 33196 35334 33206 35386
rect 33206 35334 33252 35386
rect 32956 35332 33012 35334
rect 33036 35332 33092 35334
rect 33116 35332 33172 35334
rect 33196 35332 33252 35334
rect 32956 34298 33012 34300
rect 33036 34298 33092 34300
rect 33116 34298 33172 34300
rect 33196 34298 33252 34300
rect 32956 34246 33002 34298
rect 33002 34246 33012 34298
rect 33036 34246 33066 34298
rect 33066 34246 33078 34298
rect 33078 34246 33092 34298
rect 33116 34246 33130 34298
rect 33130 34246 33142 34298
rect 33142 34246 33172 34298
rect 33196 34246 33206 34298
rect 33206 34246 33252 34298
rect 32956 34244 33012 34246
rect 33036 34244 33092 34246
rect 33116 34244 33172 34246
rect 33196 34244 33252 34246
rect 28906 33224 28962 33280
rect 32956 33210 33012 33212
rect 33036 33210 33092 33212
rect 33116 33210 33172 33212
rect 33196 33210 33252 33212
rect 32956 33158 33002 33210
rect 33002 33158 33012 33210
rect 33036 33158 33066 33210
rect 33066 33158 33078 33210
rect 33078 33158 33092 33210
rect 33116 33158 33130 33210
rect 33130 33158 33142 33210
rect 33142 33158 33172 33210
rect 33196 33158 33206 33210
rect 33206 33158 33252 33210
rect 32956 33156 33012 33158
rect 33036 33156 33092 33158
rect 33116 33156 33172 33158
rect 33196 33156 33252 33158
rect 27956 32666 28012 32668
rect 28036 32666 28092 32668
rect 28116 32666 28172 32668
rect 28196 32666 28252 32668
rect 27956 32614 28002 32666
rect 28002 32614 28012 32666
rect 28036 32614 28066 32666
rect 28066 32614 28078 32666
rect 28078 32614 28092 32666
rect 28116 32614 28130 32666
rect 28130 32614 28142 32666
rect 28142 32614 28172 32666
rect 28196 32614 28206 32666
rect 28206 32614 28252 32666
rect 27956 32612 28012 32614
rect 28036 32612 28092 32614
rect 28116 32612 28172 32614
rect 28196 32612 28252 32614
rect 32956 32122 33012 32124
rect 33036 32122 33092 32124
rect 33116 32122 33172 32124
rect 33196 32122 33252 32124
rect 32956 32070 33002 32122
rect 33002 32070 33012 32122
rect 33036 32070 33066 32122
rect 33066 32070 33078 32122
rect 33078 32070 33092 32122
rect 33116 32070 33130 32122
rect 33130 32070 33142 32122
rect 33142 32070 33172 32122
rect 33196 32070 33206 32122
rect 33206 32070 33252 32122
rect 32956 32068 33012 32070
rect 33036 32068 33092 32070
rect 33116 32068 33172 32070
rect 33196 32068 33252 32070
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 3422 8744 3478 8800
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3422 1808 3478 1864
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 9862 2372 9918 2408
rect 9862 2352 9864 2372
rect 9864 2352 9916 2372
rect 9916 2352 9918 2372
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 20258 3596 20314 3632
rect 20258 3576 20260 3596
rect 20260 3576 20312 3596
rect 20312 3576 20314 3596
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27956 31578 28012 31580
rect 28036 31578 28092 31580
rect 28116 31578 28172 31580
rect 28196 31578 28252 31580
rect 27956 31526 28002 31578
rect 28002 31526 28012 31578
rect 28036 31526 28066 31578
rect 28066 31526 28078 31578
rect 28078 31526 28092 31578
rect 28116 31526 28130 31578
rect 28130 31526 28142 31578
rect 28142 31526 28172 31578
rect 28196 31526 28206 31578
rect 28206 31526 28252 31578
rect 27956 31524 28012 31526
rect 28036 31524 28092 31526
rect 28116 31524 28172 31526
rect 28196 31524 28252 31526
rect 27956 30490 28012 30492
rect 28036 30490 28092 30492
rect 28116 30490 28172 30492
rect 28196 30490 28252 30492
rect 27956 30438 28002 30490
rect 28002 30438 28012 30490
rect 28036 30438 28066 30490
rect 28066 30438 28078 30490
rect 28078 30438 28092 30490
rect 28116 30438 28130 30490
rect 28130 30438 28142 30490
rect 28142 30438 28172 30490
rect 28196 30438 28206 30490
rect 28206 30438 28252 30490
rect 27956 30436 28012 30438
rect 28036 30436 28092 30438
rect 28116 30436 28172 30438
rect 28196 30436 28252 30438
rect 27956 29402 28012 29404
rect 28036 29402 28092 29404
rect 28116 29402 28172 29404
rect 28196 29402 28252 29404
rect 27956 29350 28002 29402
rect 28002 29350 28012 29402
rect 28036 29350 28066 29402
rect 28066 29350 28078 29402
rect 28078 29350 28092 29402
rect 28116 29350 28130 29402
rect 28130 29350 28142 29402
rect 28142 29350 28172 29402
rect 28196 29350 28206 29402
rect 28206 29350 28252 29402
rect 27956 29348 28012 29350
rect 28036 29348 28092 29350
rect 28116 29348 28172 29350
rect 28196 29348 28252 29350
rect 27956 28314 28012 28316
rect 28036 28314 28092 28316
rect 28116 28314 28172 28316
rect 28196 28314 28252 28316
rect 27956 28262 28002 28314
rect 28002 28262 28012 28314
rect 28036 28262 28066 28314
rect 28066 28262 28078 28314
rect 28078 28262 28092 28314
rect 28116 28262 28130 28314
rect 28130 28262 28142 28314
rect 28142 28262 28172 28314
rect 28196 28262 28206 28314
rect 28206 28262 28252 28314
rect 27956 28260 28012 28262
rect 28036 28260 28092 28262
rect 28116 28260 28172 28262
rect 28196 28260 28252 28262
rect 25318 5072 25374 5128
rect 27956 27226 28012 27228
rect 28036 27226 28092 27228
rect 28116 27226 28172 27228
rect 28196 27226 28252 27228
rect 27956 27174 28002 27226
rect 28002 27174 28012 27226
rect 28036 27174 28066 27226
rect 28066 27174 28078 27226
rect 28078 27174 28092 27226
rect 28116 27174 28130 27226
rect 28130 27174 28142 27226
rect 28142 27174 28172 27226
rect 28196 27174 28206 27226
rect 28206 27174 28252 27226
rect 27956 27172 28012 27174
rect 28036 27172 28092 27174
rect 28116 27172 28172 27174
rect 28196 27172 28252 27174
rect 27956 26138 28012 26140
rect 28036 26138 28092 26140
rect 28116 26138 28172 26140
rect 28196 26138 28252 26140
rect 27956 26086 28002 26138
rect 28002 26086 28012 26138
rect 28036 26086 28066 26138
rect 28066 26086 28078 26138
rect 28078 26086 28092 26138
rect 28116 26086 28130 26138
rect 28130 26086 28142 26138
rect 28142 26086 28172 26138
rect 28196 26086 28206 26138
rect 28206 26086 28252 26138
rect 27956 26084 28012 26086
rect 28036 26084 28092 26086
rect 28116 26084 28172 26086
rect 28196 26084 28252 26086
rect 27956 25050 28012 25052
rect 28036 25050 28092 25052
rect 28116 25050 28172 25052
rect 28196 25050 28252 25052
rect 27956 24998 28002 25050
rect 28002 24998 28012 25050
rect 28036 24998 28066 25050
rect 28066 24998 28078 25050
rect 28078 24998 28092 25050
rect 28116 24998 28130 25050
rect 28130 24998 28142 25050
rect 28142 24998 28172 25050
rect 28196 24998 28206 25050
rect 28206 24998 28252 25050
rect 27956 24996 28012 24998
rect 28036 24996 28092 24998
rect 28116 24996 28172 24998
rect 28196 24996 28252 24998
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 26974 14356 26976 14376
rect 26976 14356 27028 14376
rect 27028 14356 27030 14376
rect 26974 14320 27030 14356
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 28262 14764 28264 14784
rect 28264 14764 28316 14784
rect 28316 14764 28318 14784
rect 28262 14728 28318 14764
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27618 12416 27674 12472
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27802 12416 27858 12472
rect 28170 12316 28172 12336
rect 28172 12316 28224 12336
rect 28224 12316 28226 12336
rect 28170 12280 28226 12316
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 28354 11736 28410 11792
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 28630 10648 28686 10704
rect 32956 31034 33012 31036
rect 33036 31034 33092 31036
rect 33116 31034 33172 31036
rect 33196 31034 33252 31036
rect 32956 30982 33002 31034
rect 33002 30982 33012 31034
rect 33036 30982 33066 31034
rect 33066 30982 33078 31034
rect 33078 30982 33092 31034
rect 33116 30982 33130 31034
rect 33130 30982 33142 31034
rect 33142 30982 33172 31034
rect 33196 30982 33206 31034
rect 33206 30982 33252 31034
rect 32956 30980 33012 30982
rect 33036 30980 33092 30982
rect 33116 30980 33172 30982
rect 33196 30980 33252 30982
rect 32956 29946 33012 29948
rect 33036 29946 33092 29948
rect 33116 29946 33172 29948
rect 33196 29946 33252 29948
rect 32956 29894 33002 29946
rect 33002 29894 33012 29946
rect 33036 29894 33066 29946
rect 33066 29894 33078 29946
rect 33078 29894 33092 29946
rect 33116 29894 33130 29946
rect 33130 29894 33142 29946
rect 33142 29894 33172 29946
rect 33196 29894 33206 29946
rect 33206 29894 33252 29946
rect 32956 29892 33012 29894
rect 33036 29892 33092 29894
rect 33116 29892 33172 29894
rect 33196 29892 33252 29894
rect 32956 28858 33012 28860
rect 33036 28858 33092 28860
rect 33116 28858 33172 28860
rect 33196 28858 33252 28860
rect 32956 28806 33002 28858
rect 33002 28806 33012 28858
rect 33036 28806 33066 28858
rect 33066 28806 33078 28858
rect 33078 28806 33092 28858
rect 33116 28806 33130 28858
rect 33130 28806 33142 28858
rect 33142 28806 33172 28858
rect 33196 28806 33206 28858
rect 33206 28806 33252 28858
rect 32956 28804 33012 28806
rect 33036 28804 33092 28806
rect 33116 28804 33172 28806
rect 33196 28804 33252 28806
rect 29090 12860 29092 12880
rect 29092 12860 29144 12880
rect 29144 12860 29146 12880
rect 29090 12824 29146 12860
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 29642 10920 29698 10976
rect 30930 17196 30986 17232
rect 30930 17176 30932 17196
rect 30932 17176 30984 17196
rect 30984 17176 30986 17196
rect 29918 11192 29974 11248
rect 30470 12824 30526 12880
rect 30286 9424 30342 9480
rect 30562 11192 30618 11248
rect 30746 10648 30802 10704
rect 31850 24928 31906 24984
rect 32034 17584 32090 17640
rect 31390 11192 31446 11248
rect 31666 12280 31722 12336
rect 32586 24692 32588 24712
rect 32588 24692 32640 24712
rect 32640 24692 32642 24712
rect 32586 24656 32642 24692
rect 32956 27770 33012 27772
rect 33036 27770 33092 27772
rect 33116 27770 33172 27772
rect 33196 27770 33252 27772
rect 32956 27718 33002 27770
rect 33002 27718 33012 27770
rect 33036 27718 33066 27770
rect 33066 27718 33078 27770
rect 33078 27718 33092 27770
rect 33116 27718 33130 27770
rect 33130 27718 33142 27770
rect 33142 27718 33172 27770
rect 33196 27718 33206 27770
rect 33206 27718 33252 27770
rect 32956 27716 33012 27718
rect 33036 27716 33092 27718
rect 33116 27716 33172 27718
rect 33196 27716 33252 27718
rect 32956 26682 33012 26684
rect 33036 26682 33092 26684
rect 33116 26682 33172 26684
rect 33196 26682 33252 26684
rect 32956 26630 33002 26682
rect 33002 26630 33012 26682
rect 33036 26630 33066 26682
rect 33066 26630 33078 26682
rect 33078 26630 33092 26682
rect 33116 26630 33130 26682
rect 33130 26630 33142 26682
rect 33142 26630 33172 26682
rect 33196 26630 33206 26682
rect 33206 26630 33252 26682
rect 32956 26628 33012 26630
rect 33036 26628 33092 26630
rect 33116 26628 33172 26630
rect 33196 26628 33252 26630
rect 33046 25744 33102 25800
rect 32956 25594 33012 25596
rect 33036 25594 33092 25596
rect 33116 25594 33172 25596
rect 33196 25594 33252 25596
rect 32956 25542 33002 25594
rect 33002 25542 33012 25594
rect 33036 25542 33066 25594
rect 33066 25542 33078 25594
rect 33078 25542 33092 25594
rect 33116 25542 33130 25594
rect 33130 25542 33142 25594
rect 33142 25542 33172 25594
rect 33196 25542 33206 25594
rect 33206 25542 33252 25594
rect 32956 25540 33012 25542
rect 33036 25540 33092 25542
rect 33116 25540 33172 25542
rect 33196 25540 33252 25542
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32126 9036 32182 9072
rect 32126 9016 32128 9036
rect 32128 9016 32180 9036
rect 32180 9016 32182 9036
rect 32586 11076 32642 11112
rect 32586 11056 32588 11076
rect 32588 11056 32640 11076
rect 32640 11056 32642 11076
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 37956 52250 38012 52252
rect 38036 52250 38092 52252
rect 38116 52250 38172 52252
rect 38196 52250 38252 52252
rect 37956 52198 38002 52250
rect 38002 52198 38012 52250
rect 38036 52198 38066 52250
rect 38066 52198 38078 52250
rect 38078 52198 38092 52250
rect 38116 52198 38130 52250
rect 38130 52198 38142 52250
rect 38142 52198 38172 52250
rect 38196 52198 38206 52250
rect 38206 52198 38252 52250
rect 37956 52196 38012 52198
rect 38036 52196 38092 52198
rect 38116 52196 38172 52198
rect 38196 52196 38252 52198
rect 37956 51162 38012 51164
rect 38036 51162 38092 51164
rect 38116 51162 38172 51164
rect 38196 51162 38252 51164
rect 37956 51110 38002 51162
rect 38002 51110 38012 51162
rect 38036 51110 38066 51162
rect 38066 51110 38078 51162
rect 38078 51110 38092 51162
rect 38116 51110 38130 51162
rect 38130 51110 38142 51162
rect 38142 51110 38172 51162
rect 38196 51110 38206 51162
rect 38206 51110 38252 51162
rect 37956 51108 38012 51110
rect 38036 51108 38092 51110
rect 38116 51108 38172 51110
rect 38196 51108 38252 51110
rect 34518 29008 34574 29064
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 33966 17176 34022 17232
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 33230 9560 33286 9616
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32586 8880 32642 8936
rect 33506 9016 33562 9072
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 37956 50074 38012 50076
rect 38036 50074 38092 50076
rect 38116 50074 38172 50076
rect 38196 50074 38252 50076
rect 37956 50022 38002 50074
rect 38002 50022 38012 50074
rect 38036 50022 38066 50074
rect 38066 50022 38078 50074
rect 38078 50022 38092 50074
rect 38116 50022 38130 50074
rect 38130 50022 38142 50074
rect 38142 50022 38172 50074
rect 38196 50022 38206 50074
rect 38206 50022 38252 50074
rect 37956 50020 38012 50022
rect 38036 50020 38092 50022
rect 38116 50020 38172 50022
rect 38196 50020 38252 50022
rect 37956 48986 38012 48988
rect 38036 48986 38092 48988
rect 38116 48986 38172 48988
rect 38196 48986 38252 48988
rect 37956 48934 38002 48986
rect 38002 48934 38012 48986
rect 38036 48934 38066 48986
rect 38066 48934 38078 48986
rect 38078 48934 38092 48986
rect 38116 48934 38130 48986
rect 38130 48934 38142 48986
rect 38142 48934 38172 48986
rect 38196 48934 38206 48986
rect 38206 48934 38252 48986
rect 37956 48932 38012 48934
rect 38036 48932 38092 48934
rect 38116 48932 38172 48934
rect 38196 48932 38252 48934
rect 37956 47898 38012 47900
rect 38036 47898 38092 47900
rect 38116 47898 38172 47900
rect 38196 47898 38252 47900
rect 37956 47846 38002 47898
rect 38002 47846 38012 47898
rect 38036 47846 38066 47898
rect 38066 47846 38078 47898
rect 38078 47846 38092 47898
rect 38116 47846 38130 47898
rect 38130 47846 38142 47898
rect 38142 47846 38172 47898
rect 38196 47846 38206 47898
rect 38206 47846 38252 47898
rect 37956 47844 38012 47846
rect 38036 47844 38092 47846
rect 38116 47844 38172 47846
rect 38196 47844 38252 47846
rect 37956 46810 38012 46812
rect 38036 46810 38092 46812
rect 38116 46810 38172 46812
rect 38196 46810 38252 46812
rect 37956 46758 38002 46810
rect 38002 46758 38012 46810
rect 38036 46758 38066 46810
rect 38066 46758 38078 46810
rect 38078 46758 38092 46810
rect 38116 46758 38130 46810
rect 38130 46758 38142 46810
rect 38142 46758 38172 46810
rect 38196 46758 38206 46810
rect 38206 46758 38252 46810
rect 37956 46756 38012 46758
rect 38036 46756 38092 46758
rect 38116 46756 38172 46758
rect 38196 46756 38252 46758
rect 37956 45722 38012 45724
rect 38036 45722 38092 45724
rect 38116 45722 38172 45724
rect 38196 45722 38252 45724
rect 37956 45670 38002 45722
rect 38002 45670 38012 45722
rect 38036 45670 38066 45722
rect 38066 45670 38078 45722
rect 38078 45670 38092 45722
rect 38116 45670 38130 45722
rect 38130 45670 38142 45722
rect 38142 45670 38172 45722
rect 38196 45670 38206 45722
rect 38206 45670 38252 45722
rect 37956 45668 38012 45670
rect 38036 45668 38092 45670
rect 38116 45668 38172 45670
rect 38196 45668 38252 45670
rect 37956 44634 38012 44636
rect 38036 44634 38092 44636
rect 38116 44634 38172 44636
rect 38196 44634 38252 44636
rect 37956 44582 38002 44634
rect 38002 44582 38012 44634
rect 38036 44582 38066 44634
rect 38066 44582 38078 44634
rect 38078 44582 38092 44634
rect 38116 44582 38130 44634
rect 38130 44582 38142 44634
rect 38142 44582 38172 44634
rect 38196 44582 38206 44634
rect 38206 44582 38252 44634
rect 37956 44580 38012 44582
rect 38036 44580 38092 44582
rect 38116 44580 38172 44582
rect 38196 44580 38252 44582
rect 37956 43546 38012 43548
rect 38036 43546 38092 43548
rect 38116 43546 38172 43548
rect 38196 43546 38252 43548
rect 37956 43494 38002 43546
rect 38002 43494 38012 43546
rect 38036 43494 38066 43546
rect 38066 43494 38078 43546
rect 38078 43494 38092 43546
rect 38116 43494 38130 43546
rect 38130 43494 38142 43546
rect 38142 43494 38172 43546
rect 38196 43494 38206 43546
rect 38206 43494 38252 43546
rect 37956 43492 38012 43494
rect 38036 43492 38092 43494
rect 38116 43492 38172 43494
rect 38196 43492 38252 43494
rect 37956 42458 38012 42460
rect 38036 42458 38092 42460
rect 38116 42458 38172 42460
rect 38196 42458 38252 42460
rect 37956 42406 38002 42458
rect 38002 42406 38012 42458
rect 38036 42406 38066 42458
rect 38066 42406 38078 42458
rect 38078 42406 38092 42458
rect 38116 42406 38130 42458
rect 38130 42406 38142 42458
rect 38142 42406 38172 42458
rect 38196 42406 38206 42458
rect 38206 42406 38252 42458
rect 37956 42404 38012 42406
rect 38036 42404 38092 42406
rect 38116 42404 38172 42406
rect 38196 42404 38252 42406
rect 35714 29008 35770 29064
rect 34242 10920 34298 10976
rect 35254 26324 35256 26344
rect 35256 26324 35308 26344
rect 35308 26324 35310 26344
rect 35254 26288 35310 26324
rect 34426 8472 34482 8528
rect 34794 9288 34850 9344
rect 35990 29552 36046 29608
rect 35990 27276 35992 27296
rect 35992 27276 36044 27296
rect 36044 27276 36046 27296
rect 35990 27240 36046 27276
rect 35622 24656 35678 24712
rect 35346 11076 35402 11112
rect 35346 11056 35348 11076
rect 35348 11056 35400 11076
rect 35400 11056 35402 11076
rect 35254 9560 35310 9616
rect 36266 11756 36322 11792
rect 36266 11736 36268 11756
rect 36268 11736 36320 11756
rect 36320 11736 36322 11756
rect 36082 10684 36084 10704
rect 36084 10684 36136 10704
rect 36136 10684 36138 10704
rect 36082 10648 36138 10684
rect 37956 41370 38012 41372
rect 38036 41370 38092 41372
rect 38116 41370 38172 41372
rect 38196 41370 38252 41372
rect 37956 41318 38002 41370
rect 38002 41318 38012 41370
rect 38036 41318 38066 41370
rect 38066 41318 38078 41370
rect 38078 41318 38092 41370
rect 38116 41318 38130 41370
rect 38130 41318 38142 41370
rect 38142 41318 38172 41370
rect 38196 41318 38206 41370
rect 38206 41318 38252 41370
rect 37956 41316 38012 41318
rect 38036 41316 38092 41318
rect 38116 41316 38172 41318
rect 38196 41316 38252 41318
rect 37956 40282 38012 40284
rect 38036 40282 38092 40284
rect 38116 40282 38172 40284
rect 38196 40282 38252 40284
rect 37956 40230 38002 40282
rect 38002 40230 38012 40282
rect 38036 40230 38066 40282
rect 38066 40230 38078 40282
rect 38078 40230 38092 40282
rect 38116 40230 38130 40282
rect 38130 40230 38142 40282
rect 38142 40230 38172 40282
rect 38196 40230 38206 40282
rect 38206 40230 38252 40282
rect 37956 40228 38012 40230
rect 38036 40228 38092 40230
rect 38116 40228 38172 40230
rect 38196 40228 38252 40230
rect 37956 39194 38012 39196
rect 38036 39194 38092 39196
rect 38116 39194 38172 39196
rect 38196 39194 38252 39196
rect 37956 39142 38002 39194
rect 38002 39142 38012 39194
rect 38036 39142 38066 39194
rect 38066 39142 38078 39194
rect 38078 39142 38092 39194
rect 38116 39142 38130 39194
rect 38130 39142 38142 39194
rect 38142 39142 38172 39194
rect 38196 39142 38206 39194
rect 38206 39142 38252 39194
rect 37956 39140 38012 39142
rect 38036 39140 38092 39142
rect 38116 39140 38172 39142
rect 38196 39140 38252 39142
rect 37956 38106 38012 38108
rect 38036 38106 38092 38108
rect 38116 38106 38172 38108
rect 38196 38106 38252 38108
rect 37956 38054 38002 38106
rect 38002 38054 38012 38106
rect 38036 38054 38066 38106
rect 38066 38054 38078 38106
rect 38078 38054 38092 38106
rect 38116 38054 38130 38106
rect 38130 38054 38142 38106
rect 38142 38054 38172 38106
rect 38196 38054 38206 38106
rect 38206 38054 38252 38106
rect 37956 38052 38012 38054
rect 38036 38052 38092 38054
rect 38116 38052 38172 38054
rect 38196 38052 38252 38054
rect 37956 37018 38012 37020
rect 38036 37018 38092 37020
rect 38116 37018 38172 37020
rect 38196 37018 38252 37020
rect 37956 36966 38002 37018
rect 38002 36966 38012 37018
rect 38036 36966 38066 37018
rect 38066 36966 38078 37018
rect 38078 36966 38092 37018
rect 38116 36966 38130 37018
rect 38130 36966 38142 37018
rect 38142 36966 38172 37018
rect 38196 36966 38206 37018
rect 38206 36966 38252 37018
rect 37956 36964 38012 36966
rect 38036 36964 38092 36966
rect 38116 36964 38172 36966
rect 38196 36964 38252 36966
rect 37956 35930 38012 35932
rect 38036 35930 38092 35932
rect 38116 35930 38172 35932
rect 38196 35930 38252 35932
rect 37956 35878 38002 35930
rect 38002 35878 38012 35930
rect 38036 35878 38066 35930
rect 38066 35878 38078 35930
rect 38078 35878 38092 35930
rect 38116 35878 38130 35930
rect 38130 35878 38142 35930
rect 38142 35878 38172 35930
rect 38196 35878 38206 35930
rect 38206 35878 38252 35930
rect 37956 35876 38012 35878
rect 38036 35876 38092 35878
rect 38116 35876 38172 35878
rect 38196 35876 38252 35878
rect 37956 34842 38012 34844
rect 38036 34842 38092 34844
rect 38116 34842 38172 34844
rect 38196 34842 38252 34844
rect 37956 34790 38002 34842
rect 38002 34790 38012 34842
rect 38036 34790 38066 34842
rect 38066 34790 38078 34842
rect 38078 34790 38092 34842
rect 38116 34790 38130 34842
rect 38130 34790 38142 34842
rect 38142 34790 38172 34842
rect 38196 34790 38206 34842
rect 38206 34790 38252 34842
rect 37956 34788 38012 34790
rect 38036 34788 38092 34790
rect 38116 34788 38172 34790
rect 38196 34788 38252 34790
rect 37956 33754 38012 33756
rect 38036 33754 38092 33756
rect 38116 33754 38172 33756
rect 38196 33754 38252 33756
rect 37956 33702 38002 33754
rect 38002 33702 38012 33754
rect 38036 33702 38066 33754
rect 38066 33702 38078 33754
rect 38078 33702 38092 33754
rect 38116 33702 38130 33754
rect 38130 33702 38142 33754
rect 38142 33702 38172 33754
rect 38196 33702 38206 33754
rect 38206 33702 38252 33754
rect 37956 33700 38012 33702
rect 38036 33700 38092 33702
rect 38116 33700 38172 33702
rect 38196 33700 38252 33702
rect 37956 32666 38012 32668
rect 38036 32666 38092 32668
rect 38116 32666 38172 32668
rect 38196 32666 38252 32668
rect 37956 32614 38002 32666
rect 38002 32614 38012 32666
rect 38036 32614 38066 32666
rect 38066 32614 38078 32666
rect 38078 32614 38092 32666
rect 38116 32614 38130 32666
rect 38130 32614 38142 32666
rect 38142 32614 38172 32666
rect 38196 32614 38206 32666
rect 38206 32614 38252 32666
rect 37956 32612 38012 32614
rect 38036 32612 38092 32614
rect 38116 32612 38172 32614
rect 38196 32612 38252 32614
rect 37956 31578 38012 31580
rect 38036 31578 38092 31580
rect 38116 31578 38172 31580
rect 38196 31578 38252 31580
rect 37956 31526 38002 31578
rect 38002 31526 38012 31578
rect 38036 31526 38066 31578
rect 38066 31526 38078 31578
rect 38078 31526 38092 31578
rect 38116 31526 38130 31578
rect 38130 31526 38142 31578
rect 38142 31526 38172 31578
rect 38196 31526 38206 31578
rect 38206 31526 38252 31578
rect 37956 31524 38012 31526
rect 38036 31524 38092 31526
rect 38116 31524 38172 31526
rect 38196 31524 38252 31526
rect 37956 30490 38012 30492
rect 38036 30490 38092 30492
rect 38116 30490 38172 30492
rect 38196 30490 38252 30492
rect 37956 30438 38002 30490
rect 38002 30438 38012 30490
rect 38036 30438 38066 30490
rect 38066 30438 38078 30490
rect 38078 30438 38092 30490
rect 38116 30438 38130 30490
rect 38130 30438 38142 30490
rect 38142 30438 38172 30490
rect 38196 30438 38206 30490
rect 38206 30438 38252 30490
rect 37956 30436 38012 30438
rect 38036 30436 38092 30438
rect 38116 30436 38172 30438
rect 38196 30436 38252 30438
rect 37956 29402 38012 29404
rect 38036 29402 38092 29404
rect 38116 29402 38172 29404
rect 38196 29402 38252 29404
rect 37956 29350 38002 29402
rect 38002 29350 38012 29402
rect 38036 29350 38066 29402
rect 38066 29350 38078 29402
rect 38078 29350 38092 29402
rect 38116 29350 38130 29402
rect 38130 29350 38142 29402
rect 38142 29350 38172 29402
rect 38196 29350 38206 29402
rect 38206 29350 38252 29402
rect 37956 29348 38012 29350
rect 38036 29348 38092 29350
rect 38116 29348 38172 29350
rect 38196 29348 38252 29350
rect 37956 28314 38012 28316
rect 38036 28314 38092 28316
rect 38116 28314 38172 28316
rect 38196 28314 38252 28316
rect 37956 28262 38002 28314
rect 38002 28262 38012 28314
rect 38036 28262 38066 28314
rect 38066 28262 38078 28314
rect 38078 28262 38092 28314
rect 38116 28262 38130 28314
rect 38130 28262 38142 28314
rect 38142 28262 38172 28314
rect 38196 28262 38206 28314
rect 38206 28262 38252 28314
rect 37956 28260 38012 28262
rect 38036 28260 38092 28262
rect 38116 28260 38172 28262
rect 38196 28260 38252 28262
rect 36818 14320 36874 14376
rect 37956 27226 38012 27228
rect 38036 27226 38092 27228
rect 38116 27226 38172 27228
rect 38196 27226 38252 27228
rect 37956 27174 38002 27226
rect 38002 27174 38012 27226
rect 38036 27174 38066 27226
rect 38066 27174 38078 27226
rect 38078 27174 38092 27226
rect 38116 27174 38130 27226
rect 38130 27174 38142 27226
rect 38142 27174 38172 27226
rect 38196 27174 38206 27226
rect 38206 27174 38252 27226
rect 37956 27172 38012 27174
rect 38036 27172 38092 27174
rect 38116 27172 38172 27174
rect 38196 27172 38252 27174
rect 37956 26138 38012 26140
rect 38036 26138 38092 26140
rect 38116 26138 38172 26140
rect 38196 26138 38252 26140
rect 37956 26086 38002 26138
rect 38002 26086 38012 26138
rect 38036 26086 38066 26138
rect 38066 26086 38078 26138
rect 38078 26086 38092 26138
rect 38116 26086 38130 26138
rect 38130 26086 38142 26138
rect 38142 26086 38172 26138
rect 38196 26086 38206 26138
rect 38206 26086 38252 26138
rect 37956 26084 38012 26086
rect 38036 26084 38092 26086
rect 38116 26084 38172 26086
rect 38196 26084 38252 26086
rect 37956 25050 38012 25052
rect 38036 25050 38092 25052
rect 38116 25050 38172 25052
rect 38196 25050 38252 25052
rect 37956 24998 38002 25050
rect 38002 24998 38012 25050
rect 38036 24998 38066 25050
rect 38066 24998 38078 25050
rect 38078 24998 38092 25050
rect 38116 24998 38130 25050
rect 38130 24998 38142 25050
rect 38142 24998 38172 25050
rect 38196 24998 38206 25050
rect 38206 24998 38252 25050
rect 37956 24996 38012 24998
rect 38036 24996 38092 24998
rect 38116 24996 38172 24998
rect 38196 24996 38252 24998
rect 40590 33360 40646 33416
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37830 23568 37886 23624
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 36542 9424 36598 9480
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37370 9288 37426 9344
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 38290 12144 38346 12200
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 38290 11600 38346 11656
rect 38290 11192 38346 11248
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 41234 33360 41290 33416
rect 42956 53882 43012 53884
rect 43036 53882 43092 53884
rect 43116 53882 43172 53884
rect 43196 53882 43252 53884
rect 42956 53830 43002 53882
rect 43002 53830 43012 53882
rect 43036 53830 43066 53882
rect 43066 53830 43078 53882
rect 43078 53830 43092 53882
rect 43116 53830 43130 53882
rect 43130 53830 43142 53882
rect 43142 53830 43172 53882
rect 43196 53830 43206 53882
rect 43206 53830 43252 53882
rect 42956 53828 43012 53830
rect 43036 53828 43092 53830
rect 43116 53828 43172 53830
rect 43196 53828 43252 53830
rect 42956 52794 43012 52796
rect 43036 52794 43092 52796
rect 43116 52794 43172 52796
rect 43196 52794 43252 52796
rect 42956 52742 43002 52794
rect 43002 52742 43012 52794
rect 43036 52742 43066 52794
rect 43066 52742 43078 52794
rect 43078 52742 43092 52794
rect 43116 52742 43130 52794
rect 43130 52742 43142 52794
rect 43142 52742 43172 52794
rect 43196 52742 43206 52794
rect 43206 52742 43252 52794
rect 42956 52740 43012 52742
rect 43036 52740 43092 52742
rect 43116 52740 43172 52742
rect 43196 52740 43252 52742
rect 42956 51706 43012 51708
rect 43036 51706 43092 51708
rect 43116 51706 43172 51708
rect 43196 51706 43252 51708
rect 42956 51654 43002 51706
rect 43002 51654 43012 51706
rect 43036 51654 43066 51706
rect 43066 51654 43078 51706
rect 43078 51654 43092 51706
rect 43116 51654 43130 51706
rect 43130 51654 43142 51706
rect 43142 51654 43172 51706
rect 43196 51654 43206 51706
rect 43206 51654 43252 51706
rect 42956 51652 43012 51654
rect 43036 51652 43092 51654
rect 43116 51652 43172 51654
rect 43196 51652 43252 51654
rect 42956 50618 43012 50620
rect 43036 50618 43092 50620
rect 43116 50618 43172 50620
rect 43196 50618 43252 50620
rect 42956 50566 43002 50618
rect 43002 50566 43012 50618
rect 43036 50566 43066 50618
rect 43066 50566 43078 50618
rect 43078 50566 43092 50618
rect 43116 50566 43130 50618
rect 43130 50566 43142 50618
rect 43142 50566 43172 50618
rect 43196 50566 43206 50618
rect 43206 50566 43252 50618
rect 42956 50564 43012 50566
rect 43036 50564 43092 50566
rect 43116 50564 43172 50566
rect 43196 50564 43252 50566
rect 42956 49530 43012 49532
rect 43036 49530 43092 49532
rect 43116 49530 43172 49532
rect 43196 49530 43252 49532
rect 42956 49478 43002 49530
rect 43002 49478 43012 49530
rect 43036 49478 43066 49530
rect 43066 49478 43078 49530
rect 43078 49478 43092 49530
rect 43116 49478 43130 49530
rect 43130 49478 43142 49530
rect 43142 49478 43172 49530
rect 43196 49478 43206 49530
rect 43206 49478 43252 49530
rect 42956 49476 43012 49478
rect 43036 49476 43092 49478
rect 43116 49476 43172 49478
rect 43196 49476 43252 49478
rect 42956 48442 43012 48444
rect 43036 48442 43092 48444
rect 43116 48442 43172 48444
rect 43196 48442 43252 48444
rect 42956 48390 43002 48442
rect 43002 48390 43012 48442
rect 43036 48390 43066 48442
rect 43066 48390 43078 48442
rect 43078 48390 43092 48442
rect 43116 48390 43130 48442
rect 43130 48390 43142 48442
rect 43142 48390 43172 48442
rect 43196 48390 43206 48442
rect 43206 48390 43252 48442
rect 42956 48388 43012 48390
rect 43036 48388 43092 48390
rect 43116 48388 43172 48390
rect 43196 48388 43252 48390
rect 42956 47354 43012 47356
rect 43036 47354 43092 47356
rect 43116 47354 43172 47356
rect 43196 47354 43252 47356
rect 42956 47302 43002 47354
rect 43002 47302 43012 47354
rect 43036 47302 43066 47354
rect 43066 47302 43078 47354
rect 43078 47302 43092 47354
rect 43116 47302 43130 47354
rect 43130 47302 43142 47354
rect 43142 47302 43172 47354
rect 43196 47302 43206 47354
rect 43206 47302 43252 47354
rect 42956 47300 43012 47302
rect 43036 47300 43092 47302
rect 43116 47300 43172 47302
rect 43196 47300 43252 47302
rect 42956 46266 43012 46268
rect 43036 46266 43092 46268
rect 43116 46266 43172 46268
rect 43196 46266 43252 46268
rect 42956 46214 43002 46266
rect 43002 46214 43012 46266
rect 43036 46214 43066 46266
rect 43066 46214 43078 46266
rect 43078 46214 43092 46266
rect 43116 46214 43130 46266
rect 43130 46214 43142 46266
rect 43142 46214 43172 46266
rect 43196 46214 43206 46266
rect 43206 46214 43252 46266
rect 42956 46212 43012 46214
rect 43036 46212 43092 46214
rect 43116 46212 43172 46214
rect 43196 46212 43252 46214
rect 42956 45178 43012 45180
rect 43036 45178 43092 45180
rect 43116 45178 43172 45180
rect 43196 45178 43252 45180
rect 42956 45126 43002 45178
rect 43002 45126 43012 45178
rect 43036 45126 43066 45178
rect 43066 45126 43078 45178
rect 43078 45126 43092 45178
rect 43116 45126 43130 45178
rect 43130 45126 43142 45178
rect 43142 45126 43172 45178
rect 43196 45126 43206 45178
rect 43206 45126 43252 45178
rect 42956 45124 43012 45126
rect 43036 45124 43092 45126
rect 43116 45124 43172 45126
rect 43196 45124 43252 45126
rect 42956 44090 43012 44092
rect 43036 44090 43092 44092
rect 43116 44090 43172 44092
rect 43196 44090 43252 44092
rect 42956 44038 43002 44090
rect 43002 44038 43012 44090
rect 43036 44038 43066 44090
rect 43066 44038 43078 44090
rect 43078 44038 43092 44090
rect 43116 44038 43130 44090
rect 43130 44038 43142 44090
rect 43142 44038 43172 44090
rect 43196 44038 43206 44090
rect 43206 44038 43252 44090
rect 42956 44036 43012 44038
rect 43036 44036 43092 44038
rect 43116 44036 43172 44038
rect 43196 44036 43252 44038
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 40590 19488 40646 19544
rect 42956 43002 43012 43004
rect 43036 43002 43092 43004
rect 43116 43002 43172 43004
rect 43196 43002 43252 43004
rect 42956 42950 43002 43002
rect 43002 42950 43012 43002
rect 43036 42950 43066 43002
rect 43066 42950 43078 43002
rect 43078 42950 43092 43002
rect 43116 42950 43130 43002
rect 43130 42950 43142 43002
rect 43142 42950 43172 43002
rect 43196 42950 43206 43002
rect 43206 42950 43252 43002
rect 42956 42948 43012 42950
rect 43036 42948 43092 42950
rect 43116 42948 43172 42950
rect 43196 42948 43252 42950
rect 42956 41914 43012 41916
rect 43036 41914 43092 41916
rect 43116 41914 43172 41916
rect 43196 41914 43252 41916
rect 42956 41862 43002 41914
rect 43002 41862 43012 41914
rect 43036 41862 43066 41914
rect 43066 41862 43078 41914
rect 43078 41862 43092 41914
rect 43116 41862 43130 41914
rect 43130 41862 43142 41914
rect 43142 41862 43172 41914
rect 43196 41862 43206 41914
rect 43206 41862 43252 41914
rect 42956 41860 43012 41862
rect 43036 41860 43092 41862
rect 43116 41860 43172 41862
rect 43196 41860 43252 41862
rect 42956 40826 43012 40828
rect 43036 40826 43092 40828
rect 43116 40826 43172 40828
rect 43196 40826 43252 40828
rect 42956 40774 43002 40826
rect 43002 40774 43012 40826
rect 43036 40774 43066 40826
rect 43066 40774 43078 40826
rect 43078 40774 43092 40826
rect 43116 40774 43130 40826
rect 43130 40774 43142 40826
rect 43142 40774 43172 40826
rect 43196 40774 43206 40826
rect 43206 40774 43252 40826
rect 42956 40772 43012 40774
rect 43036 40772 43092 40774
rect 43116 40772 43172 40774
rect 43196 40772 43252 40774
rect 42956 39738 43012 39740
rect 43036 39738 43092 39740
rect 43116 39738 43172 39740
rect 43196 39738 43252 39740
rect 42956 39686 43002 39738
rect 43002 39686 43012 39738
rect 43036 39686 43066 39738
rect 43066 39686 43078 39738
rect 43078 39686 43092 39738
rect 43116 39686 43130 39738
rect 43130 39686 43142 39738
rect 43142 39686 43172 39738
rect 43196 39686 43206 39738
rect 43206 39686 43252 39738
rect 42956 39684 43012 39686
rect 43036 39684 43092 39686
rect 43116 39684 43172 39686
rect 43196 39684 43252 39686
rect 42956 38650 43012 38652
rect 43036 38650 43092 38652
rect 43116 38650 43172 38652
rect 43196 38650 43252 38652
rect 42956 38598 43002 38650
rect 43002 38598 43012 38650
rect 43036 38598 43066 38650
rect 43066 38598 43078 38650
rect 43078 38598 43092 38650
rect 43116 38598 43130 38650
rect 43130 38598 43142 38650
rect 43142 38598 43172 38650
rect 43196 38598 43206 38650
rect 43206 38598 43252 38650
rect 42956 38596 43012 38598
rect 43036 38596 43092 38598
rect 43116 38596 43172 38598
rect 43196 38596 43252 38598
rect 42956 37562 43012 37564
rect 43036 37562 43092 37564
rect 43116 37562 43172 37564
rect 43196 37562 43252 37564
rect 42956 37510 43002 37562
rect 43002 37510 43012 37562
rect 43036 37510 43066 37562
rect 43066 37510 43078 37562
rect 43078 37510 43092 37562
rect 43116 37510 43130 37562
rect 43130 37510 43142 37562
rect 43142 37510 43172 37562
rect 43196 37510 43206 37562
rect 43206 37510 43252 37562
rect 42956 37508 43012 37510
rect 43036 37508 43092 37510
rect 43116 37508 43172 37510
rect 43196 37508 43252 37510
rect 42956 36474 43012 36476
rect 43036 36474 43092 36476
rect 43116 36474 43172 36476
rect 43196 36474 43252 36476
rect 42956 36422 43002 36474
rect 43002 36422 43012 36474
rect 43036 36422 43066 36474
rect 43066 36422 43078 36474
rect 43078 36422 43092 36474
rect 43116 36422 43130 36474
rect 43130 36422 43142 36474
rect 43142 36422 43172 36474
rect 43196 36422 43206 36474
rect 43206 36422 43252 36474
rect 42956 36420 43012 36422
rect 43036 36420 43092 36422
rect 43116 36420 43172 36422
rect 43196 36420 43252 36422
rect 42956 35386 43012 35388
rect 43036 35386 43092 35388
rect 43116 35386 43172 35388
rect 43196 35386 43252 35388
rect 42956 35334 43002 35386
rect 43002 35334 43012 35386
rect 43036 35334 43066 35386
rect 43066 35334 43078 35386
rect 43078 35334 43092 35386
rect 43116 35334 43130 35386
rect 43130 35334 43142 35386
rect 43142 35334 43172 35386
rect 43196 35334 43206 35386
rect 43206 35334 43252 35386
rect 42956 35332 43012 35334
rect 43036 35332 43092 35334
rect 43116 35332 43172 35334
rect 43196 35332 43252 35334
rect 42956 34298 43012 34300
rect 43036 34298 43092 34300
rect 43116 34298 43172 34300
rect 43196 34298 43252 34300
rect 42956 34246 43002 34298
rect 43002 34246 43012 34298
rect 43036 34246 43066 34298
rect 43066 34246 43078 34298
rect 43078 34246 43092 34298
rect 43116 34246 43130 34298
rect 43130 34246 43142 34298
rect 43142 34246 43172 34298
rect 43196 34246 43206 34298
rect 43206 34246 43252 34298
rect 42956 34244 43012 34246
rect 43036 34244 43092 34246
rect 43116 34244 43172 34246
rect 43196 34244 43252 34246
rect 42956 33210 43012 33212
rect 43036 33210 43092 33212
rect 43116 33210 43172 33212
rect 43196 33210 43252 33212
rect 42956 33158 43002 33210
rect 43002 33158 43012 33210
rect 43036 33158 43066 33210
rect 43066 33158 43078 33210
rect 43078 33158 43092 33210
rect 43116 33158 43130 33210
rect 43130 33158 43142 33210
rect 43142 33158 43172 33210
rect 43196 33158 43206 33210
rect 43206 33158 43252 33210
rect 42956 33156 43012 33158
rect 43036 33156 43092 33158
rect 43116 33156 43172 33158
rect 43196 33156 43252 33158
rect 42956 32122 43012 32124
rect 43036 32122 43092 32124
rect 43116 32122 43172 32124
rect 43196 32122 43252 32124
rect 42956 32070 43002 32122
rect 43002 32070 43012 32122
rect 43036 32070 43066 32122
rect 43066 32070 43078 32122
rect 43078 32070 43092 32122
rect 43116 32070 43130 32122
rect 43130 32070 43142 32122
rect 43142 32070 43172 32122
rect 43196 32070 43206 32122
rect 43206 32070 43252 32122
rect 42956 32068 43012 32070
rect 43036 32068 43092 32070
rect 43116 32068 43172 32070
rect 43196 32068 43252 32070
rect 42956 31034 43012 31036
rect 43036 31034 43092 31036
rect 43116 31034 43172 31036
rect 43196 31034 43252 31036
rect 42956 30982 43002 31034
rect 43002 30982 43012 31034
rect 43036 30982 43066 31034
rect 43066 30982 43078 31034
rect 43078 30982 43092 31034
rect 43116 30982 43130 31034
rect 43130 30982 43142 31034
rect 43142 30982 43172 31034
rect 43196 30982 43206 31034
rect 43206 30982 43252 31034
rect 42956 30980 43012 30982
rect 43036 30980 43092 30982
rect 43116 30980 43172 30982
rect 43196 30980 43252 30982
rect 42956 29946 43012 29948
rect 43036 29946 43092 29948
rect 43116 29946 43172 29948
rect 43196 29946 43252 29948
rect 42956 29894 43002 29946
rect 43002 29894 43012 29946
rect 43036 29894 43066 29946
rect 43066 29894 43078 29946
rect 43078 29894 43092 29946
rect 43116 29894 43130 29946
rect 43130 29894 43142 29946
rect 43142 29894 43172 29946
rect 43196 29894 43206 29946
rect 43206 29894 43252 29946
rect 42956 29892 43012 29894
rect 43036 29892 43092 29894
rect 43116 29892 43172 29894
rect 43196 29892 43252 29894
rect 42956 28858 43012 28860
rect 43036 28858 43092 28860
rect 43116 28858 43172 28860
rect 43196 28858 43252 28860
rect 42956 28806 43002 28858
rect 43002 28806 43012 28858
rect 43036 28806 43066 28858
rect 43066 28806 43078 28858
rect 43078 28806 43092 28858
rect 43116 28806 43130 28858
rect 43130 28806 43142 28858
rect 43142 28806 43172 28858
rect 43196 28806 43206 28858
rect 43206 28806 43252 28858
rect 42956 28804 43012 28806
rect 43036 28804 43092 28806
rect 43116 28804 43172 28806
rect 43196 28804 43252 28806
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 40498 8880 40554 8936
rect 40866 8472 40922 8528
rect 42956 27770 43012 27772
rect 43036 27770 43092 27772
rect 43116 27770 43172 27772
rect 43196 27770 43252 27772
rect 42956 27718 43002 27770
rect 43002 27718 43012 27770
rect 43036 27718 43066 27770
rect 43066 27718 43078 27770
rect 43078 27718 43092 27770
rect 43116 27718 43130 27770
rect 43130 27718 43142 27770
rect 43142 27718 43172 27770
rect 43196 27718 43206 27770
rect 43206 27718 43252 27770
rect 42956 27716 43012 27718
rect 43036 27716 43092 27718
rect 43116 27716 43172 27718
rect 43196 27716 43252 27718
rect 42956 26682 43012 26684
rect 43036 26682 43092 26684
rect 43116 26682 43172 26684
rect 43196 26682 43252 26684
rect 42956 26630 43002 26682
rect 43002 26630 43012 26682
rect 43036 26630 43066 26682
rect 43066 26630 43078 26682
rect 43078 26630 43092 26682
rect 43116 26630 43130 26682
rect 43130 26630 43142 26682
rect 43142 26630 43172 26682
rect 43196 26630 43206 26682
rect 43206 26630 43252 26682
rect 42956 26628 43012 26630
rect 43036 26628 43092 26630
rect 43116 26628 43172 26630
rect 43196 26628 43252 26630
rect 42956 25594 43012 25596
rect 43036 25594 43092 25596
rect 43116 25594 43172 25596
rect 43196 25594 43252 25596
rect 42956 25542 43002 25594
rect 43002 25542 43012 25594
rect 43036 25542 43066 25594
rect 43066 25542 43078 25594
rect 43078 25542 43092 25594
rect 43116 25542 43130 25594
rect 43130 25542 43142 25594
rect 43142 25542 43172 25594
rect 43196 25542 43206 25594
rect 43206 25542 43252 25594
rect 42956 25540 43012 25542
rect 43036 25540 43092 25542
rect 43116 25540 43172 25542
rect 43196 25540 43252 25542
rect 42982 25064 43038 25120
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 43902 19488 43958 19544
rect 49146 54576 49202 54632
rect 47956 53338 48012 53340
rect 48036 53338 48092 53340
rect 48116 53338 48172 53340
rect 48196 53338 48252 53340
rect 47956 53286 48002 53338
rect 48002 53286 48012 53338
rect 48036 53286 48066 53338
rect 48066 53286 48078 53338
rect 48078 53286 48092 53338
rect 48116 53286 48130 53338
rect 48130 53286 48142 53338
rect 48142 53286 48172 53338
rect 48196 53286 48206 53338
rect 48206 53286 48252 53338
rect 47956 53284 48012 53286
rect 48036 53284 48092 53286
rect 48116 53284 48172 53286
rect 48196 53284 48252 53286
rect 47956 52250 48012 52252
rect 48036 52250 48092 52252
rect 48116 52250 48172 52252
rect 48196 52250 48252 52252
rect 47956 52198 48002 52250
rect 48002 52198 48012 52250
rect 48036 52198 48066 52250
rect 48066 52198 48078 52250
rect 48078 52198 48092 52250
rect 48116 52198 48130 52250
rect 48130 52198 48142 52250
rect 48142 52198 48172 52250
rect 48196 52198 48206 52250
rect 48206 52198 48252 52250
rect 47956 52196 48012 52198
rect 48036 52196 48092 52198
rect 48116 52196 48172 52198
rect 48196 52196 48252 52198
rect 47956 51162 48012 51164
rect 48036 51162 48092 51164
rect 48116 51162 48172 51164
rect 48196 51162 48252 51164
rect 47956 51110 48002 51162
rect 48002 51110 48012 51162
rect 48036 51110 48066 51162
rect 48066 51110 48078 51162
rect 48078 51110 48092 51162
rect 48116 51110 48130 51162
rect 48130 51110 48142 51162
rect 48142 51110 48172 51162
rect 48196 51110 48206 51162
rect 48206 51110 48252 51162
rect 47956 51108 48012 51110
rect 48036 51108 48092 51110
rect 48116 51108 48172 51110
rect 48196 51108 48252 51110
rect 47956 50074 48012 50076
rect 48036 50074 48092 50076
rect 48116 50074 48172 50076
rect 48196 50074 48252 50076
rect 47956 50022 48002 50074
rect 48002 50022 48012 50074
rect 48036 50022 48066 50074
rect 48066 50022 48078 50074
rect 48078 50022 48092 50074
rect 48116 50022 48130 50074
rect 48130 50022 48142 50074
rect 48142 50022 48172 50074
rect 48196 50022 48206 50074
rect 48206 50022 48252 50074
rect 47956 50020 48012 50022
rect 48036 50020 48092 50022
rect 48116 50020 48172 50022
rect 48196 50020 48252 50022
rect 47956 48986 48012 48988
rect 48036 48986 48092 48988
rect 48116 48986 48172 48988
rect 48196 48986 48252 48988
rect 47956 48934 48002 48986
rect 48002 48934 48012 48986
rect 48036 48934 48066 48986
rect 48066 48934 48078 48986
rect 48078 48934 48092 48986
rect 48116 48934 48130 48986
rect 48130 48934 48142 48986
rect 48142 48934 48172 48986
rect 48196 48934 48206 48986
rect 48206 48934 48252 48986
rect 47956 48932 48012 48934
rect 48036 48932 48092 48934
rect 48116 48932 48172 48934
rect 48196 48932 48252 48934
rect 47956 47898 48012 47900
rect 48036 47898 48092 47900
rect 48116 47898 48172 47900
rect 48196 47898 48252 47900
rect 47956 47846 48002 47898
rect 48002 47846 48012 47898
rect 48036 47846 48066 47898
rect 48066 47846 48078 47898
rect 48078 47846 48092 47898
rect 48116 47846 48130 47898
rect 48130 47846 48142 47898
rect 48142 47846 48172 47898
rect 48196 47846 48206 47898
rect 48206 47846 48252 47898
rect 47956 47844 48012 47846
rect 48036 47844 48092 47846
rect 48116 47844 48172 47846
rect 48196 47844 48252 47846
rect 47956 46810 48012 46812
rect 48036 46810 48092 46812
rect 48116 46810 48172 46812
rect 48196 46810 48252 46812
rect 47956 46758 48002 46810
rect 48002 46758 48012 46810
rect 48036 46758 48066 46810
rect 48066 46758 48078 46810
rect 48078 46758 48092 46810
rect 48116 46758 48130 46810
rect 48130 46758 48142 46810
rect 48142 46758 48172 46810
rect 48196 46758 48206 46810
rect 48206 46758 48252 46810
rect 47956 46756 48012 46758
rect 48036 46756 48092 46758
rect 48116 46756 48172 46758
rect 48196 46756 48252 46758
rect 47956 45722 48012 45724
rect 48036 45722 48092 45724
rect 48116 45722 48172 45724
rect 48196 45722 48252 45724
rect 47956 45670 48002 45722
rect 48002 45670 48012 45722
rect 48036 45670 48066 45722
rect 48066 45670 48078 45722
rect 48078 45670 48092 45722
rect 48116 45670 48130 45722
rect 48130 45670 48142 45722
rect 48142 45670 48172 45722
rect 48196 45670 48206 45722
rect 48206 45670 48252 45722
rect 47956 45668 48012 45670
rect 48036 45668 48092 45670
rect 48116 45668 48172 45670
rect 48196 45668 48252 45670
rect 47956 44634 48012 44636
rect 48036 44634 48092 44636
rect 48116 44634 48172 44636
rect 48196 44634 48252 44636
rect 47956 44582 48002 44634
rect 48002 44582 48012 44634
rect 48036 44582 48066 44634
rect 48066 44582 48078 44634
rect 48078 44582 48092 44634
rect 48116 44582 48130 44634
rect 48130 44582 48142 44634
rect 48142 44582 48172 44634
rect 48196 44582 48206 44634
rect 48206 44582 48252 44634
rect 47956 44580 48012 44582
rect 48036 44580 48092 44582
rect 48116 44580 48172 44582
rect 48196 44580 48252 44582
rect 47956 43546 48012 43548
rect 48036 43546 48092 43548
rect 48116 43546 48172 43548
rect 48196 43546 48252 43548
rect 47956 43494 48002 43546
rect 48002 43494 48012 43546
rect 48036 43494 48066 43546
rect 48066 43494 48078 43546
rect 48078 43494 48092 43546
rect 48116 43494 48130 43546
rect 48130 43494 48142 43546
rect 48142 43494 48172 43546
rect 48196 43494 48206 43546
rect 48206 43494 48252 43546
rect 47956 43492 48012 43494
rect 48036 43492 48092 43494
rect 48116 43492 48172 43494
rect 48196 43492 48252 43494
rect 47956 42458 48012 42460
rect 48036 42458 48092 42460
rect 48116 42458 48172 42460
rect 48196 42458 48252 42460
rect 47956 42406 48002 42458
rect 48002 42406 48012 42458
rect 48036 42406 48066 42458
rect 48066 42406 48078 42458
rect 48078 42406 48092 42458
rect 48116 42406 48130 42458
rect 48130 42406 48142 42458
rect 48142 42406 48172 42458
rect 48196 42406 48206 42458
rect 48206 42406 48252 42458
rect 47956 42404 48012 42406
rect 48036 42404 48092 42406
rect 48116 42404 48172 42406
rect 48196 42404 48252 42406
rect 47956 41370 48012 41372
rect 48036 41370 48092 41372
rect 48116 41370 48172 41372
rect 48196 41370 48252 41372
rect 47956 41318 48002 41370
rect 48002 41318 48012 41370
rect 48036 41318 48066 41370
rect 48066 41318 48078 41370
rect 48078 41318 48092 41370
rect 48116 41318 48130 41370
rect 48130 41318 48142 41370
rect 48142 41318 48172 41370
rect 48196 41318 48206 41370
rect 48206 41318 48252 41370
rect 47956 41316 48012 41318
rect 48036 41316 48092 41318
rect 48116 41316 48172 41318
rect 48196 41316 48252 41318
rect 47956 40282 48012 40284
rect 48036 40282 48092 40284
rect 48116 40282 48172 40284
rect 48196 40282 48252 40284
rect 47956 40230 48002 40282
rect 48002 40230 48012 40282
rect 48036 40230 48066 40282
rect 48066 40230 48078 40282
rect 48078 40230 48092 40282
rect 48116 40230 48130 40282
rect 48130 40230 48142 40282
rect 48142 40230 48172 40282
rect 48196 40230 48206 40282
rect 48206 40230 48252 40282
rect 47956 40228 48012 40230
rect 48036 40228 48092 40230
rect 48116 40228 48172 40230
rect 48196 40228 48252 40230
rect 47956 39194 48012 39196
rect 48036 39194 48092 39196
rect 48116 39194 48172 39196
rect 48196 39194 48252 39196
rect 47956 39142 48002 39194
rect 48002 39142 48012 39194
rect 48036 39142 48066 39194
rect 48066 39142 48078 39194
rect 48078 39142 48092 39194
rect 48116 39142 48130 39194
rect 48130 39142 48142 39194
rect 48142 39142 48172 39194
rect 48196 39142 48206 39194
rect 48206 39142 48252 39194
rect 47956 39140 48012 39142
rect 48036 39140 48092 39142
rect 48116 39140 48172 39142
rect 48196 39140 48252 39142
rect 47956 38106 48012 38108
rect 48036 38106 48092 38108
rect 48116 38106 48172 38108
rect 48196 38106 48252 38108
rect 47956 38054 48002 38106
rect 48002 38054 48012 38106
rect 48036 38054 48066 38106
rect 48066 38054 48078 38106
rect 48078 38054 48092 38106
rect 48116 38054 48130 38106
rect 48130 38054 48142 38106
rect 48142 38054 48172 38106
rect 48196 38054 48206 38106
rect 48206 38054 48252 38106
rect 47956 38052 48012 38054
rect 48036 38052 48092 38054
rect 48116 38052 48172 38054
rect 48196 38052 48252 38054
rect 47956 37018 48012 37020
rect 48036 37018 48092 37020
rect 48116 37018 48172 37020
rect 48196 37018 48252 37020
rect 47956 36966 48002 37018
rect 48002 36966 48012 37018
rect 48036 36966 48066 37018
rect 48066 36966 48078 37018
rect 48078 36966 48092 37018
rect 48116 36966 48130 37018
rect 48130 36966 48142 37018
rect 48142 36966 48172 37018
rect 48196 36966 48206 37018
rect 48206 36966 48252 37018
rect 47956 36964 48012 36966
rect 48036 36964 48092 36966
rect 48116 36964 48172 36966
rect 48196 36964 48252 36966
rect 47956 35930 48012 35932
rect 48036 35930 48092 35932
rect 48116 35930 48172 35932
rect 48196 35930 48252 35932
rect 47956 35878 48002 35930
rect 48002 35878 48012 35930
rect 48036 35878 48066 35930
rect 48066 35878 48078 35930
rect 48078 35878 48092 35930
rect 48116 35878 48130 35930
rect 48130 35878 48142 35930
rect 48142 35878 48172 35930
rect 48196 35878 48206 35930
rect 48206 35878 48252 35930
rect 47956 35876 48012 35878
rect 48036 35876 48092 35878
rect 48116 35876 48172 35878
rect 48196 35876 48252 35878
rect 47956 34842 48012 34844
rect 48036 34842 48092 34844
rect 48116 34842 48172 34844
rect 48196 34842 48252 34844
rect 47956 34790 48002 34842
rect 48002 34790 48012 34842
rect 48036 34790 48066 34842
rect 48066 34790 48078 34842
rect 48078 34790 48092 34842
rect 48116 34790 48130 34842
rect 48130 34790 48142 34842
rect 48142 34790 48172 34842
rect 48196 34790 48206 34842
rect 48206 34790 48252 34842
rect 47956 34788 48012 34790
rect 48036 34788 48092 34790
rect 48116 34788 48172 34790
rect 48196 34788 48252 34790
rect 47956 33754 48012 33756
rect 48036 33754 48092 33756
rect 48116 33754 48172 33756
rect 48196 33754 48252 33756
rect 47956 33702 48002 33754
rect 48002 33702 48012 33754
rect 48036 33702 48066 33754
rect 48066 33702 48078 33754
rect 48078 33702 48092 33754
rect 48116 33702 48130 33754
rect 48130 33702 48142 33754
rect 48142 33702 48172 33754
rect 48196 33702 48206 33754
rect 48206 33702 48252 33754
rect 47956 33700 48012 33702
rect 48036 33700 48092 33702
rect 48116 33700 48172 33702
rect 48196 33700 48252 33702
rect 45558 25100 45560 25120
rect 45560 25100 45612 25120
rect 45612 25100 45614 25120
rect 45558 25064 45614 25100
rect 47956 32666 48012 32668
rect 48036 32666 48092 32668
rect 48116 32666 48172 32668
rect 48196 32666 48252 32668
rect 47956 32614 48002 32666
rect 48002 32614 48012 32666
rect 48036 32614 48066 32666
rect 48066 32614 48078 32666
rect 48078 32614 48092 32666
rect 48116 32614 48130 32666
rect 48130 32614 48142 32666
rect 48142 32614 48172 32666
rect 48196 32614 48206 32666
rect 48206 32614 48252 32666
rect 47956 32612 48012 32614
rect 48036 32612 48092 32614
rect 48116 32612 48172 32614
rect 48196 32612 48252 32614
rect 47956 31578 48012 31580
rect 48036 31578 48092 31580
rect 48116 31578 48172 31580
rect 48196 31578 48252 31580
rect 47956 31526 48002 31578
rect 48002 31526 48012 31578
rect 48036 31526 48066 31578
rect 48066 31526 48078 31578
rect 48078 31526 48092 31578
rect 48116 31526 48130 31578
rect 48130 31526 48142 31578
rect 48142 31526 48172 31578
rect 48196 31526 48206 31578
rect 48206 31526 48252 31578
rect 47956 31524 48012 31526
rect 48036 31524 48092 31526
rect 48116 31524 48172 31526
rect 48196 31524 48252 31526
rect 47956 30490 48012 30492
rect 48036 30490 48092 30492
rect 48116 30490 48172 30492
rect 48196 30490 48252 30492
rect 47956 30438 48002 30490
rect 48002 30438 48012 30490
rect 48036 30438 48066 30490
rect 48066 30438 48078 30490
rect 48078 30438 48092 30490
rect 48116 30438 48130 30490
rect 48130 30438 48142 30490
rect 48142 30438 48172 30490
rect 48196 30438 48206 30490
rect 48206 30438 48252 30490
rect 47956 30436 48012 30438
rect 48036 30436 48092 30438
rect 48116 30436 48172 30438
rect 48196 30436 48252 30438
rect 47956 29402 48012 29404
rect 48036 29402 48092 29404
rect 48116 29402 48172 29404
rect 48196 29402 48252 29404
rect 47956 29350 48002 29402
rect 48002 29350 48012 29402
rect 48036 29350 48066 29402
rect 48066 29350 48078 29402
rect 48078 29350 48092 29402
rect 48116 29350 48130 29402
rect 48130 29350 48142 29402
rect 48142 29350 48172 29402
rect 48196 29350 48206 29402
rect 48206 29350 48252 29402
rect 47956 29348 48012 29350
rect 48036 29348 48092 29350
rect 48116 29348 48172 29350
rect 48196 29348 48252 29350
rect 47956 28314 48012 28316
rect 48036 28314 48092 28316
rect 48116 28314 48172 28316
rect 48196 28314 48252 28316
rect 47956 28262 48002 28314
rect 48002 28262 48012 28314
rect 48036 28262 48066 28314
rect 48066 28262 48078 28314
rect 48078 28262 48092 28314
rect 48116 28262 48130 28314
rect 48130 28262 48142 28314
rect 48142 28262 48172 28314
rect 48196 28262 48206 28314
rect 48206 28262 48252 28314
rect 47956 28260 48012 28262
rect 48036 28260 48092 28262
rect 48116 28260 48172 28262
rect 48196 28260 48252 28262
rect 47956 27226 48012 27228
rect 48036 27226 48092 27228
rect 48116 27226 48172 27228
rect 48196 27226 48252 27228
rect 47956 27174 48002 27226
rect 48002 27174 48012 27226
rect 48036 27174 48066 27226
rect 48066 27174 48078 27226
rect 48078 27174 48092 27226
rect 48116 27174 48130 27226
rect 48130 27174 48142 27226
rect 48142 27174 48172 27226
rect 48196 27174 48206 27226
rect 48206 27174 48252 27226
rect 47956 27172 48012 27174
rect 48036 27172 48092 27174
rect 48116 27172 48172 27174
rect 48196 27172 48252 27174
rect 47956 26138 48012 26140
rect 48036 26138 48092 26140
rect 48116 26138 48172 26140
rect 48196 26138 48252 26140
rect 47956 26086 48002 26138
rect 48002 26086 48012 26138
rect 48036 26086 48066 26138
rect 48066 26086 48078 26138
rect 48078 26086 48092 26138
rect 48116 26086 48130 26138
rect 48130 26086 48142 26138
rect 48142 26086 48172 26138
rect 48196 26086 48206 26138
rect 48206 26086 48252 26138
rect 47956 26084 48012 26086
rect 48036 26084 48092 26086
rect 48116 26084 48172 26086
rect 48196 26084 48252 26086
rect 47956 25050 48012 25052
rect 48036 25050 48092 25052
rect 48116 25050 48172 25052
rect 48196 25050 48252 25052
rect 47956 24998 48002 25050
rect 48002 24998 48012 25050
rect 48036 24998 48066 25050
rect 48066 24998 48078 25050
rect 48078 24998 48092 25050
rect 48116 24998 48130 25050
rect 48130 24998 48142 25050
rect 48142 24998 48172 25050
rect 48196 24998 48206 25050
rect 48206 24998 48252 25050
rect 47956 24996 48012 24998
rect 48036 24996 48092 24998
rect 48116 24996 48172 24998
rect 48196 24996 48252 24998
rect 48502 26016 48558 26072
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 49054 53760 49110 53816
rect 49054 52944 49110 53000
rect 48962 52128 49018 52184
rect 48962 51332 49018 51368
rect 48962 51312 48964 51332
rect 48964 51312 49016 51332
rect 49016 51312 49018 51332
rect 48962 50496 49018 50552
rect 49146 49680 49202 49736
rect 49146 48864 49202 48920
rect 49146 48068 49202 48104
rect 49146 48048 49148 48068
rect 49148 48048 49200 48068
rect 49200 48048 49202 48068
rect 49330 47232 49386 47288
rect 49330 46416 49386 46472
rect 49330 45600 49386 45656
rect 49330 44820 49332 44840
rect 49332 44820 49384 44840
rect 49384 44820 49386 44840
rect 49330 44784 49386 44820
rect 49146 43968 49202 44024
rect 49146 43152 49202 43208
rect 49146 42336 49202 42392
rect 49146 41540 49202 41576
rect 49146 41520 49148 41540
rect 49148 41520 49200 41540
rect 49200 41520 49202 41540
rect 49146 37440 49202 37496
rect 49146 36624 49202 36680
rect 49146 25236 49148 25256
rect 49148 25236 49200 25256
rect 49200 25236 49202 25256
rect 49146 25200 49202 25236
rect 49146 24384 49202 24440
rect 49146 23604 49148 23624
rect 49148 23604 49200 23624
rect 49200 23604 49202 23624
rect 49146 23568 49202 23604
rect 49146 22752 49202 22808
rect 49146 21972 49148 21992
rect 49148 21972 49200 21992
rect 49200 21972 49202 21992
rect 49146 21936 49202 21972
rect 49146 21120 49202 21176
rect 49146 20340 49148 20360
rect 49148 20340 49200 20360
rect 49200 20340 49202 20360
rect 49146 20304 49202 20340
rect 49146 19488 49202 19544
rect 49146 18708 49148 18728
rect 49148 18708 49200 18728
rect 49200 18708 49202 18728
rect 49146 18672 49202 18708
rect 49146 17856 49202 17912
rect 49146 17076 49148 17096
rect 49148 17076 49200 17096
rect 49200 17076 49202 17096
rect 49146 17040 49202 17076
rect 49146 16224 49202 16280
rect 49146 15444 49148 15464
rect 49148 15444 49200 15464
rect 49200 15444 49202 15464
rect 49146 15408 49202 15444
rect 49146 14592 49202 14648
rect 49330 40704 49386 40760
rect 49330 39888 49386 39944
rect 49330 39072 49386 39128
rect 49330 38292 49332 38312
rect 49332 38292 49384 38312
rect 49384 38292 49386 38312
rect 49330 38256 49386 38292
rect 49330 35808 49386 35864
rect 49330 35028 49332 35048
rect 49332 35028 49384 35048
rect 49384 35028 49386 35048
rect 49330 34992 49386 35028
rect 49330 34176 49386 34232
rect 49330 33360 49386 33416
rect 49330 32544 49386 32600
rect 49330 31764 49332 31784
rect 49332 31764 49384 31784
rect 49384 31764 49386 31784
rect 49330 31728 49386 31764
rect 49330 30912 49386 30968
rect 49330 30096 49386 30152
rect 49330 29280 49386 29336
rect 49330 28500 49332 28520
rect 49332 28500 49384 28520
rect 49384 28500 49386 28520
rect 49330 28464 49386 28500
rect 49330 27648 49386 27704
rect 49330 26832 49386 26888
rect 49974 29552 50030 29608
rect 50434 25744 50490 25800
rect 49146 13812 49148 13832
rect 49148 13812 49200 13832
rect 49200 13812 49202 13832
rect 49146 13776 49202 13812
rect 49146 12960 49202 13016
rect 49146 12180 49148 12200
rect 49148 12180 49200 12200
rect 49200 12180 49202 12200
rect 49146 12144 49202 12180
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 49146 11328 49202 11384
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49146 10548 49148 10568
rect 49148 10548 49200 10568
rect 49200 10548 49202 10568
rect 49146 10512 49202 10548
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 49146 9696 49202 9752
rect 49146 8900 49202 8936
rect 49146 8880 49148 8900
rect 49148 8880 49200 8900
rect 49200 8880 49202 8900
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 49146 8064 49202 8120
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 7284 49148 7304
rect 49148 7284 49200 7304
rect 49200 7284 49202 7304
rect 49146 7248 49202 7284
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 49146 6432 49202 6488
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 5636 49202 5672
rect 49146 5616 49148 5636
rect 49148 5616 49200 5636
rect 49200 5616 49202 5636
rect 49146 4800 49202 4856
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47858 2352 47914 2408
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
rect 49146 4020 49148 4040
rect 49148 4020 49200 4040
rect 49200 4020 49202 4040
rect 49146 3984 49202 4020
rect 49146 3168 49202 3224
rect 49238 1536 49294 1592
rect 48686 720 48742 776
<< metal3 >>
rect 48405 56266 48471 56269
rect 50200 56266 51000 56296
rect 48405 56264 51000 56266
rect 48405 56208 48410 56264
rect 48466 56208 51000 56264
rect 48405 56206 51000 56208
rect 48405 56203 48471 56206
rect 50200 56176 51000 56206
rect 48221 55450 48287 55453
rect 50200 55450 51000 55480
rect 48221 55448 51000 55450
rect 48221 55392 48226 55448
rect 48282 55392 51000 55448
rect 48221 55390 51000 55392
rect 48221 55387 48287 55390
rect 50200 55360 51000 55390
rect 49141 54634 49207 54637
rect 50200 54634 51000 54664
rect 49141 54632 51000 54634
rect 49141 54576 49146 54632
rect 49202 54576 51000 54632
rect 49141 54574 51000 54576
rect 49141 54571 49207 54574
rect 50200 54544 51000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 27946 54432 28262 54433
rect 27946 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28262 54432
rect 27946 54367 28262 54368
rect 37946 54432 38262 54433
rect 37946 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38262 54432
rect 37946 54367 38262 54368
rect 47946 54432 48262 54433
rect 47946 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48262 54432
rect 47946 54367 48262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 32946 53888 33262 53889
rect 32946 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33262 53888
rect 32946 53823 33262 53824
rect 42946 53888 43262 53889
rect 42946 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43262 53888
rect 42946 53823 43262 53824
rect 49049 53818 49115 53821
rect 50200 53818 51000 53848
rect 49049 53816 51000 53818
rect 49049 53760 49054 53816
rect 49110 53760 51000 53816
rect 49049 53758 51000 53760
rect 49049 53755 49115 53758
rect 50200 53728 51000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 27946 53344 28262 53345
rect 27946 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28262 53344
rect 27946 53279 28262 53280
rect 37946 53344 38262 53345
rect 37946 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38262 53344
rect 37946 53279 38262 53280
rect 47946 53344 48262 53345
rect 47946 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48262 53344
rect 47946 53279 48262 53280
rect 49049 53002 49115 53005
rect 50200 53002 51000 53032
rect 49049 53000 51000 53002
rect 49049 52944 49054 53000
rect 49110 52944 51000 53000
rect 49049 52942 51000 52944
rect 49049 52939 49115 52942
rect 50200 52912 51000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 32946 52800 33262 52801
rect 32946 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33262 52800
rect 32946 52735 33262 52736
rect 42946 52800 43262 52801
rect 42946 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43262 52800
rect 42946 52735 43262 52736
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 27946 52256 28262 52257
rect 27946 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28262 52256
rect 27946 52191 28262 52192
rect 37946 52256 38262 52257
rect 37946 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38262 52256
rect 37946 52191 38262 52192
rect 47946 52256 48262 52257
rect 47946 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48262 52256
rect 47946 52191 48262 52192
rect 48957 52186 49023 52189
rect 50200 52186 51000 52216
rect 48957 52184 51000 52186
rect 48957 52128 48962 52184
rect 49018 52128 51000 52184
rect 48957 52126 51000 52128
rect 48957 52123 49023 52126
rect 50200 52096 51000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 32946 51712 33262 51713
rect 32946 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33262 51712
rect 32946 51647 33262 51648
rect 42946 51712 43262 51713
rect 42946 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43262 51712
rect 42946 51647 43262 51648
rect 48957 51370 49023 51373
rect 50200 51370 51000 51400
rect 48957 51368 51000 51370
rect 48957 51312 48962 51368
rect 49018 51312 51000 51368
rect 48957 51310 51000 51312
rect 48957 51307 49023 51310
rect 50200 51280 51000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 27946 51168 28262 51169
rect 27946 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28262 51168
rect 27946 51103 28262 51104
rect 37946 51168 38262 51169
rect 37946 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38262 51168
rect 37946 51103 38262 51104
rect 47946 51168 48262 51169
rect 47946 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48262 51168
rect 47946 51103 48262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 32946 50624 33262 50625
rect 32946 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33262 50624
rect 32946 50559 33262 50560
rect 42946 50624 43262 50625
rect 42946 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43262 50624
rect 42946 50559 43262 50560
rect 48957 50554 49023 50557
rect 50200 50554 51000 50584
rect 48957 50552 51000 50554
rect 48957 50496 48962 50552
rect 49018 50496 51000 50552
rect 48957 50494 51000 50496
rect 48957 50491 49023 50494
rect 50200 50464 51000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 27946 50080 28262 50081
rect 27946 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28262 50080
rect 27946 50015 28262 50016
rect 37946 50080 38262 50081
rect 37946 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38262 50080
rect 37946 50015 38262 50016
rect 47946 50080 48262 50081
rect 47946 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48262 50080
rect 47946 50015 48262 50016
rect 49141 49738 49207 49741
rect 50200 49738 51000 49768
rect 49141 49736 51000 49738
rect 49141 49680 49146 49736
rect 49202 49680 51000 49736
rect 49141 49678 51000 49680
rect 49141 49675 49207 49678
rect 50200 49648 51000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 32946 49536 33262 49537
rect 32946 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33262 49536
rect 32946 49471 33262 49472
rect 42946 49536 43262 49537
rect 42946 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43262 49536
rect 42946 49471 43262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 27946 48992 28262 48993
rect 27946 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28262 48992
rect 27946 48927 28262 48928
rect 37946 48992 38262 48993
rect 37946 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38262 48992
rect 37946 48927 38262 48928
rect 47946 48992 48262 48993
rect 47946 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48262 48992
rect 47946 48927 48262 48928
rect 49141 48922 49207 48925
rect 50200 48922 51000 48952
rect 49141 48920 51000 48922
rect 49141 48864 49146 48920
rect 49202 48864 51000 48920
rect 49141 48862 51000 48864
rect 49141 48859 49207 48862
rect 50200 48832 51000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 32946 48448 33262 48449
rect 32946 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33262 48448
rect 32946 48383 33262 48384
rect 42946 48448 43262 48449
rect 42946 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43262 48448
rect 42946 48383 43262 48384
rect 49141 48106 49207 48109
rect 50200 48106 51000 48136
rect 49141 48104 51000 48106
rect 49141 48048 49146 48104
rect 49202 48048 51000 48104
rect 49141 48046 51000 48048
rect 49141 48043 49207 48046
rect 50200 48016 51000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 27946 47904 28262 47905
rect 27946 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28262 47904
rect 27946 47839 28262 47840
rect 37946 47904 38262 47905
rect 37946 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38262 47904
rect 37946 47839 38262 47840
rect 47946 47904 48262 47905
rect 47946 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48262 47904
rect 47946 47839 48262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 32946 47360 33262 47361
rect 32946 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33262 47360
rect 32946 47295 33262 47296
rect 42946 47360 43262 47361
rect 42946 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43262 47360
rect 42946 47295 43262 47296
rect 49325 47290 49391 47293
rect 50200 47290 51000 47320
rect 49325 47288 51000 47290
rect 49325 47232 49330 47288
rect 49386 47232 51000 47288
rect 49325 47230 51000 47232
rect 49325 47227 49391 47230
rect 50200 47200 51000 47230
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 27946 46816 28262 46817
rect 27946 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28262 46816
rect 27946 46751 28262 46752
rect 37946 46816 38262 46817
rect 37946 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38262 46816
rect 37946 46751 38262 46752
rect 47946 46816 48262 46817
rect 47946 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48262 46816
rect 47946 46751 48262 46752
rect 49325 46474 49391 46477
rect 50200 46474 51000 46504
rect 49325 46472 51000 46474
rect 49325 46416 49330 46472
rect 49386 46416 51000 46472
rect 49325 46414 51000 46416
rect 49325 46411 49391 46414
rect 50200 46384 51000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 32946 46272 33262 46273
rect 32946 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33262 46272
rect 32946 46207 33262 46208
rect 42946 46272 43262 46273
rect 42946 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43262 46272
rect 42946 46207 43262 46208
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 27946 45728 28262 45729
rect 27946 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28262 45728
rect 27946 45663 28262 45664
rect 37946 45728 38262 45729
rect 37946 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38262 45728
rect 37946 45663 38262 45664
rect 47946 45728 48262 45729
rect 47946 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48262 45728
rect 47946 45663 48262 45664
rect 49325 45658 49391 45661
rect 50200 45658 51000 45688
rect 49325 45656 51000 45658
rect 49325 45600 49330 45656
rect 49386 45600 51000 45656
rect 49325 45598 51000 45600
rect 49325 45595 49391 45598
rect 50200 45568 51000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 32946 45184 33262 45185
rect 32946 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33262 45184
rect 32946 45119 33262 45120
rect 42946 45184 43262 45185
rect 42946 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43262 45184
rect 42946 45119 43262 45120
rect 49325 44842 49391 44845
rect 50200 44842 51000 44872
rect 49325 44840 51000 44842
rect 49325 44784 49330 44840
rect 49386 44784 51000 44840
rect 49325 44782 51000 44784
rect 49325 44779 49391 44782
rect 50200 44752 51000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 27946 44640 28262 44641
rect 27946 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28262 44640
rect 27946 44575 28262 44576
rect 37946 44640 38262 44641
rect 37946 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38262 44640
rect 37946 44575 38262 44576
rect 47946 44640 48262 44641
rect 47946 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48262 44640
rect 47946 44575 48262 44576
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 32946 44096 33262 44097
rect 32946 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33262 44096
rect 32946 44031 33262 44032
rect 42946 44096 43262 44097
rect 42946 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43262 44096
rect 42946 44031 43262 44032
rect 49141 44026 49207 44029
rect 50200 44026 51000 44056
rect 49141 44024 51000 44026
rect 49141 43968 49146 44024
rect 49202 43968 51000 44024
rect 49141 43966 51000 43968
rect 49141 43963 49207 43966
rect 50200 43936 51000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 27946 43552 28262 43553
rect 27946 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28262 43552
rect 27946 43487 28262 43488
rect 37946 43552 38262 43553
rect 37946 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38262 43552
rect 37946 43487 38262 43488
rect 47946 43552 48262 43553
rect 47946 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48262 43552
rect 47946 43487 48262 43488
rect 49141 43210 49207 43213
rect 50200 43210 51000 43240
rect 49141 43208 51000 43210
rect 49141 43152 49146 43208
rect 49202 43152 51000 43208
rect 49141 43150 51000 43152
rect 49141 43147 49207 43150
rect 50200 43120 51000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 32946 43008 33262 43009
rect 32946 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33262 43008
rect 32946 42943 33262 42944
rect 42946 43008 43262 43009
rect 42946 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43262 43008
rect 42946 42943 43262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 27946 42464 28262 42465
rect 27946 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28262 42464
rect 27946 42399 28262 42400
rect 37946 42464 38262 42465
rect 37946 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38262 42464
rect 37946 42399 38262 42400
rect 47946 42464 48262 42465
rect 47946 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48262 42464
rect 47946 42399 48262 42400
rect 49141 42394 49207 42397
rect 50200 42394 51000 42424
rect 49141 42392 51000 42394
rect 49141 42336 49146 42392
rect 49202 42336 51000 42392
rect 49141 42334 51000 42336
rect 49141 42331 49207 42334
rect 50200 42304 51000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 32946 41920 33262 41921
rect 32946 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33262 41920
rect 32946 41855 33262 41856
rect 42946 41920 43262 41921
rect 42946 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43262 41920
rect 42946 41855 43262 41856
rect 49141 41578 49207 41581
rect 50200 41578 51000 41608
rect 49141 41576 51000 41578
rect 49141 41520 49146 41576
rect 49202 41520 51000 41576
rect 49141 41518 51000 41520
rect 49141 41515 49207 41518
rect 50200 41488 51000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 27946 41376 28262 41377
rect 27946 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28262 41376
rect 27946 41311 28262 41312
rect 37946 41376 38262 41377
rect 37946 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38262 41376
rect 37946 41311 38262 41312
rect 47946 41376 48262 41377
rect 47946 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48262 41376
rect 47946 41311 48262 41312
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 32946 40832 33262 40833
rect 32946 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33262 40832
rect 32946 40767 33262 40768
rect 42946 40832 43262 40833
rect 42946 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43262 40832
rect 42946 40767 43262 40768
rect 49325 40762 49391 40765
rect 50200 40762 51000 40792
rect 49325 40760 51000 40762
rect 49325 40704 49330 40760
rect 49386 40704 51000 40760
rect 49325 40702 51000 40704
rect 49325 40699 49391 40702
rect 50200 40672 51000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 27946 40288 28262 40289
rect 27946 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28262 40288
rect 27946 40223 28262 40224
rect 37946 40288 38262 40289
rect 37946 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38262 40288
rect 37946 40223 38262 40224
rect 47946 40288 48262 40289
rect 47946 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48262 40288
rect 47946 40223 48262 40224
rect 49325 39946 49391 39949
rect 50200 39946 51000 39976
rect 49325 39944 51000 39946
rect 49325 39888 49330 39944
rect 49386 39888 51000 39944
rect 49325 39886 51000 39888
rect 49325 39883 49391 39886
rect 50200 39856 51000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 32946 39744 33262 39745
rect 32946 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33262 39744
rect 32946 39679 33262 39680
rect 42946 39744 43262 39745
rect 42946 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43262 39744
rect 42946 39679 43262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 27946 39200 28262 39201
rect 27946 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28262 39200
rect 27946 39135 28262 39136
rect 37946 39200 38262 39201
rect 37946 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38262 39200
rect 37946 39135 38262 39136
rect 47946 39200 48262 39201
rect 47946 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48262 39200
rect 47946 39135 48262 39136
rect 49325 39130 49391 39133
rect 50200 39130 51000 39160
rect 49325 39128 51000 39130
rect 49325 39072 49330 39128
rect 49386 39072 51000 39128
rect 49325 39070 51000 39072
rect 49325 39067 49391 39070
rect 50200 39040 51000 39070
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 32946 38656 33262 38657
rect 32946 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33262 38656
rect 32946 38591 33262 38592
rect 42946 38656 43262 38657
rect 42946 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43262 38656
rect 42946 38591 43262 38592
rect 49325 38314 49391 38317
rect 50200 38314 51000 38344
rect 49325 38312 51000 38314
rect 49325 38256 49330 38312
rect 49386 38256 51000 38312
rect 49325 38254 51000 38256
rect 49325 38251 49391 38254
rect 50200 38224 51000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 27946 38112 28262 38113
rect 27946 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28262 38112
rect 27946 38047 28262 38048
rect 37946 38112 38262 38113
rect 37946 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38262 38112
rect 37946 38047 38262 38048
rect 47946 38112 48262 38113
rect 47946 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48262 38112
rect 47946 38047 48262 38048
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 32946 37568 33262 37569
rect 32946 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33262 37568
rect 32946 37503 33262 37504
rect 42946 37568 43262 37569
rect 42946 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43262 37568
rect 42946 37503 43262 37504
rect 49141 37498 49207 37501
rect 50200 37498 51000 37528
rect 49141 37496 51000 37498
rect 49141 37440 49146 37496
rect 49202 37440 51000 37496
rect 49141 37438 51000 37440
rect 49141 37435 49207 37438
rect 50200 37408 51000 37438
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 27946 37024 28262 37025
rect 27946 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28262 37024
rect 27946 36959 28262 36960
rect 37946 37024 38262 37025
rect 37946 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38262 37024
rect 37946 36959 38262 36960
rect 47946 37024 48262 37025
rect 47946 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48262 37024
rect 47946 36959 48262 36960
rect 49141 36682 49207 36685
rect 50200 36682 51000 36712
rect 49141 36680 51000 36682
rect 49141 36624 49146 36680
rect 49202 36624 51000 36680
rect 49141 36622 51000 36624
rect 49141 36619 49207 36622
rect 50200 36592 51000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 32946 36480 33262 36481
rect 32946 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33262 36480
rect 32946 36415 33262 36416
rect 42946 36480 43262 36481
rect 42946 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43262 36480
rect 42946 36415 43262 36416
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 27946 35936 28262 35937
rect 27946 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28262 35936
rect 27946 35871 28262 35872
rect 37946 35936 38262 35937
rect 37946 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38262 35936
rect 37946 35871 38262 35872
rect 47946 35936 48262 35937
rect 47946 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48262 35936
rect 47946 35871 48262 35872
rect 49325 35866 49391 35869
rect 50200 35866 51000 35896
rect 49325 35864 51000 35866
rect 49325 35808 49330 35864
rect 49386 35808 51000 35864
rect 49325 35806 51000 35808
rect 49325 35803 49391 35806
rect 50200 35776 51000 35806
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 32946 35392 33262 35393
rect 32946 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33262 35392
rect 32946 35327 33262 35328
rect 42946 35392 43262 35393
rect 42946 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43262 35392
rect 42946 35327 43262 35328
rect 49325 35050 49391 35053
rect 50200 35050 51000 35080
rect 49325 35048 51000 35050
rect 49325 34992 49330 35048
rect 49386 34992 51000 35048
rect 49325 34990 51000 34992
rect 49325 34987 49391 34990
rect 50200 34960 51000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 27946 34848 28262 34849
rect 27946 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28262 34848
rect 27946 34783 28262 34784
rect 37946 34848 38262 34849
rect 37946 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38262 34848
rect 37946 34783 38262 34784
rect 47946 34848 48262 34849
rect 47946 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48262 34848
rect 47946 34783 48262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 32946 34304 33262 34305
rect 32946 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33262 34304
rect 32946 34239 33262 34240
rect 42946 34304 43262 34305
rect 42946 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43262 34304
rect 42946 34239 43262 34240
rect 49325 34234 49391 34237
rect 50200 34234 51000 34264
rect 49325 34232 51000 34234
rect 49325 34176 49330 34232
rect 49386 34176 51000 34232
rect 49325 34174 51000 34176
rect 49325 34171 49391 34174
rect 50200 34144 51000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 27946 33760 28262 33761
rect 27946 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28262 33760
rect 27946 33695 28262 33696
rect 37946 33760 38262 33761
rect 37946 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38262 33760
rect 37946 33695 38262 33696
rect 47946 33760 48262 33761
rect 47946 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48262 33760
rect 47946 33695 48262 33696
rect 26182 33628 26188 33692
rect 26252 33690 26258 33692
rect 27521 33690 27587 33693
rect 26252 33688 27587 33690
rect 26252 33632 27526 33688
rect 27582 33632 27587 33688
rect 26252 33630 27587 33632
rect 26252 33628 26258 33630
rect 27521 33627 27587 33630
rect 40585 33418 40651 33421
rect 41229 33418 41295 33421
rect 31158 33416 41295 33418
rect 31158 33360 40590 33416
rect 40646 33360 41234 33416
rect 41290 33360 41295 33416
rect 31158 33358 41295 33360
rect 28574 33220 28580 33284
rect 28644 33282 28650 33284
rect 28901 33282 28967 33285
rect 31158 33282 31218 33358
rect 40585 33355 40651 33358
rect 41229 33355 41295 33358
rect 49325 33418 49391 33421
rect 50200 33418 51000 33448
rect 49325 33416 51000 33418
rect 49325 33360 49330 33416
rect 49386 33360 51000 33416
rect 49325 33358 51000 33360
rect 49325 33355 49391 33358
rect 50200 33328 51000 33358
rect 28644 33280 31218 33282
rect 28644 33224 28906 33280
rect 28962 33224 31218 33280
rect 28644 33222 31218 33224
rect 28644 33220 28650 33222
rect 28901 33219 28967 33222
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 32946 33216 33262 33217
rect 32946 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33262 33216
rect 32946 33151 33262 33152
rect 42946 33216 43262 33217
rect 42946 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43262 33216
rect 42946 33151 43262 33152
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 27946 32672 28262 32673
rect 27946 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28262 32672
rect 27946 32607 28262 32608
rect 37946 32672 38262 32673
rect 37946 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38262 32672
rect 37946 32607 38262 32608
rect 47946 32672 48262 32673
rect 47946 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48262 32672
rect 47946 32607 48262 32608
rect 49325 32602 49391 32605
rect 50200 32602 51000 32632
rect 49325 32600 51000 32602
rect 49325 32544 49330 32600
rect 49386 32544 51000 32600
rect 49325 32542 51000 32544
rect 49325 32539 49391 32542
rect 50200 32512 51000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 32946 32128 33262 32129
rect 32946 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33262 32128
rect 32946 32063 33262 32064
rect 42946 32128 43262 32129
rect 42946 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43262 32128
rect 42946 32063 43262 32064
rect 49325 31786 49391 31789
rect 50200 31786 51000 31816
rect 49325 31784 51000 31786
rect 49325 31728 49330 31784
rect 49386 31728 51000 31784
rect 49325 31726 51000 31728
rect 49325 31723 49391 31726
rect 50200 31696 51000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 27946 31584 28262 31585
rect 27946 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28262 31584
rect 27946 31519 28262 31520
rect 37946 31584 38262 31585
rect 37946 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38262 31584
rect 37946 31519 38262 31520
rect 47946 31584 48262 31585
rect 47946 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48262 31584
rect 47946 31519 48262 31520
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 32946 31040 33262 31041
rect 32946 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33262 31040
rect 32946 30975 33262 30976
rect 42946 31040 43262 31041
rect 42946 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43262 31040
rect 42946 30975 43262 30976
rect 49325 30970 49391 30973
rect 50200 30970 51000 31000
rect 49325 30968 51000 30970
rect 49325 30912 49330 30968
rect 49386 30912 51000 30968
rect 49325 30910 51000 30912
rect 49325 30907 49391 30910
rect 50200 30880 51000 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 27946 30496 28262 30497
rect 27946 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28262 30496
rect 27946 30431 28262 30432
rect 37946 30496 38262 30497
rect 37946 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38262 30496
rect 37946 30431 38262 30432
rect 47946 30496 48262 30497
rect 47946 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48262 30496
rect 47946 30431 48262 30432
rect 49325 30154 49391 30157
rect 50200 30154 51000 30184
rect 49325 30152 51000 30154
rect 49325 30096 49330 30152
rect 49386 30096 51000 30152
rect 49325 30094 51000 30096
rect 49325 30091 49391 30094
rect 50200 30064 51000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 32946 29952 33262 29953
rect 32946 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33262 29952
rect 32946 29887 33262 29888
rect 42946 29952 43262 29953
rect 42946 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43262 29952
rect 42946 29887 43262 29888
rect 35985 29610 36051 29613
rect 49969 29610 50035 29613
rect 35985 29608 50035 29610
rect 35985 29552 35990 29608
rect 36046 29552 49974 29608
rect 50030 29552 50035 29608
rect 35985 29550 50035 29552
rect 35985 29547 36051 29550
rect 49969 29547 50035 29550
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 27946 29408 28262 29409
rect 27946 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28262 29408
rect 27946 29343 28262 29344
rect 37946 29408 38262 29409
rect 37946 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38262 29408
rect 37946 29343 38262 29344
rect 47946 29408 48262 29409
rect 47946 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48262 29408
rect 47946 29343 48262 29344
rect 49325 29338 49391 29341
rect 50200 29338 51000 29368
rect 49325 29336 51000 29338
rect 49325 29280 49330 29336
rect 49386 29280 51000 29336
rect 49325 29278 51000 29280
rect 49325 29275 49391 29278
rect 50200 29248 51000 29278
rect 34513 29066 34579 29069
rect 35382 29066 35388 29068
rect 34513 29064 35388 29066
rect 34513 29008 34518 29064
rect 34574 29008 35388 29064
rect 34513 29006 35388 29008
rect 34513 29003 34579 29006
rect 35382 29004 35388 29006
rect 35452 29066 35458 29068
rect 35709 29066 35775 29069
rect 35452 29064 35775 29066
rect 35452 29008 35714 29064
rect 35770 29008 35775 29064
rect 35452 29006 35775 29008
rect 35452 29004 35458 29006
rect 35709 29003 35775 29006
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 32946 28864 33262 28865
rect 32946 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33262 28864
rect 32946 28799 33262 28800
rect 42946 28864 43262 28865
rect 42946 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43262 28864
rect 42946 28799 43262 28800
rect 49325 28522 49391 28525
rect 50200 28522 51000 28552
rect 49325 28520 51000 28522
rect 49325 28464 49330 28520
rect 49386 28464 51000 28520
rect 49325 28462 51000 28464
rect 49325 28459 49391 28462
rect 50200 28432 51000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 27946 28320 28262 28321
rect 27946 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28262 28320
rect 27946 28255 28262 28256
rect 37946 28320 38262 28321
rect 37946 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38262 28320
rect 37946 28255 38262 28256
rect 47946 28320 48262 28321
rect 47946 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48262 28320
rect 47946 28255 48262 28256
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 32946 27776 33262 27777
rect 32946 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33262 27776
rect 32946 27711 33262 27712
rect 42946 27776 43262 27777
rect 42946 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43262 27776
rect 42946 27711 43262 27712
rect 49325 27706 49391 27709
rect 50200 27706 51000 27736
rect 49325 27704 51000 27706
rect 49325 27648 49330 27704
rect 49386 27648 51000 27704
rect 49325 27646 51000 27648
rect 49325 27643 49391 27646
rect 50200 27616 51000 27646
rect 35985 27298 36051 27301
rect 36118 27298 36124 27300
rect 35985 27296 36124 27298
rect 35985 27240 35990 27296
rect 36046 27240 36124 27296
rect 35985 27238 36124 27240
rect 35985 27235 36051 27238
rect 36118 27236 36124 27238
rect 36188 27236 36194 27300
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 27946 27232 28262 27233
rect 27946 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28262 27232
rect 27946 27167 28262 27168
rect 37946 27232 38262 27233
rect 37946 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38262 27232
rect 37946 27167 38262 27168
rect 47946 27232 48262 27233
rect 47946 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48262 27232
rect 47946 27167 48262 27168
rect 49325 26890 49391 26893
rect 50200 26890 51000 26920
rect 49325 26888 51000 26890
rect 49325 26832 49330 26888
rect 49386 26832 51000 26888
rect 49325 26830 51000 26832
rect 49325 26827 49391 26830
rect 50200 26800 51000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 32946 26688 33262 26689
rect 32946 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33262 26688
rect 32946 26623 33262 26624
rect 42946 26688 43262 26689
rect 42946 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43262 26688
rect 42946 26623 43262 26624
rect 35249 26346 35315 26349
rect 35382 26346 35388 26348
rect 35249 26344 35388 26346
rect 35249 26288 35254 26344
rect 35310 26288 35388 26344
rect 35249 26286 35388 26288
rect 35249 26283 35315 26286
rect 35382 26284 35388 26286
rect 35452 26284 35458 26348
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 27946 26144 28262 26145
rect 27946 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28262 26144
rect 27946 26079 28262 26080
rect 37946 26144 38262 26145
rect 37946 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38262 26144
rect 37946 26079 38262 26080
rect 47946 26144 48262 26145
rect 47946 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48262 26144
rect 47946 26079 48262 26080
rect 48497 26074 48563 26077
rect 50200 26074 51000 26104
rect 48497 26072 51000 26074
rect 48497 26016 48502 26072
rect 48558 26016 51000 26072
rect 48497 26014 51000 26016
rect 48497 26011 48563 26014
rect 50200 25984 51000 26014
rect 33041 25802 33107 25805
rect 50429 25802 50495 25805
rect 33041 25800 50495 25802
rect 33041 25744 33046 25800
rect 33102 25744 50434 25800
rect 50490 25744 50495 25800
rect 33041 25742 50495 25744
rect 33041 25739 33107 25742
rect 50429 25739 50495 25742
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 32946 25600 33262 25601
rect 32946 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33262 25600
rect 32946 25535 33262 25536
rect 42946 25600 43262 25601
rect 42946 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43262 25600
rect 42946 25535 43262 25536
rect 49141 25258 49207 25261
rect 50200 25258 51000 25288
rect 49141 25256 51000 25258
rect 49141 25200 49146 25256
rect 49202 25200 51000 25256
rect 49141 25198 51000 25200
rect 49141 25195 49207 25198
rect 50200 25168 51000 25198
rect 42977 25122 43043 25125
rect 45553 25122 45619 25125
rect 42977 25120 45619 25122
rect 42977 25064 42982 25120
rect 43038 25064 45558 25120
rect 45614 25064 45619 25120
rect 42977 25062 45619 25064
rect 42977 25059 43043 25062
rect 45553 25059 45619 25062
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 27946 25056 28262 25057
rect 27946 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28262 25056
rect 27946 24991 28262 24992
rect 37946 25056 38262 25057
rect 37946 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38262 25056
rect 37946 24991 38262 24992
rect 47946 25056 48262 25057
rect 47946 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48262 25056
rect 47946 24991 48262 24992
rect 31845 24988 31911 24989
rect 31845 24984 31892 24988
rect 31956 24986 31962 24988
rect 31845 24928 31850 24984
rect 31845 24924 31892 24928
rect 31956 24926 32002 24986
rect 31956 24924 31962 24926
rect 31845 24923 31911 24924
rect 32581 24714 32647 24717
rect 35617 24714 35683 24717
rect 32581 24712 35683 24714
rect 32581 24656 32586 24712
rect 32642 24656 35622 24712
rect 35678 24656 35683 24712
rect 32581 24654 35683 24656
rect 32581 24651 32647 24654
rect 35617 24651 35683 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 49141 24442 49207 24445
rect 50200 24442 51000 24472
rect 49141 24440 51000 24442
rect 49141 24384 49146 24440
rect 49202 24384 51000 24440
rect 49141 24382 51000 24384
rect 49141 24379 49207 24382
rect 50200 24352 51000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 37590 23564 37596 23628
rect 37660 23626 37666 23628
rect 37825 23626 37891 23629
rect 37660 23624 37891 23626
rect 37660 23568 37830 23624
rect 37886 23568 37891 23624
rect 37660 23566 37891 23568
rect 37660 23564 37666 23566
rect 37825 23563 37891 23566
rect 49141 23626 49207 23629
rect 50200 23626 51000 23656
rect 49141 23624 51000 23626
rect 49141 23568 49146 23624
rect 49202 23568 51000 23624
rect 49141 23566 51000 23568
rect 49141 23563 49207 23566
rect 50200 23536 51000 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 49141 22810 49207 22813
rect 50200 22810 51000 22840
rect 49141 22808 51000 22810
rect 49141 22752 49146 22808
rect 49202 22752 51000 22808
rect 49141 22750 51000 22752
rect 49141 22747 49207 22750
rect 50200 22720 51000 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 49141 21994 49207 21997
rect 50200 21994 51000 22024
rect 49141 21992 51000 21994
rect 49141 21936 49146 21992
rect 49202 21936 51000 21992
rect 49141 21934 51000 21936
rect 49141 21931 49207 21934
rect 50200 21904 51000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 49141 21178 49207 21181
rect 50200 21178 51000 21208
rect 49141 21176 51000 21178
rect 49141 21120 49146 21176
rect 49202 21120 51000 21176
rect 49141 21118 51000 21120
rect 49141 21115 49207 21118
rect 50200 21088 51000 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 49141 20362 49207 20365
rect 50200 20362 51000 20392
rect 49141 20360 51000 20362
rect 49141 20304 49146 20360
rect 49202 20304 51000 20360
rect 49141 20302 51000 20304
rect 49141 20299 49207 20302
rect 50200 20272 51000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 40585 19546 40651 19549
rect 43897 19546 43963 19549
rect 40585 19544 43963 19546
rect 40585 19488 40590 19544
rect 40646 19488 43902 19544
rect 43958 19488 43963 19544
rect 40585 19486 43963 19488
rect 40585 19483 40651 19486
rect 43897 19483 43963 19486
rect 49141 19546 49207 19549
rect 50200 19546 51000 19576
rect 49141 19544 51000 19546
rect 49141 19488 49146 19544
rect 49202 19488 51000 19544
rect 49141 19486 51000 19488
rect 49141 19483 49207 19486
rect 50200 19456 51000 19486
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 49141 18730 49207 18733
rect 50200 18730 51000 18760
rect 49141 18728 51000 18730
rect 49141 18672 49146 18728
rect 49202 18672 51000 18728
rect 49141 18670 51000 18672
rect 49141 18667 49207 18670
rect 50200 18640 51000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 49141 17914 49207 17917
rect 50200 17914 51000 17944
rect 49141 17912 51000 17914
rect 49141 17856 49146 17912
rect 49202 17856 51000 17912
rect 49141 17854 51000 17856
rect 49141 17851 49207 17854
rect 50200 17824 51000 17854
rect 31886 17580 31892 17644
rect 31956 17642 31962 17644
rect 32029 17642 32095 17645
rect 31956 17640 32095 17642
rect 31956 17584 32034 17640
rect 32090 17584 32095 17640
rect 31956 17582 32095 17584
rect 31956 17580 31962 17582
rect 32029 17579 32095 17582
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 30925 17234 30991 17237
rect 33961 17234 34027 17237
rect 30925 17232 34027 17234
rect 30925 17176 30930 17232
rect 30986 17176 33966 17232
rect 34022 17176 34027 17232
rect 30925 17174 34027 17176
rect 30925 17171 30991 17174
rect 33961 17171 34027 17174
rect 49141 17098 49207 17101
rect 50200 17098 51000 17128
rect 49141 17096 51000 17098
rect 49141 17040 49146 17096
rect 49202 17040 51000 17096
rect 49141 17038 51000 17040
rect 49141 17035 49207 17038
rect 50200 17008 51000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 49141 16282 49207 16285
rect 50200 16282 51000 16312
rect 49141 16280 51000 16282
rect 49141 16224 49146 16280
rect 49202 16224 51000 16280
rect 49141 16222 51000 16224
rect 49141 16219 49207 16222
rect 50200 16192 51000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 49141 15466 49207 15469
rect 50200 15466 51000 15496
rect 49141 15464 51000 15466
rect 49141 15408 49146 15464
rect 49202 15408 51000 15464
rect 49141 15406 51000 15408
rect 49141 15403 49207 15406
rect 50200 15376 51000 15406
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 27654 14724 27660 14788
rect 27724 14786 27730 14788
rect 28257 14786 28323 14789
rect 27724 14784 28323 14786
rect 27724 14728 28262 14784
rect 28318 14728 28323 14784
rect 27724 14726 28323 14728
rect 27724 14724 27730 14726
rect 28257 14723 28323 14726
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 49141 14650 49207 14653
rect 50200 14650 51000 14680
rect 49141 14648 51000 14650
rect 49141 14592 49146 14648
rect 49202 14592 51000 14648
rect 49141 14590 51000 14592
rect 49141 14587 49207 14590
rect 50200 14560 51000 14590
rect 26969 14378 27035 14381
rect 36813 14378 36879 14381
rect 26969 14376 36879 14378
rect 26969 14320 26974 14376
rect 27030 14320 36818 14376
rect 36874 14320 36879 14376
rect 26969 14318 36879 14320
rect 26969 14315 27035 14318
rect 36813 14315 36879 14318
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 49141 13834 49207 13837
rect 50200 13834 51000 13864
rect 49141 13832 51000 13834
rect 49141 13776 49146 13832
rect 49202 13776 51000 13832
rect 49141 13774 51000 13776
rect 49141 13771 49207 13774
rect 50200 13744 51000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 49141 13018 49207 13021
rect 50200 13018 51000 13048
rect 49141 13016 51000 13018
rect 49141 12960 49146 13016
rect 49202 12960 51000 13016
rect 49141 12958 51000 12960
rect 49141 12955 49207 12958
rect 50200 12928 51000 12958
rect 29085 12882 29151 12885
rect 30465 12882 30531 12885
rect 29085 12880 30531 12882
rect 29085 12824 29090 12880
rect 29146 12824 30470 12880
rect 30526 12824 30531 12880
rect 29085 12822 30531 12824
rect 29085 12819 29151 12822
rect 30465 12819 30531 12822
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 27613 12474 27679 12477
rect 27797 12474 27863 12477
rect 27613 12472 27863 12474
rect 27613 12416 27618 12472
rect 27674 12416 27802 12472
rect 27858 12416 27863 12472
rect 27613 12414 27863 12416
rect 27613 12411 27679 12414
rect 27797 12411 27863 12414
rect 28165 12338 28231 12341
rect 31661 12338 31727 12341
rect 28165 12336 31727 12338
rect 28165 12280 28170 12336
rect 28226 12280 31666 12336
rect 31722 12280 31727 12336
rect 28165 12278 31727 12280
rect 28165 12275 28231 12278
rect 31661 12275 31727 12278
rect 38285 12202 38351 12205
rect 49141 12202 49207 12205
rect 50200 12202 51000 12232
rect 38285 12200 38394 12202
rect 38285 12144 38290 12200
rect 38346 12144 38394 12200
rect 38285 12139 38394 12144
rect 49141 12200 51000 12202
rect 49141 12144 49146 12200
rect 49202 12144 51000 12200
rect 49141 12142 51000 12144
rect 49141 12139 49207 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 28349 11794 28415 11797
rect 36261 11794 36327 11797
rect 28349 11792 36327 11794
rect 28349 11736 28354 11792
rect 28410 11736 36266 11792
rect 36322 11736 36327 11792
rect 28349 11734 36327 11736
rect 28349 11731 28415 11734
rect 36261 11731 36327 11734
rect 38334 11661 38394 12139
rect 50200 12112 51000 12142
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 38285 11656 38394 11661
rect 38285 11600 38290 11656
rect 38346 11600 38394 11656
rect 38285 11598 38394 11600
rect 38285 11595 38351 11598
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 49141 11386 49207 11389
rect 50200 11386 51000 11416
rect 49141 11384 51000 11386
rect 49141 11328 49146 11384
rect 49202 11328 51000 11384
rect 49141 11326 51000 11328
rect 49141 11323 49207 11326
rect 50200 11296 51000 11326
rect 29913 11250 29979 11253
rect 30557 11250 30623 11253
rect 29913 11248 30623 11250
rect 29913 11192 29918 11248
rect 29974 11192 30562 11248
rect 30618 11192 30623 11248
rect 29913 11190 30623 11192
rect 29913 11187 29979 11190
rect 30557 11187 30623 11190
rect 31385 11250 31451 11253
rect 38285 11250 38351 11253
rect 31385 11248 38351 11250
rect 31385 11192 31390 11248
rect 31446 11192 38290 11248
rect 38346 11192 38351 11248
rect 31385 11190 38351 11192
rect 31385 11187 31451 11190
rect 38285 11187 38351 11190
rect 32438 11052 32444 11116
rect 32508 11114 32514 11116
rect 32581 11114 32647 11117
rect 32508 11112 32647 11114
rect 32508 11056 32586 11112
rect 32642 11056 32647 11112
rect 32508 11054 32647 11056
rect 32508 11052 32514 11054
rect 32581 11051 32647 11054
rect 35341 11114 35407 11117
rect 36118 11114 36124 11116
rect 35341 11112 36124 11114
rect 35341 11056 35346 11112
rect 35402 11056 36124 11112
rect 35341 11054 36124 11056
rect 35341 11051 35407 11054
rect 36118 11052 36124 11054
rect 36188 11052 36194 11116
rect 29637 10978 29703 10981
rect 34237 10978 34303 10981
rect 29637 10976 34303 10978
rect 29637 10920 29642 10976
rect 29698 10920 34242 10976
rect 34298 10920 34303 10976
rect 29637 10918 34303 10920
rect 29637 10915 29703 10918
rect 34237 10915 34303 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 28625 10706 28691 10709
rect 30741 10706 30807 10709
rect 35382 10706 35388 10708
rect 28625 10704 35388 10706
rect 28625 10648 28630 10704
rect 28686 10648 30746 10704
rect 30802 10648 35388 10704
rect 28625 10646 35388 10648
rect 28625 10643 28691 10646
rect 30741 10643 30807 10646
rect 35382 10644 35388 10646
rect 35452 10706 35458 10708
rect 36077 10706 36143 10709
rect 35452 10704 36143 10706
rect 35452 10648 36082 10704
rect 36138 10648 36143 10704
rect 35452 10646 36143 10648
rect 35452 10644 35458 10646
rect 36077 10643 36143 10646
rect 49141 10570 49207 10573
rect 50200 10570 51000 10600
rect 49141 10568 51000 10570
rect 49141 10512 49146 10568
rect 49202 10512 51000 10568
rect 49141 10510 51000 10512
rect 49141 10507 49207 10510
rect 50200 10480 51000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 49141 9754 49207 9757
rect 50200 9754 51000 9784
rect 49141 9752 51000 9754
rect 49141 9696 49146 9752
rect 49202 9696 51000 9752
rect 49141 9694 51000 9696
rect 49141 9691 49207 9694
rect 50200 9664 51000 9694
rect 33225 9618 33291 9621
rect 35249 9618 35315 9621
rect 33225 9616 35315 9618
rect 33225 9560 33230 9616
rect 33286 9560 35254 9616
rect 35310 9560 35315 9616
rect 33225 9558 35315 9560
rect 33225 9555 33291 9558
rect 35249 9555 35315 9558
rect 30281 9482 30347 9485
rect 36537 9482 36603 9485
rect 30281 9480 36603 9482
rect 30281 9424 30286 9480
rect 30342 9424 36542 9480
rect 36598 9424 36603 9480
rect 30281 9422 36603 9424
rect 30281 9419 30347 9422
rect 36537 9419 36603 9422
rect 34789 9346 34855 9349
rect 37365 9346 37431 9349
rect 34789 9344 37431 9346
rect 34789 9288 34794 9344
rect 34850 9288 37370 9344
rect 37426 9288 37431 9344
rect 34789 9286 37431 9288
rect 34789 9283 34855 9286
rect 37365 9283 37431 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 32121 9074 32187 9077
rect 33501 9074 33567 9077
rect 32121 9072 33567 9074
rect 32121 9016 32126 9072
rect 32182 9016 33506 9072
rect 33562 9016 33567 9072
rect 32121 9014 33567 9016
rect 32121 9011 32187 9014
rect 33501 9011 33567 9014
rect 32581 8938 32647 8941
rect 40493 8938 40559 8941
rect 32581 8936 40559 8938
rect 32581 8880 32586 8936
rect 32642 8880 40498 8936
rect 40554 8880 40559 8936
rect 32581 8878 40559 8880
rect 32581 8875 32647 8878
rect 40493 8875 40559 8878
rect 49141 8938 49207 8941
rect 50200 8938 51000 8968
rect 49141 8936 51000 8938
rect 49141 8880 49146 8936
rect 49202 8880 51000 8936
rect 49141 8878 51000 8880
rect 49141 8875 49207 8878
rect 50200 8848 51000 8878
rect 0 8802 800 8832
rect 3417 8802 3483 8805
rect 0 8800 3483 8802
rect 0 8744 3422 8800
rect 3478 8744 3483 8800
rect 0 8742 3483 8744
rect 0 8712 800 8742
rect 3417 8739 3483 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 34421 8530 34487 8533
rect 40861 8530 40927 8533
rect 34421 8528 40927 8530
rect 34421 8472 34426 8528
rect 34482 8472 40866 8528
rect 40922 8472 40927 8528
rect 34421 8470 40927 8472
rect 34421 8467 34487 8470
rect 40861 8467 40927 8470
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 49141 8122 49207 8125
rect 50200 8122 51000 8152
rect 49141 8120 51000 8122
rect 49141 8064 49146 8120
rect 49202 8064 51000 8120
rect 49141 8062 51000 8064
rect 49141 8059 49207 8062
rect 50200 8032 51000 8062
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 49141 7306 49207 7309
rect 50200 7306 51000 7336
rect 49141 7304 51000 7306
rect 49141 7248 49146 7304
rect 49202 7248 51000 7304
rect 49141 7246 51000 7248
rect 49141 7243 49207 7246
rect 50200 7216 51000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 26182 6762 26188 6764
rect 6870 6702 26188 6762
rect 0 6490 800 6520
rect 6870 6490 6930 6702
rect 26182 6700 26188 6702
rect 26252 6700 26258 6764
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 0 6430 6930 6490
rect 49141 6490 49207 6493
rect 50200 6490 51000 6520
rect 49141 6488 51000 6490
rect 49141 6432 49146 6488
rect 49202 6432 51000 6488
rect 49141 6430 51000 6432
rect 0 6400 800 6430
rect 49141 6427 49207 6430
rect 50200 6400 51000 6430
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5674 49207 5677
rect 50200 5674 51000 5704
rect 49141 5672 51000 5674
rect 49141 5616 49146 5672
rect 49202 5616 51000 5672
rect 49141 5614 51000 5616
rect 49141 5611 49207 5614
rect 50200 5584 51000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 25313 5130 25379 5133
rect 37590 5130 37596 5132
rect 25313 5128 37596 5130
rect 25313 5072 25318 5128
rect 25374 5072 37596 5128
rect 25313 5070 37596 5072
rect 25313 5067 25379 5070
rect 37590 5068 37596 5070
rect 37660 5068 37666 5132
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 49141 4858 49207 4861
rect 50200 4858 51000 4888
rect 49141 4856 51000 4858
rect 49141 4800 49146 4856
rect 49202 4800 51000 4856
rect 49141 4798 51000 4800
rect 49141 4795 49207 4798
rect 50200 4768 51000 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 0 4178 800 4208
rect 28574 4178 28580 4180
rect 0 4118 28580 4178
rect 0 4088 800 4118
rect 28574 4116 28580 4118
rect 28644 4116 28650 4180
rect 49141 4042 49207 4045
rect 50200 4042 51000 4072
rect 49141 4040 51000 4042
rect 49141 3984 49146 4040
rect 49202 3984 51000 4040
rect 49141 3982 51000 3984
rect 49141 3979 49207 3982
rect 50200 3952 51000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 20253 3634 20319 3637
rect 32438 3634 32444 3636
rect 20253 3632 32444 3634
rect 20253 3576 20258 3632
rect 20314 3576 32444 3632
rect 20253 3574 32444 3576
rect 20253 3571 20319 3574
rect 32438 3572 32444 3574
rect 32508 3572 32514 3636
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 49141 3226 49207 3229
rect 50200 3226 51000 3256
rect 49141 3224 51000 3226
rect 49141 3168 49146 3224
rect 49202 3168 51000 3224
rect 49141 3166 51000 3168
rect 49141 3163 49207 3166
rect 50200 3136 51000 3166
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 9857 2410 9923 2413
rect 27654 2410 27660 2412
rect 9857 2408 27660 2410
rect 9857 2352 9862 2408
rect 9918 2352 27660 2408
rect 9857 2350 27660 2352
rect 9857 2347 9923 2350
rect 27654 2348 27660 2350
rect 27724 2348 27730 2412
rect 47853 2410 47919 2413
rect 50200 2410 51000 2440
rect 47853 2408 51000 2410
rect 47853 2352 47858 2408
rect 47914 2352 51000 2408
rect 47853 2350 51000 2352
rect 47853 2347 47919 2350
rect 50200 2320 51000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 1866 800 1896
rect 3417 1866 3483 1869
rect 0 1864 3483 1866
rect 0 1808 3422 1864
rect 3478 1808 3483 1864
rect 0 1806 3483 1808
rect 0 1776 800 1806
rect 3417 1803 3483 1806
rect 49233 1594 49299 1597
rect 50200 1594 51000 1624
rect 49233 1592 51000 1594
rect 49233 1536 49238 1592
rect 49294 1536 51000 1592
rect 49233 1534 51000 1536
rect 49233 1531 49299 1534
rect 50200 1504 51000 1534
rect 48681 778 48747 781
rect 50200 778 51000 808
rect 48681 776 51000 778
rect 48681 720 48686 776
rect 48742 720 51000 776
rect 48681 718 51000 720
rect 48681 715 48747 718
rect 50200 688 51000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 27952 54428 28016 54432
rect 27952 54372 27956 54428
rect 27956 54372 28012 54428
rect 28012 54372 28016 54428
rect 27952 54368 28016 54372
rect 28032 54428 28096 54432
rect 28032 54372 28036 54428
rect 28036 54372 28092 54428
rect 28092 54372 28096 54428
rect 28032 54368 28096 54372
rect 28112 54428 28176 54432
rect 28112 54372 28116 54428
rect 28116 54372 28172 54428
rect 28172 54372 28176 54428
rect 28112 54368 28176 54372
rect 28192 54428 28256 54432
rect 28192 54372 28196 54428
rect 28196 54372 28252 54428
rect 28252 54372 28256 54428
rect 28192 54368 28256 54372
rect 37952 54428 38016 54432
rect 37952 54372 37956 54428
rect 37956 54372 38012 54428
rect 38012 54372 38016 54428
rect 37952 54368 38016 54372
rect 38032 54428 38096 54432
rect 38032 54372 38036 54428
rect 38036 54372 38092 54428
rect 38092 54372 38096 54428
rect 38032 54368 38096 54372
rect 38112 54428 38176 54432
rect 38112 54372 38116 54428
rect 38116 54372 38172 54428
rect 38172 54372 38176 54428
rect 38112 54368 38176 54372
rect 38192 54428 38256 54432
rect 38192 54372 38196 54428
rect 38196 54372 38252 54428
rect 38252 54372 38256 54428
rect 38192 54368 38256 54372
rect 47952 54428 48016 54432
rect 47952 54372 47956 54428
rect 47956 54372 48012 54428
rect 48012 54372 48016 54428
rect 47952 54368 48016 54372
rect 48032 54428 48096 54432
rect 48032 54372 48036 54428
rect 48036 54372 48092 54428
rect 48092 54372 48096 54428
rect 48032 54368 48096 54372
rect 48112 54428 48176 54432
rect 48112 54372 48116 54428
rect 48116 54372 48172 54428
rect 48172 54372 48176 54428
rect 48112 54368 48176 54372
rect 48192 54428 48256 54432
rect 48192 54372 48196 54428
rect 48196 54372 48252 54428
rect 48252 54372 48256 54428
rect 48192 54368 48256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 32952 53884 33016 53888
rect 32952 53828 32956 53884
rect 32956 53828 33012 53884
rect 33012 53828 33016 53884
rect 32952 53824 33016 53828
rect 33032 53884 33096 53888
rect 33032 53828 33036 53884
rect 33036 53828 33092 53884
rect 33092 53828 33096 53884
rect 33032 53824 33096 53828
rect 33112 53884 33176 53888
rect 33112 53828 33116 53884
rect 33116 53828 33172 53884
rect 33172 53828 33176 53884
rect 33112 53824 33176 53828
rect 33192 53884 33256 53888
rect 33192 53828 33196 53884
rect 33196 53828 33252 53884
rect 33252 53828 33256 53884
rect 33192 53824 33256 53828
rect 42952 53884 43016 53888
rect 42952 53828 42956 53884
rect 42956 53828 43012 53884
rect 43012 53828 43016 53884
rect 42952 53824 43016 53828
rect 43032 53884 43096 53888
rect 43032 53828 43036 53884
rect 43036 53828 43092 53884
rect 43092 53828 43096 53884
rect 43032 53824 43096 53828
rect 43112 53884 43176 53888
rect 43112 53828 43116 53884
rect 43116 53828 43172 53884
rect 43172 53828 43176 53884
rect 43112 53824 43176 53828
rect 43192 53884 43256 53888
rect 43192 53828 43196 53884
rect 43196 53828 43252 53884
rect 43252 53828 43256 53884
rect 43192 53824 43256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 27952 53340 28016 53344
rect 27952 53284 27956 53340
rect 27956 53284 28012 53340
rect 28012 53284 28016 53340
rect 27952 53280 28016 53284
rect 28032 53340 28096 53344
rect 28032 53284 28036 53340
rect 28036 53284 28092 53340
rect 28092 53284 28096 53340
rect 28032 53280 28096 53284
rect 28112 53340 28176 53344
rect 28112 53284 28116 53340
rect 28116 53284 28172 53340
rect 28172 53284 28176 53340
rect 28112 53280 28176 53284
rect 28192 53340 28256 53344
rect 28192 53284 28196 53340
rect 28196 53284 28252 53340
rect 28252 53284 28256 53340
rect 28192 53280 28256 53284
rect 37952 53340 38016 53344
rect 37952 53284 37956 53340
rect 37956 53284 38012 53340
rect 38012 53284 38016 53340
rect 37952 53280 38016 53284
rect 38032 53340 38096 53344
rect 38032 53284 38036 53340
rect 38036 53284 38092 53340
rect 38092 53284 38096 53340
rect 38032 53280 38096 53284
rect 38112 53340 38176 53344
rect 38112 53284 38116 53340
rect 38116 53284 38172 53340
rect 38172 53284 38176 53340
rect 38112 53280 38176 53284
rect 38192 53340 38256 53344
rect 38192 53284 38196 53340
rect 38196 53284 38252 53340
rect 38252 53284 38256 53340
rect 38192 53280 38256 53284
rect 47952 53340 48016 53344
rect 47952 53284 47956 53340
rect 47956 53284 48012 53340
rect 48012 53284 48016 53340
rect 47952 53280 48016 53284
rect 48032 53340 48096 53344
rect 48032 53284 48036 53340
rect 48036 53284 48092 53340
rect 48092 53284 48096 53340
rect 48032 53280 48096 53284
rect 48112 53340 48176 53344
rect 48112 53284 48116 53340
rect 48116 53284 48172 53340
rect 48172 53284 48176 53340
rect 48112 53280 48176 53284
rect 48192 53340 48256 53344
rect 48192 53284 48196 53340
rect 48196 53284 48252 53340
rect 48252 53284 48256 53340
rect 48192 53280 48256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 32952 52796 33016 52800
rect 32952 52740 32956 52796
rect 32956 52740 33012 52796
rect 33012 52740 33016 52796
rect 32952 52736 33016 52740
rect 33032 52796 33096 52800
rect 33032 52740 33036 52796
rect 33036 52740 33092 52796
rect 33092 52740 33096 52796
rect 33032 52736 33096 52740
rect 33112 52796 33176 52800
rect 33112 52740 33116 52796
rect 33116 52740 33172 52796
rect 33172 52740 33176 52796
rect 33112 52736 33176 52740
rect 33192 52796 33256 52800
rect 33192 52740 33196 52796
rect 33196 52740 33252 52796
rect 33252 52740 33256 52796
rect 33192 52736 33256 52740
rect 42952 52796 43016 52800
rect 42952 52740 42956 52796
rect 42956 52740 43012 52796
rect 43012 52740 43016 52796
rect 42952 52736 43016 52740
rect 43032 52796 43096 52800
rect 43032 52740 43036 52796
rect 43036 52740 43092 52796
rect 43092 52740 43096 52796
rect 43032 52736 43096 52740
rect 43112 52796 43176 52800
rect 43112 52740 43116 52796
rect 43116 52740 43172 52796
rect 43172 52740 43176 52796
rect 43112 52736 43176 52740
rect 43192 52796 43256 52800
rect 43192 52740 43196 52796
rect 43196 52740 43252 52796
rect 43252 52740 43256 52796
rect 43192 52736 43256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 27952 52252 28016 52256
rect 27952 52196 27956 52252
rect 27956 52196 28012 52252
rect 28012 52196 28016 52252
rect 27952 52192 28016 52196
rect 28032 52252 28096 52256
rect 28032 52196 28036 52252
rect 28036 52196 28092 52252
rect 28092 52196 28096 52252
rect 28032 52192 28096 52196
rect 28112 52252 28176 52256
rect 28112 52196 28116 52252
rect 28116 52196 28172 52252
rect 28172 52196 28176 52252
rect 28112 52192 28176 52196
rect 28192 52252 28256 52256
rect 28192 52196 28196 52252
rect 28196 52196 28252 52252
rect 28252 52196 28256 52252
rect 28192 52192 28256 52196
rect 37952 52252 38016 52256
rect 37952 52196 37956 52252
rect 37956 52196 38012 52252
rect 38012 52196 38016 52252
rect 37952 52192 38016 52196
rect 38032 52252 38096 52256
rect 38032 52196 38036 52252
rect 38036 52196 38092 52252
rect 38092 52196 38096 52252
rect 38032 52192 38096 52196
rect 38112 52252 38176 52256
rect 38112 52196 38116 52252
rect 38116 52196 38172 52252
rect 38172 52196 38176 52252
rect 38112 52192 38176 52196
rect 38192 52252 38256 52256
rect 38192 52196 38196 52252
rect 38196 52196 38252 52252
rect 38252 52196 38256 52252
rect 38192 52192 38256 52196
rect 47952 52252 48016 52256
rect 47952 52196 47956 52252
rect 47956 52196 48012 52252
rect 48012 52196 48016 52252
rect 47952 52192 48016 52196
rect 48032 52252 48096 52256
rect 48032 52196 48036 52252
rect 48036 52196 48092 52252
rect 48092 52196 48096 52252
rect 48032 52192 48096 52196
rect 48112 52252 48176 52256
rect 48112 52196 48116 52252
rect 48116 52196 48172 52252
rect 48172 52196 48176 52252
rect 48112 52192 48176 52196
rect 48192 52252 48256 52256
rect 48192 52196 48196 52252
rect 48196 52196 48252 52252
rect 48252 52196 48256 52252
rect 48192 52192 48256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 32952 51708 33016 51712
rect 32952 51652 32956 51708
rect 32956 51652 33012 51708
rect 33012 51652 33016 51708
rect 32952 51648 33016 51652
rect 33032 51708 33096 51712
rect 33032 51652 33036 51708
rect 33036 51652 33092 51708
rect 33092 51652 33096 51708
rect 33032 51648 33096 51652
rect 33112 51708 33176 51712
rect 33112 51652 33116 51708
rect 33116 51652 33172 51708
rect 33172 51652 33176 51708
rect 33112 51648 33176 51652
rect 33192 51708 33256 51712
rect 33192 51652 33196 51708
rect 33196 51652 33252 51708
rect 33252 51652 33256 51708
rect 33192 51648 33256 51652
rect 42952 51708 43016 51712
rect 42952 51652 42956 51708
rect 42956 51652 43012 51708
rect 43012 51652 43016 51708
rect 42952 51648 43016 51652
rect 43032 51708 43096 51712
rect 43032 51652 43036 51708
rect 43036 51652 43092 51708
rect 43092 51652 43096 51708
rect 43032 51648 43096 51652
rect 43112 51708 43176 51712
rect 43112 51652 43116 51708
rect 43116 51652 43172 51708
rect 43172 51652 43176 51708
rect 43112 51648 43176 51652
rect 43192 51708 43256 51712
rect 43192 51652 43196 51708
rect 43196 51652 43252 51708
rect 43252 51652 43256 51708
rect 43192 51648 43256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 27952 51164 28016 51168
rect 27952 51108 27956 51164
rect 27956 51108 28012 51164
rect 28012 51108 28016 51164
rect 27952 51104 28016 51108
rect 28032 51164 28096 51168
rect 28032 51108 28036 51164
rect 28036 51108 28092 51164
rect 28092 51108 28096 51164
rect 28032 51104 28096 51108
rect 28112 51164 28176 51168
rect 28112 51108 28116 51164
rect 28116 51108 28172 51164
rect 28172 51108 28176 51164
rect 28112 51104 28176 51108
rect 28192 51164 28256 51168
rect 28192 51108 28196 51164
rect 28196 51108 28252 51164
rect 28252 51108 28256 51164
rect 28192 51104 28256 51108
rect 37952 51164 38016 51168
rect 37952 51108 37956 51164
rect 37956 51108 38012 51164
rect 38012 51108 38016 51164
rect 37952 51104 38016 51108
rect 38032 51164 38096 51168
rect 38032 51108 38036 51164
rect 38036 51108 38092 51164
rect 38092 51108 38096 51164
rect 38032 51104 38096 51108
rect 38112 51164 38176 51168
rect 38112 51108 38116 51164
rect 38116 51108 38172 51164
rect 38172 51108 38176 51164
rect 38112 51104 38176 51108
rect 38192 51164 38256 51168
rect 38192 51108 38196 51164
rect 38196 51108 38252 51164
rect 38252 51108 38256 51164
rect 38192 51104 38256 51108
rect 47952 51164 48016 51168
rect 47952 51108 47956 51164
rect 47956 51108 48012 51164
rect 48012 51108 48016 51164
rect 47952 51104 48016 51108
rect 48032 51164 48096 51168
rect 48032 51108 48036 51164
rect 48036 51108 48092 51164
rect 48092 51108 48096 51164
rect 48032 51104 48096 51108
rect 48112 51164 48176 51168
rect 48112 51108 48116 51164
rect 48116 51108 48172 51164
rect 48172 51108 48176 51164
rect 48112 51104 48176 51108
rect 48192 51164 48256 51168
rect 48192 51108 48196 51164
rect 48196 51108 48252 51164
rect 48252 51108 48256 51164
rect 48192 51104 48256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 32952 50620 33016 50624
rect 32952 50564 32956 50620
rect 32956 50564 33012 50620
rect 33012 50564 33016 50620
rect 32952 50560 33016 50564
rect 33032 50620 33096 50624
rect 33032 50564 33036 50620
rect 33036 50564 33092 50620
rect 33092 50564 33096 50620
rect 33032 50560 33096 50564
rect 33112 50620 33176 50624
rect 33112 50564 33116 50620
rect 33116 50564 33172 50620
rect 33172 50564 33176 50620
rect 33112 50560 33176 50564
rect 33192 50620 33256 50624
rect 33192 50564 33196 50620
rect 33196 50564 33252 50620
rect 33252 50564 33256 50620
rect 33192 50560 33256 50564
rect 42952 50620 43016 50624
rect 42952 50564 42956 50620
rect 42956 50564 43012 50620
rect 43012 50564 43016 50620
rect 42952 50560 43016 50564
rect 43032 50620 43096 50624
rect 43032 50564 43036 50620
rect 43036 50564 43092 50620
rect 43092 50564 43096 50620
rect 43032 50560 43096 50564
rect 43112 50620 43176 50624
rect 43112 50564 43116 50620
rect 43116 50564 43172 50620
rect 43172 50564 43176 50620
rect 43112 50560 43176 50564
rect 43192 50620 43256 50624
rect 43192 50564 43196 50620
rect 43196 50564 43252 50620
rect 43252 50564 43256 50620
rect 43192 50560 43256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 27952 50076 28016 50080
rect 27952 50020 27956 50076
rect 27956 50020 28012 50076
rect 28012 50020 28016 50076
rect 27952 50016 28016 50020
rect 28032 50076 28096 50080
rect 28032 50020 28036 50076
rect 28036 50020 28092 50076
rect 28092 50020 28096 50076
rect 28032 50016 28096 50020
rect 28112 50076 28176 50080
rect 28112 50020 28116 50076
rect 28116 50020 28172 50076
rect 28172 50020 28176 50076
rect 28112 50016 28176 50020
rect 28192 50076 28256 50080
rect 28192 50020 28196 50076
rect 28196 50020 28252 50076
rect 28252 50020 28256 50076
rect 28192 50016 28256 50020
rect 37952 50076 38016 50080
rect 37952 50020 37956 50076
rect 37956 50020 38012 50076
rect 38012 50020 38016 50076
rect 37952 50016 38016 50020
rect 38032 50076 38096 50080
rect 38032 50020 38036 50076
rect 38036 50020 38092 50076
rect 38092 50020 38096 50076
rect 38032 50016 38096 50020
rect 38112 50076 38176 50080
rect 38112 50020 38116 50076
rect 38116 50020 38172 50076
rect 38172 50020 38176 50076
rect 38112 50016 38176 50020
rect 38192 50076 38256 50080
rect 38192 50020 38196 50076
rect 38196 50020 38252 50076
rect 38252 50020 38256 50076
rect 38192 50016 38256 50020
rect 47952 50076 48016 50080
rect 47952 50020 47956 50076
rect 47956 50020 48012 50076
rect 48012 50020 48016 50076
rect 47952 50016 48016 50020
rect 48032 50076 48096 50080
rect 48032 50020 48036 50076
rect 48036 50020 48092 50076
rect 48092 50020 48096 50076
rect 48032 50016 48096 50020
rect 48112 50076 48176 50080
rect 48112 50020 48116 50076
rect 48116 50020 48172 50076
rect 48172 50020 48176 50076
rect 48112 50016 48176 50020
rect 48192 50076 48256 50080
rect 48192 50020 48196 50076
rect 48196 50020 48252 50076
rect 48252 50020 48256 50076
rect 48192 50016 48256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 32952 49532 33016 49536
rect 32952 49476 32956 49532
rect 32956 49476 33012 49532
rect 33012 49476 33016 49532
rect 32952 49472 33016 49476
rect 33032 49532 33096 49536
rect 33032 49476 33036 49532
rect 33036 49476 33092 49532
rect 33092 49476 33096 49532
rect 33032 49472 33096 49476
rect 33112 49532 33176 49536
rect 33112 49476 33116 49532
rect 33116 49476 33172 49532
rect 33172 49476 33176 49532
rect 33112 49472 33176 49476
rect 33192 49532 33256 49536
rect 33192 49476 33196 49532
rect 33196 49476 33252 49532
rect 33252 49476 33256 49532
rect 33192 49472 33256 49476
rect 42952 49532 43016 49536
rect 42952 49476 42956 49532
rect 42956 49476 43012 49532
rect 43012 49476 43016 49532
rect 42952 49472 43016 49476
rect 43032 49532 43096 49536
rect 43032 49476 43036 49532
rect 43036 49476 43092 49532
rect 43092 49476 43096 49532
rect 43032 49472 43096 49476
rect 43112 49532 43176 49536
rect 43112 49476 43116 49532
rect 43116 49476 43172 49532
rect 43172 49476 43176 49532
rect 43112 49472 43176 49476
rect 43192 49532 43256 49536
rect 43192 49476 43196 49532
rect 43196 49476 43252 49532
rect 43252 49476 43256 49532
rect 43192 49472 43256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 27952 48988 28016 48992
rect 27952 48932 27956 48988
rect 27956 48932 28012 48988
rect 28012 48932 28016 48988
rect 27952 48928 28016 48932
rect 28032 48988 28096 48992
rect 28032 48932 28036 48988
rect 28036 48932 28092 48988
rect 28092 48932 28096 48988
rect 28032 48928 28096 48932
rect 28112 48988 28176 48992
rect 28112 48932 28116 48988
rect 28116 48932 28172 48988
rect 28172 48932 28176 48988
rect 28112 48928 28176 48932
rect 28192 48988 28256 48992
rect 28192 48932 28196 48988
rect 28196 48932 28252 48988
rect 28252 48932 28256 48988
rect 28192 48928 28256 48932
rect 37952 48988 38016 48992
rect 37952 48932 37956 48988
rect 37956 48932 38012 48988
rect 38012 48932 38016 48988
rect 37952 48928 38016 48932
rect 38032 48988 38096 48992
rect 38032 48932 38036 48988
rect 38036 48932 38092 48988
rect 38092 48932 38096 48988
rect 38032 48928 38096 48932
rect 38112 48988 38176 48992
rect 38112 48932 38116 48988
rect 38116 48932 38172 48988
rect 38172 48932 38176 48988
rect 38112 48928 38176 48932
rect 38192 48988 38256 48992
rect 38192 48932 38196 48988
rect 38196 48932 38252 48988
rect 38252 48932 38256 48988
rect 38192 48928 38256 48932
rect 47952 48988 48016 48992
rect 47952 48932 47956 48988
rect 47956 48932 48012 48988
rect 48012 48932 48016 48988
rect 47952 48928 48016 48932
rect 48032 48988 48096 48992
rect 48032 48932 48036 48988
rect 48036 48932 48092 48988
rect 48092 48932 48096 48988
rect 48032 48928 48096 48932
rect 48112 48988 48176 48992
rect 48112 48932 48116 48988
rect 48116 48932 48172 48988
rect 48172 48932 48176 48988
rect 48112 48928 48176 48932
rect 48192 48988 48256 48992
rect 48192 48932 48196 48988
rect 48196 48932 48252 48988
rect 48252 48932 48256 48988
rect 48192 48928 48256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 32952 48444 33016 48448
rect 32952 48388 32956 48444
rect 32956 48388 33012 48444
rect 33012 48388 33016 48444
rect 32952 48384 33016 48388
rect 33032 48444 33096 48448
rect 33032 48388 33036 48444
rect 33036 48388 33092 48444
rect 33092 48388 33096 48444
rect 33032 48384 33096 48388
rect 33112 48444 33176 48448
rect 33112 48388 33116 48444
rect 33116 48388 33172 48444
rect 33172 48388 33176 48444
rect 33112 48384 33176 48388
rect 33192 48444 33256 48448
rect 33192 48388 33196 48444
rect 33196 48388 33252 48444
rect 33252 48388 33256 48444
rect 33192 48384 33256 48388
rect 42952 48444 43016 48448
rect 42952 48388 42956 48444
rect 42956 48388 43012 48444
rect 43012 48388 43016 48444
rect 42952 48384 43016 48388
rect 43032 48444 43096 48448
rect 43032 48388 43036 48444
rect 43036 48388 43092 48444
rect 43092 48388 43096 48444
rect 43032 48384 43096 48388
rect 43112 48444 43176 48448
rect 43112 48388 43116 48444
rect 43116 48388 43172 48444
rect 43172 48388 43176 48444
rect 43112 48384 43176 48388
rect 43192 48444 43256 48448
rect 43192 48388 43196 48444
rect 43196 48388 43252 48444
rect 43252 48388 43256 48444
rect 43192 48384 43256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 27952 47900 28016 47904
rect 27952 47844 27956 47900
rect 27956 47844 28012 47900
rect 28012 47844 28016 47900
rect 27952 47840 28016 47844
rect 28032 47900 28096 47904
rect 28032 47844 28036 47900
rect 28036 47844 28092 47900
rect 28092 47844 28096 47900
rect 28032 47840 28096 47844
rect 28112 47900 28176 47904
rect 28112 47844 28116 47900
rect 28116 47844 28172 47900
rect 28172 47844 28176 47900
rect 28112 47840 28176 47844
rect 28192 47900 28256 47904
rect 28192 47844 28196 47900
rect 28196 47844 28252 47900
rect 28252 47844 28256 47900
rect 28192 47840 28256 47844
rect 37952 47900 38016 47904
rect 37952 47844 37956 47900
rect 37956 47844 38012 47900
rect 38012 47844 38016 47900
rect 37952 47840 38016 47844
rect 38032 47900 38096 47904
rect 38032 47844 38036 47900
rect 38036 47844 38092 47900
rect 38092 47844 38096 47900
rect 38032 47840 38096 47844
rect 38112 47900 38176 47904
rect 38112 47844 38116 47900
rect 38116 47844 38172 47900
rect 38172 47844 38176 47900
rect 38112 47840 38176 47844
rect 38192 47900 38256 47904
rect 38192 47844 38196 47900
rect 38196 47844 38252 47900
rect 38252 47844 38256 47900
rect 38192 47840 38256 47844
rect 47952 47900 48016 47904
rect 47952 47844 47956 47900
rect 47956 47844 48012 47900
rect 48012 47844 48016 47900
rect 47952 47840 48016 47844
rect 48032 47900 48096 47904
rect 48032 47844 48036 47900
rect 48036 47844 48092 47900
rect 48092 47844 48096 47900
rect 48032 47840 48096 47844
rect 48112 47900 48176 47904
rect 48112 47844 48116 47900
rect 48116 47844 48172 47900
rect 48172 47844 48176 47900
rect 48112 47840 48176 47844
rect 48192 47900 48256 47904
rect 48192 47844 48196 47900
rect 48196 47844 48252 47900
rect 48252 47844 48256 47900
rect 48192 47840 48256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 32952 47356 33016 47360
rect 32952 47300 32956 47356
rect 32956 47300 33012 47356
rect 33012 47300 33016 47356
rect 32952 47296 33016 47300
rect 33032 47356 33096 47360
rect 33032 47300 33036 47356
rect 33036 47300 33092 47356
rect 33092 47300 33096 47356
rect 33032 47296 33096 47300
rect 33112 47356 33176 47360
rect 33112 47300 33116 47356
rect 33116 47300 33172 47356
rect 33172 47300 33176 47356
rect 33112 47296 33176 47300
rect 33192 47356 33256 47360
rect 33192 47300 33196 47356
rect 33196 47300 33252 47356
rect 33252 47300 33256 47356
rect 33192 47296 33256 47300
rect 42952 47356 43016 47360
rect 42952 47300 42956 47356
rect 42956 47300 43012 47356
rect 43012 47300 43016 47356
rect 42952 47296 43016 47300
rect 43032 47356 43096 47360
rect 43032 47300 43036 47356
rect 43036 47300 43092 47356
rect 43092 47300 43096 47356
rect 43032 47296 43096 47300
rect 43112 47356 43176 47360
rect 43112 47300 43116 47356
rect 43116 47300 43172 47356
rect 43172 47300 43176 47356
rect 43112 47296 43176 47300
rect 43192 47356 43256 47360
rect 43192 47300 43196 47356
rect 43196 47300 43252 47356
rect 43252 47300 43256 47356
rect 43192 47296 43256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 27952 46812 28016 46816
rect 27952 46756 27956 46812
rect 27956 46756 28012 46812
rect 28012 46756 28016 46812
rect 27952 46752 28016 46756
rect 28032 46812 28096 46816
rect 28032 46756 28036 46812
rect 28036 46756 28092 46812
rect 28092 46756 28096 46812
rect 28032 46752 28096 46756
rect 28112 46812 28176 46816
rect 28112 46756 28116 46812
rect 28116 46756 28172 46812
rect 28172 46756 28176 46812
rect 28112 46752 28176 46756
rect 28192 46812 28256 46816
rect 28192 46756 28196 46812
rect 28196 46756 28252 46812
rect 28252 46756 28256 46812
rect 28192 46752 28256 46756
rect 37952 46812 38016 46816
rect 37952 46756 37956 46812
rect 37956 46756 38012 46812
rect 38012 46756 38016 46812
rect 37952 46752 38016 46756
rect 38032 46812 38096 46816
rect 38032 46756 38036 46812
rect 38036 46756 38092 46812
rect 38092 46756 38096 46812
rect 38032 46752 38096 46756
rect 38112 46812 38176 46816
rect 38112 46756 38116 46812
rect 38116 46756 38172 46812
rect 38172 46756 38176 46812
rect 38112 46752 38176 46756
rect 38192 46812 38256 46816
rect 38192 46756 38196 46812
rect 38196 46756 38252 46812
rect 38252 46756 38256 46812
rect 38192 46752 38256 46756
rect 47952 46812 48016 46816
rect 47952 46756 47956 46812
rect 47956 46756 48012 46812
rect 48012 46756 48016 46812
rect 47952 46752 48016 46756
rect 48032 46812 48096 46816
rect 48032 46756 48036 46812
rect 48036 46756 48092 46812
rect 48092 46756 48096 46812
rect 48032 46752 48096 46756
rect 48112 46812 48176 46816
rect 48112 46756 48116 46812
rect 48116 46756 48172 46812
rect 48172 46756 48176 46812
rect 48112 46752 48176 46756
rect 48192 46812 48256 46816
rect 48192 46756 48196 46812
rect 48196 46756 48252 46812
rect 48252 46756 48256 46812
rect 48192 46752 48256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 32952 46268 33016 46272
rect 32952 46212 32956 46268
rect 32956 46212 33012 46268
rect 33012 46212 33016 46268
rect 32952 46208 33016 46212
rect 33032 46268 33096 46272
rect 33032 46212 33036 46268
rect 33036 46212 33092 46268
rect 33092 46212 33096 46268
rect 33032 46208 33096 46212
rect 33112 46268 33176 46272
rect 33112 46212 33116 46268
rect 33116 46212 33172 46268
rect 33172 46212 33176 46268
rect 33112 46208 33176 46212
rect 33192 46268 33256 46272
rect 33192 46212 33196 46268
rect 33196 46212 33252 46268
rect 33252 46212 33256 46268
rect 33192 46208 33256 46212
rect 42952 46268 43016 46272
rect 42952 46212 42956 46268
rect 42956 46212 43012 46268
rect 43012 46212 43016 46268
rect 42952 46208 43016 46212
rect 43032 46268 43096 46272
rect 43032 46212 43036 46268
rect 43036 46212 43092 46268
rect 43092 46212 43096 46268
rect 43032 46208 43096 46212
rect 43112 46268 43176 46272
rect 43112 46212 43116 46268
rect 43116 46212 43172 46268
rect 43172 46212 43176 46268
rect 43112 46208 43176 46212
rect 43192 46268 43256 46272
rect 43192 46212 43196 46268
rect 43196 46212 43252 46268
rect 43252 46212 43256 46268
rect 43192 46208 43256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 27952 45724 28016 45728
rect 27952 45668 27956 45724
rect 27956 45668 28012 45724
rect 28012 45668 28016 45724
rect 27952 45664 28016 45668
rect 28032 45724 28096 45728
rect 28032 45668 28036 45724
rect 28036 45668 28092 45724
rect 28092 45668 28096 45724
rect 28032 45664 28096 45668
rect 28112 45724 28176 45728
rect 28112 45668 28116 45724
rect 28116 45668 28172 45724
rect 28172 45668 28176 45724
rect 28112 45664 28176 45668
rect 28192 45724 28256 45728
rect 28192 45668 28196 45724
rect 28196 45668 28252 45724
rect 28252 45668 28256 45724
rect 28192 45664 28256 45668
rect 37952 45724 38016 45728
rect 37952 45668 37956 45724
rect 37956 45668 38012 45724
rect 38012 45668 38016 45724
rect 37952 45664 38016 45668
rect 38032 45724 38096 45728
rect 38032 45668 38036 45724
rect 38036 45668 38092 45724
rect 38092 45668 38096 45724
rect 38032 45664 38096 45668
rect 38112 45724 38176 45728
rect 38112 45668 38116 45724
rect 38116 45668 38172 45724
rect 38172 45668 38176 45724
rect 38112 45664 38176 45668
rect 38192 45724 38256 45728
rect 38192 45668 38196 45724
rect 38196 45668 38252 45724
rect 38252 45668 38256 45724
rect 38192 45664 38256 45668
rect 47952 45724 48016 45728
rect 47952 45668 47956 45724
rect 47956 45668 48012 45724
rect 48012 45668 48016 45724
rect 47952 45664 48016 45668
rect 48032 45724 48096 45728
rect 48032 45668 48036 45724
rect 48036 45668 48092 45724
rect 48092 45668 48096 45724
rect 48032 45664 48096 45668
rect 48112 45724 48176 45728
rect 48112 45668 48116 45724
rect 48116 45668 48172 45724
rect 48172 45668 48176 45724
rect 48112 45664 48176 45668
rect 48192 45724 48256 45728
rect 48192 45668 48196 45724
rect 48196 45668 48252 45724
rect 48252 45668 48256 45724
rect 48192 45664 48256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 32952 45180 33016 45184
rect 32952 45124 32956 45180
rect 32956 45124 33012 45180
rect 33012 45124 33016 45180
rect 32952 45120 33016 45124
rect 33032 45180 33096 45184
rect 33032 45124 33036 45180
rect 33036 45124 33092 45180
rect 33092 45124 33096 45180
rect 33032 45120 33096 45124
rect 33112 45180 33176 45184
rect 33112 45124 33116 45180
rect 33116 45124 33172 45180
rect 33172 45124 33176 45180
rect 33112 45120 33176 45124
rect 33192 45180 33256 45184
rect 33192 45124 33196 45180
rect 33196 45124 33252 45180
rect 33252 45124 33256 45180
rect 33192 45120 33256 45124
rect 42952 45180 43016 45184
rect 42952 45124 42956 45180
rect 42956 45124 43012 45180
rect 43012 45124 43016 45180
rect 42952 45120 43016 45124
rect 43032 45180 43096 45184
rect 43032 45124 43036 45180
rect 43036 45124 43092 45180
rect 43092 45124 43096 45180
rect 43032 45120 43096 45124
rect 43112 45180 43176 45184
rect 43112 45124 43116 45180
rect 43116 45124 43172 45180
rect 43172 45124 43176 45180
rect 43112 45120 43176 45124
rect 43192 45180 43256 45184
rect 43192 45124 43196 45180
rect 43196 45124 43252 45180
rect 43252 45124 43256 45180
rect 43192 45120 43256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 27952 44636 28016 44640
rect 27952 44580 27956 44636
rect 27956 44580 28012 44636
rect 28012 44580 28016 44636
rect 27952 44576 28016 44580
rect 28032 44636 28096 44640
rect 28032 44580 28036 44636
rect 28036 44580 28092 44636
rect 28092 44580 28096 44636
rect 28032 44576 28096 44580
rect 28112 44636 28176 44640
rect 28112 44580 28116 44636
rect 28116 44580 28172 44636
rect 28172 44580 28176 44636
rect 28112 44576 28176 44580
rect 28192 44636 28256 44640
rect 28192 44580 28196 44636
rect 28196 44580 28252 44636
rect 28252 44580 28256 44636
rect 28192 44576 28256 44580
rect 37952 44636 38016 44640
rect 37952 44580 37956 44636
rect 37956 44580 38012 44636
rect 38012 44580 38016 44636
rect 37952 44576 38016 44580
rect 38032 44636 38096 44640
rect 38032 44580 38036 44636
rect 38036 44580 38092 44636
rect 38092 44580 38096 44636
rect 38032 44576 38096 44580
rect 38112 44636 38176 44640
rect 38112 44580 38116 44636
rect 38116 44580 38172 44636
rect 38172 44580 38176 44636
rect 38112 44576 38176 44580
rect 38192 44636 38256 44640
rect 38192 44580 38196 44636
rect 38196 44580 38252 44636
rect 38252 44580 38256 44636
rect 38192 44576 38256 44580
rect 47952 44636 48016 44640
rect 47952 44580 47956 44636
rect 47956 44580 48012 44636
rect 48012 44580 48016 44636
rect 47952 44576 48016 44580
rect 48032 44636 48096 44640
rect 48032 44580 48036 44636
rect 48036 44580 48092 44636
rect 48092 44580 48096 44636
rect 48032 44576 48096 44580
rect 48112 44636 48176 44640
rect 48112 44580 48116 44636
rect 48116 44580 48172 44636
rect 48172 44580 48176 44636
rect 48112 44576 48176 44580
rect 48192 44636 48256 44640
rect 48192 44580 48196 44636
rect 48196 44580 48252 44636
rect 48252 44580 48256 44636
rect 48192 44576 48256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 32952 44092 33016 44096
rect 32952 44036 32956 44092
rect 32956 44036 33012 44092
rect 33012 44036 33016 44092
rect 32952 44032 33016 44036
rect 33032 44092 33096 44096
rect 33032 44036 33036 44092
rect 33036 44036 33092 44092
rect 33092 44036 33096 44092
rect 33032 44032 33096 44036
rect 33112 44092 33176 44096
rect 33112 44036 33116 44092
rect 33116 44036 33172 44092
rect 33172 44036 33176 44092
rect 33112 44032 33176 44036
rect 33192 44092 33256 44096
rect 33192 44036 33196 44092
rect 33196 44036 33252 44092
rect 33252 44036 33256 44092
rect 33192 44032 33256 44036
rect 42952 44092 43016 44096
rect 42952 44036 42956 44092
rect 42956 44036 43012 44092
rect 43012 44036 43016 44092
rect 42952 44032 43016 44036
rect 43032 44092 43096 44096
rect 43032 44036 43036 44092
rect 43036 44036 43092 44092
rect 43092 44036 43096 44092
rect 43032 44032 43096 44036
rect 43112 44092 43176 44096
rect 43112 44036 43116 44092
rect 43116 44036 43172 44092
rect 43172 44036 43176 44092
rect 43112 44032 43176 44036
rect 43192 44092 43256 44096
rect 43192 44036 43196 44092
rect 43196 44036 43252 44092
rect 43252 44036 43256 44092
rect 43192 44032 43256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 27952 43548 28016 43552
rect 27952 43492 27956 43548
rect 27956 43492 28012 43548
rect 28012 43492 28016 43548
rect 27952 43488 28016 43492
rect 28032 43548 28096 43552
rect 28032 43492 28036 43548
rect 28036 43492 28092 43548
rect 28092 43492 28096 43548
rect 28032 43488 28096 43492
rect 28112 43548 28176 43552
rect 28112 43492 28116 43548
rect 28116 43492 28172 43548
rect 28172 43492 28176 43548
rect 28112 43488 28176 43492
rect 28192 43548 28256 43552
rect 28192 43492 28196 43548
rect 28196 43492 28252 43548
rect 28252 43492 28256 43548
rect 28192 43488 28256 43492
rect 37952 43548 38016 43552
rect 37952 43492 37956 43548
rect 37956 43492 38012 43548
rect 38012 43492 38016 43548
rect 37952 43488 38016 43492
rect 38032 43548 38096 43552
rect 38032 43492 38036 43548
rect 38036 43492 38092 43548
rect 38092 43492 38096 43548
rect 38032 43488 38096 43492
rect 38112 43548 38176 43552
rect 38112 43492 38116 43548
rect 38116 43492 38172 43548
rect 38172 43492 38176 43548
rect 38112 43488 38176 43492
rect 38192 43548 38256 43552
rect 38192 43492 38196 43548
rect 38196 43492 38252 43548
rect 38252 43492 38256 43548
rect 38192 43488 38256 43492
rect 47952 43548 48016 43552
rect 47952 43492 47956 43548
rect 47956 43492 48012 43548
rect 48012 43492 48016 43548
rect 47952 43488 48016 43492
rect 48032 43548 48096 43552
rect 48032 43492 48036 43548
rect 48036 43492 48092 43548
rect 48092 43492 48096 43548
rect 48032 43488 48096 43492
rect 48112 43548 48176 43552
rect 48112 43492 48116 43548
rect 48116 43492 48172 43548
rect 48172 43492 48176 43548
rect 48112 43488 48176 43492
rect 48192 43548 48256 43552
rect 48192 43492 48196 43548
rect 48196 43492 48252 43548
rect 48252 43492 48256 43548
rect 48192 43488 48256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 32952 43004 33016 43008
rect 32952 42948 32956 43004
rect 32956 42948 33012 43004
rect 33012 42948 33016 43004
rect 32952 42944 33016 42948
rect 33032 43004 33096 43008
rect 33032 42948 33036 43004
rect 33036 42948 33092 43004
rect 33092 42948 33096 43004
rect 33032 42944 33096 42948
rect 33112 43004 33176 43008
rect 33112 42948 33116 43004
rect 33116 42948 33172 43004
rect 33172 42948 33176 43004
rect 33112 42944 33176 42948
rect 33192 43004 33256 43008
rect 33192 42948 33196 43004
rect 33196 42948 33252 43004
rect 33252 42948 33256 43004
rect 33192 42944 33256 42948
rect 42952 43004 43016 43008
rect 42952 42948 42956 43004
rect 42956 42948 43012 43004
rect 43012 42948 43016 43004
rect 42952 42944 43016 42948
rect 43032 43004 43096 43008
rect 43032 42948 43036 43004
rect 43036 42948 43092 43004
rect 43092 42948 43096 43004
rect 43032 42944 43096 42948
rect 43112 43004 43176 43008
rect 43112 42948 43116 43004
rect 43116 42948 43172 43004
rect 43172 42948 43176 43004
rect 43112 42944 43176 42948
rect 43192 43004 43256 43008
rect 43192 42948 43196 43004
rect 43196 42948 43252 43004
rect 43252 42948 43256 43004
rect 43192 42944 43256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 27952 42460 28016 42464
rect 27952 42404 27956 42460
rect 27956 42404 28012 42460
rect 28012 42404 28016 42460
rect 27952 42400 28016 42404
rect 28032 42460 28096 42464
rect 28032 42404 28036 42460
rect 28036 42404 28092 42460
rect 28092 42404 28096 42460
rect 28032 42400 28096 42404
rect 28112 42460 28176 42464
rect 28112 42404 28116 42460
rect 28116 42404 28172 42460
rect 28172 42404 28176 42460
rect 28112 42400 28176 42404
rect 28192 42460 28256 42464
rect 28192 42404 28196 42460
rect 28196 42404 28252 42460
rect 28252 42404 28256 42460
rect 28192 42400 28256 42404
rect 37952 42460 38016 42464
rect 37952 42404 37956 42460
rect 37956 42404 38012 42460
rect 38012 42404 38016 42460
rect 37952 42400 38016 42404
rect 38032 42460 38096 42464
rect 38032 42404 38036 42460
rect 38036 42404 38092 42460
rect 38092 42404 38096 42460
rect 38032 42400 38096 42404
rect 38112 42460 38176 42464
rect 38112 42404 38116 42460
rect 38116 42404 38172 42460
rect 38172 42404 38176 42460
rect 38112 42400 38176 42404
rect 38192 42460 38256 42464
rect 38192 42404 38196 42460
rect 38196 42404 38252 42460
rect 38252 42404 38256 42460
rect 38192 42400 38256 42404
rect 47952 42460 48016 42464
rect 47952 42404 47956 42460
rect 47956 42404 48012 42460
rect 48012 42404 48016 42460
rect 47952 42400 48016 42404
rect 48032 42460 48096 42464
rect 48032 42404 48036 42460
rect 48036 42404 48092 42460
rect 48092 42404 48096 42460
rect 48032 42400 48096 42404
rect 48112 42460 48176 42464
rect 48112 42404 48116 42460
rect 48116 42404 48172 42460
rect 48172 42404 48176 42460
rect 48112 42400 48176 42404
rect 48192 42460 48256 42464
rect 48192 42404 48196 42460
rect 48196 42404 48252 42460
rect 48252 42404 48256 42460
rect 48192 42400 48256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 32952 41916 33016 41920
rect 32952 41860 32956 41916
rect 32956 41860 33012 41916
rect 33012 41860 33016 41916
rect 32952 41856 33016 41860
rect 33032 41916 33096 41920
rect 33032 41860 33036 41916
rect 33036 41860 33092 41916
rect 33092 41860 33096 41916
rect 33032 41856 33096 41860
rect 33112 41916 33176 41920
rect 33112 41860 33116 41916
rect 33116 41860 33172 41916
rect 33172 41860 33176 41916
rect 33112 41856 33176 41860
rect 33192 41916 33256 41920
rect 33192 41860 33196 41916
rect 33196 41860 33252 41916
rect 33252 41860 33256 41916
rect 33192 41856 33256 41860
rect 42952 41916 43016 41920
rect 42952 41860 42956 41916
rect 42956 41860 43012 41916
rect 43012 41860 43016 41916
rect 42952 41856 43016 41860
rect 43032 41916 43096 41920
rect 43032 41860 43036 41916
rect 43036 41860 43092 41916
rect 43092 41860 43096 41916
rect 43032 41856 43096 41860
rect 43112 41916 43176 41920
rect 43112 41860 43116 41916
rect 43116 41860 43172 41916
rect 43172 41860 43176 41916
rect 43112 41856 43176 41860
rect 43192 41916 43256 41920
rect 43192 41860 43196 41916
rect 43196 41860 43252 41916
rect 43252 41860 43256 41916
rect 43192 41856 43256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 27952 41372 28016 41376
rect 27952 41316 27956 41372
rect 27956 41316 28012 41372
rect 28012 41316 28016 41372
rect 27952 41312 28016 41316
rect 28032 41372 28096 41376
rect 28032 41316 28036 41372
rect 28036 41316 28092 41372
rect 28092 41316 28096 41372
rect 28032 41312 28096 41316
rect 28112 41372 28176 41376
rect 28112 41316 28116 41372
rect 28116 41316 28172 41372
rect 28172 41316 28176 41372
rect 28112 41312 28176 41316
rect 28192 41372 28256 41376
rect 28192 41316 28196 41372
rect 28196 41316 28252 41372
rect 28252 41316 28256 41372
rect 28192 41312 28256 41316
rect 37952 41372 38016 41376
rect 37952 41316 37956 41372
rect 37956 41316 38012 41372
rect 38012 41316 38016 41372
rect 37952 41312 38016 41316
rect 38032 41372 38096 41376
rect 38032 41316 38036 41372
rect 38036 41316 38092 41372
rect 38092 41316 38096 41372
rect 38032 41312 38096 41316
rect 38112 41372 38176 41376
rect 38112 41316 38116 41372
rect 38116 41316 38172 41372
rect 38172 41316 38176 41372
rect 38112 41312 38176 41316
rect 38192 41372 38256 41376
rect 38192 41316 38196 41372
rect 38196 41316 38252 41372
rect 38252 41316 38256 41372
rect 38192 41312 38256 41316
rect 47952 41372 48016 41376
rect 47952 41316 47956 41372
rect 47956 41316 48012 41372
rect 48012 41316 48016 41372
rect 47952 41312 48016 41316
rect 48032 41372 48096 41376
rect 48032 41316 48036 41372
rect 48036 41316 48092 41372
rect 48092 41316 48096 41372
rect 48032 41312 48096 41316
rect 48112 41372 48176 41376
rect 48112 41316 48116 41372
rect 48116 41316 48172 41372
rect 48172 41316 48176 41372
rect 48112 41312 48176 41316
rect 48192 41372 48256 41376
rect 48192 41316 48196 41372
rect 48196 41316 48252 41372
rect 48252 41316 48256 41372
rect 48192 41312 48256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 32952 40828 33016 40832
rect 32952 40772 32956 40828
rect 32956 40772 33012 40828
rect 33012 40772 33016 40828
rect 32952 40768 33016 40772
rect 33032 40828 33096 40832
rect 33032 40772 33036 40828
rect 33036 40772 33092 40828
rect 33092 40772 33096 40828
rect 33032 40768 33096 40772
rect 33112 40828 33176 40832
rect 33112 40772 33116 40828
rect 33116 40772 33172 40828
rect 33172 40772 33176 40828
rect 33112 40768 33176 40772
rect 33192 40828 33256 40832
rect 33192 40772 33196 40828
rect 33196 40772 33252 40828
rect 33252 40772 33256 40828
rect 33192 40768 33256 40772
rect 42952 40828 43016 40832
rect 42952 40772 42956 40828
rect 42956 40772 43012 40828
rect 43012 40772 43016 40828
rect 42952 40768 43016 40772
rect 43032 40828 43096 40832
rect 43032 40772 43036 40828
rect 43036 40772 43092 40828
rect 43092 40772 43096 40828
rect 43032 40768 43096 40772
rect 43112 40828 43176 40832
rect 43112 40772 43116 40828
rect 43116 40772 43172 40828
rect 43172 40772 43176 40828
rect 43112 40768 43176 40772
rect 43192 40828 43256 40832
rect 43192 40772 43196 40828
rect 43196 40772 43252 40828
rect 43252 40772 43256 40828
rect 43192 40768 43256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 27952 40284 28016 40288
rect 27952 40228 27956 40284
rect 27956 40228 28012 40284
rect 28012 40228 28016 40284
rect 27952 40224 28016 40228
rect 28032 40284 28096 40288
rect 28032 40228 28036 40284
rect 28036 40228 28092 40284
rect 28092 40228 28096 40284
rect 28032 40224 28096 40228
rect 28112 40284 28176 40288
rect 28112 40228 28116 40284
rect 28116 40228 28172 40284
rect 28172 40228 28176 40284
rect 28112 40224 28176 40228
rect 28192 40284 28256 40288
rect 28192 40228 28196 40284
rect 28196 40228 28252 40284
rect 28252 40228 28256 40284
rect 28192 40224 28256 40228
rect 37952 40284 38016 40288
rect 37952 40228 37956 40284
rect 37956 40228 38012 40284
rect 38012 40228 38016 40284
rect 37952 40224 38016 40228
rect 38032 40284 38096 40288
rect 38032 40228 38036 40284
rect 38036 40228 38092 40284
rect 38092 40228 38096 40284
rect 38032 40224 38096 40228
rect 38112 40284 38176 40288
rect 38112 40228 38116 40284
rect 38116 40228 38172 40284
rect 38172 40228 38176 40284
rect 38112 40224 38176 40228
rect 38192 40284 38256 40288
rect 38192 40228 38196 40284
rect 38196 40228 38252 40284
rect 38252 40228 38256 40284
rect 38192 40224 38256 40228
rect 47952 40284 48016 40288
rect 47952 40228 47956 40284
rect 47956 40228 48012 40284
rect 48012 40228 48016 40284
rect 47952 40224 48016 40228
rect 48032 40284 48096 40288
rect 48032 40228 48036 40284
rect 48036 40228 48092 40284
rect 48092 40228 48096 40284
rect 48032 40224 48096 40228
rect 48112 40284 48176 40288
rect 48112 40228 48116 40284
rect 48116 40228 48172 40284
rect 48172 40228 48176 40284
rect 48112 40224 48176 40228
rect 48192 40284 48256 40288
rect 48192 40228 48196 40284
rect 48196 40228 48252 40284
rect 48252 40228 48256 40284
rect 48192 40224 48256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 32952 39740 33016 39744
rect 32952 39684 32956 39740
rect 32956 39684 33012 39740
rect 33012 39684 33016 39740
rect 32952 39680 33016 39684
rect 33032 39740 33096 39744
rect 33032 39684 33036 39740
rect 33036 39684 33092 39740
rect 33092 39684 33096 39740
rect 33032 39680 33096 39684
rect 33112 39740 33176 39744
rect 33112 39684 33116 39740
rect 33116 39684 33172 39740
rect 33172 39684 33176 39740
rect 33112 39680 33176 39684
rect 33192 39740 33256 39744
rect 33192 39684 33196 39740
rect 33196 39684 33252 39740
rect 33252 39684 33256 39740
rect 33192 39680 33256 39684
rect 42952 39740 43016 39744
rect 42952 39684 42956 39740
rect 42956 39684 43012 39740
rect 43012 39684 43016 39740
rect 42952 39680 43016 39684
rect 43032 39740 43096 39744
rect 43032 39684 43036 39740
rect 43036 39684 43092 39740
rect 43092 39684 43096 39740
rect 43032 39680 43096 39684
rect 43112 39740 43176 39744
rect 43112 39684 43116 39740
rect 43116 39684 43172 39740
rect 43172 39684 43176 39740
rect 43112 39680 43176 39684
rect 43192 39740 43256 39744
rect 43192 39684 43196 39740
rect 43196 39684 43252 39740
rect 43252 39684 43256 39740
rect 43192 39680 43256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 27952 39196 28016 39200
rect 27952 39140 27956 39196
rect 27956 39140 28012 39196
rect 28012 39140 28016 39196
rect 27952 39136 28016 39140
rect 28032 39196 28096 39200
rect 28032 39140 28036 39196
rect 28036 39140 28092 39196
rect 28092 39140 28096 39196
rect 28032 39136 28096 39140
rect 28112 39196 28176 39200
rect 28112 39140 28116 39196
rect 28116 39140 28172 39196
rect 28172 39140 28176 39196
rect 28112 39136 28176 39140
rect 28192 39196 28256 39200
rect 28192 39140 28196 39196
rect 28196 39140 28252 39196
rect 28252 39140 28256 39196
rect 28192 39136 28256 39140
rect 37952 39196 38016 39200
rect 37952 39140 37956 39196
rect 37956 39140 38012 39196
rect 38012 39140 38016 39196
rect 37952 39136 38016 39140
rect 38032 39196 38096 39200
rect 38032 39140 38036 39196
rect 38036 39140 38092 39196
rect 38092 39140 38096 39196
rect 38032 39136 38096 39140
rect 38112 39196 38176 39200
rect 38112 39140 38116 39196
rect 38116 39140 38172 39196
rect 38172 39140 38176 39196
rect 38112 39136 38176 39140
rect 38192 39196 38256 39200
rect 38192 39140 38196 39196
rect 38196 39140 38252 39196
rect 38252 39140 38256 39196
rect 38192 39136 38256 39140
rect 47952 39196 48016 39200
rect 47952 39140 47956 39196
rect 47956 39140 48012 39196
rect 48012 39140 48016 39196
rect 47952 39136 48016 39140
rect 48032 39196 48096 39200
rect 48032 39140 48036 39196
rect 48036 39140 48092 39196
rect 48092 39140 48096 39196
rect 48032 39136 48096 39140
rect 48112 39196 48176 39200
rect 48112 39140 48116 39196
rect 48116 39140 48172 39196
rect 48172 39140 48176 39196
rect 48112 39136 48176 39140
rect 48192 39196 48256 39200
rect 48192 39140 48196 39196
rect 48196 39140 48252 39196
rect 48252 39140 48256 39196
rect 48192 39136 48256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 32952 38652 33016 38656
rect 32952 38596 32956 38652
rect 32956 38596 33012 38652
rect 33012 38596 33016 38652
rect 32952 38592 33016 38596
rect 33032 38652 33096 38656
rect 33032 38596 33036 38652
rect 33036 38596 33092 38652
rect 33092 38596 33096 38652
rect 33032 38592 33096 38596
rect 33112 38652 33176 38656
rect 33112 38596 33116 38652
rect 33116 38596 33172 38652
rect 33172 38596 33176 38652
rect 33112 38592 33176 38596
rect 33192 38652 33256 38656
rect 33192 38596 33196 38652
rect 33196 38596 33252 38652
rect 33252 38596 33256 38652
rect 33192 38592 33256 38596
rect 42952 38652 43016 38656
rect 42952 38596 42956 38652
rect 42956 38596 43012 38652
rect 43012 38596 43016 38652
rect 42952 38592 43016 38596
rect 43032 38652 43096 38656
rect 43032 38596 43036 38652
rect 43036 38596 43092 38652
rect 43092 38596 43096 38652
rect 43032 38592 43096 38596
rect 43112 38652 43176 38656
rect 43112 38596 43116 38652
rect 43116 38596 43172 38652
rect 43172 38596 43176 38652
rect 43112 38592 43176 38596
rect 43192 38652 43256 38656
rect 43192 38596 43196 38652
rect 43196 38596 43252 38652
rect 43252 38596 43256 38652
rect 43192 38592 43256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 27952 38108 28016 38112
rect 27952 38052 27956 38108
rect 27956 38052 28012 38108
rect 28012 38052 28016 38108
rect 27952 38048 28016 38052
rect 28032 38108 28096 38112
rect 28032 38052 28036 38108
rect 28036 38052 28092 38108
rect 28092 38052 28096 38108
rect 28032 38048 28096 38052
rect 28112 38108 28176 38112
rect 28112 38052 28116 38108
rect 28116 38052 28172 38108
rect 28172 38052 28176 38108
rect 28112 38048 28176 38052
rect 28192 38108 28256 38112
rect 28192 38052 28196 38108
rect 28196 38052 28252 38108
rect 28252 38052 28256 38108
rect 28192 38048 28256 38052
rect 37952 38108 38016 38112
rect 37952 38052 37956 38108
rect 37956 38052 38012 38108
rect 38012 38052 38016 38108
rect 37952 38048 38016 38052
rect 38032 38108 38096 38112
rect 38032 38052 38036 38108
rect 38036 38052 38092 38108
rect 38092 38052 38096 38108
rect 38032 38048 38096 38052
rect 38112 38108 38176 38112
rect 38112 38052 38116 38108
rect 38116 38052 38172 38108
rect 38172 38052 38176 38108
rect 38112 38048 38176 38052
rect 38192 38108 38256 38112
rect 38192 38052 38196 38108
rect 38196 38052 38252 38108
rect 38252 38052 38256 38108
rect 38192 38048 38256 38052
rect 47952 38108 48016 38112
rect 47952 38052 47956 38108
rect 47956 38052 48012 38108
rect 48012 38052 48016 38108
rect 47952 38048 48016 38052
rect 48032 38108 48096 38112
rect 48032 38052 48036 38108
rect 48036 38052 48092 38108
rect 48092 38052 48096 38108
rect 48032 38048 48096 38052
rect 48112 38108 48176 38112
rect 48112 38052 48116 38108
rect 48116 38052 48172 38108
rect 48172 38052 48176 38108
rect 48112 38048 48176 38052
rect 48192 38108 48256 38112
rect 48192 38052 48196 38108
rect 48196 38052 48252 38108
rect 48252 38052 48256 38108
rect 48192 38048 48256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 32952 37564 33016 37568
rect 32952 37508 32956 37564
rect 32956 37508 33012 37564
rect 33012 37508 33016 37564
rect 32952 37504 33016 37508
rect 33032 37564 33096 37568
rect 33032 37508 33036 37564
rect 33036 37508 33092 37564
rect 33092 37508 33096 37564
rect 33032 37504 33096 37508
rect 33112 37564 33176 37568
rect 33112 37508 33116 37564
rect 33116 37508 33172 37564
rect 33172 37508 33176 37564
rect 33112 37504 33176 37508
rect 33192 37564 33256 37568
rect 33192 37508 33196 37564
rect 33196 37508 33252 37564
rect 33252 37508 33256 37564
rect 33192 37504 33256 37508
rect 42952 37564 43016 37568
rect 42952 37508 42956 37564
rect 42956 37508 43012 37564
rect 43012 37508 43016 37564
rect 42952 37504 43016 37508
rect 43032 37564 43096 37568
rect 43032 37508 43036 37564
rect 43036 37508 43092 37564
rect 43092 37508 43096 37564
rect 43032 37504 43096 37508
rect 43112 37564 43176 37568
rect 43112 37508 43116 37564
rect 43116 37508 43172 37564
rect 43172 37508 43176 37564
rect 43112 37504 43176 37508
rect 43192 37564 43256 37568
rect 43192 37508 43196 37564
rect 43196 37508 43252 37564
rect 43252 37508 43256 37564
rect 43192 37504 43256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 27952 37020 28016 37024
rect 27952 36964 27956 37020
rect 27956 36964 28012 37020
rect 28012 36964 28016 37020
rect 27952 36960 28016 36964
rect 28032 37020 28096 37024
rect 28032 36964 28036 37020
rect 28036 36964 28092 37020
rect 28092 36964 28096 37020
rect 28032 36960 28096 36964
rect 28112 37020 28176 37024
rect 28112 36964 28116 37020
rect 28116 36964 28172 37020
rect 28172 36964 28176 37020
rect 28112 36960 28176 36964
rect 28192 37020 28256 37024
rect 28192 36964 28196 37020
rect 28196 36964 28252 37020
rect 28252 36964 28256 37020
rect 28192 36960 28256 36964
rect 37952 37020 38016 37024
rect 37952 36964 37956 37020
rect 37956 36964 38012 37020
rect 38012 36964 38016 37020
rect 37952 36960 38016 36964
rect 38032 37020 38096 37024
rect 38032 36964 38036 37020
rect 38036 36964 38092 37020
rect 38092 36964 38096 37020
rect 38032 36960 38096 36964
rect 38112 37020 38176 37024
rect 38112 36964 38116 37020
rect 38116 36964 38172 37020
rect 38172 36964 38176 37020
rect 38112 36960 38176 36964
rect 38192 37020 38256 37024
rect 38192 36964 38196 37020
rect 38196 36964 38252 37020
rect 38252 36964 38256 37020
rect 38192 36960 38256 36964
rect 47952 37020 48016 37024
rect 47952 36964 47956 37020
rect 47956 36964 48012 37020
rect 48012 36964 48016 37020
rect 47952 36960 48016 36964
rect 48032 37020 48096 37024
rect 48032 36964 48036 37020
rect 48036 36964 48092 37020
rect 48092 36964 48096 37020
rect 48032 36960 48096 36964
rect 48112 37020 48176 37024
rect 48112 36964 48116 37020
rect 48116 36964 48172 37020
rect 48172 36964 48176 37020
rect 48112 36960 48176 36964
rect 48192 37020 48256 37024
rect 48192 36964 48196 37020
rect 48196 36964 48252 37020
rect 48252 36964 48256 37020
rect 48192 36960 48256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 32952 36476 33016 36480
rect 32952 36420 32956 36476
rect 32956 36420 33012 36476
rect 33012 36420 33016 36476
rect 32952 36416 33016 36420
rect 33032 36476 33096 36480
rect 33032 36420 33036 36476
rect 33036 36420 33092 36476
rect 33092 36420 33096 36476
rect 33032 36416 33096 36420
rect 33112 36476 33176 36480
rect 33112 36420 33116 36476
rect 33116 36420 33172 36476
rect 33172 36420 33176 36476
rect 33112 36416 33176 36420
rect 33192 36476 33256 36480
rect 33192 36420 33196 36476
rect 33196 36420 33252 36476
rect 33252 36420 33256 36476
rect 33192 36416 33256 36420
rect 42952 36476 43016 36480
rect 42952 36420 42956 36476
rect 42956 36420 43012 36476
rect 43012 36420 43016 36476
rect 42952 36416 43016 36420
rect 43032 36476 43096 36480
rect 43032 36420 43036 36476
rect 43036 36420 43092 36476
rect 43092 36420 43096 36476
rect 43032 36416 43096 36420
rect 43112 36476 43176 36480
rect 43112 36420 43116 36476
rect 43116 36420 43172 36476
rect 43172 36420 43176 36476
rect 43112 36416 43176 36420
rect 43192 36476 43256 36480
rect 43192 36420 43196 36476
rect 43196 36420 43252 36476
rect 43252 36420 43256 36476
rect 43192 36416 43256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 27952 35932 28016 35936
rect 27952 35876 27956 35932
rect 27956 35876 28012 35932
rect 28012 35876 28016 35932
rect 27952 35872 28016 35876
rect 28032 35932 28096 35936
rect 28032 35876 28036 35932
rect 28036 35876 28092 35932
rect 28092 35876 28096 35932
rect 28032 35872 28096 35876
rect 28112 35932 28176 35936
rect 28112 35876 28116 35932
rect 28116 35876 28172 35932
rect 28172 35876 28176 35932
rect 28112 35872 28176 35876
rect 28192 35932 28256 35936
rect 28192 35876 28196 35932
rect 28196 35876 28252 35932
rect 28252 35876 28256 35932
rect 28192 35872 28256 35876
rect 37952 35932 38016 35936
rect 37952 35876 37956 35932
rect 37956 35876 38012 35932
rect 38012 35876 38016 35932
rect 37952 35872 38016 35876
rect 38032 35932 38096 35936
rect 38032 35876 38036 35932
rect 38036 35876 38092 35932
rect 38092 35876 38096 35932
rect 38032 35872 38096 35876
rect 38112 35932 38176 35936
rect 38112 35876 38116 35932
rect 38116 35876 38172 35932
rect 38172 35876 38176 35932
rect 38112 35872 38176 35876
rect 38192 35932 38256 35936
rect 38192 35876 38196 35932
rect 38196 35876 38252 35932
rect 38252 35876 38256 35932
rect 38192 35872 38256 35876
rect 47952 35932 48016 35936
rect 47952 35876 47956 35932
rect 47956 35876 48012 35932
rect 48012 35876 48016 35932
rect 47952 35872 48016 35876
rect 48032 35932 48096 35936
rect 48032 35876 48036 35932
rect 48036 35876 48092 35932
rect 48092 35876 48096 35932
rect 48032 35872 48096 35876
rect 48112 35932 48176 35936
rect 48112 35876 48116 35932
rect 48116 35876 48172 35932
rect 48172 35876 48176 35932
rect 48112 35872 48176 35876
rect 48192 35932 48256 35936
rect 48192 35876 48196 35932
rect 48196 35876 48252 35932
rect 48252 35876 48256 35932
rect 48192 35872 48256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 32952 35388 33016 35392
rect 32952 35332 32956 35388
rect 32956 35332 33012 35388
rect 33012 35332 33016 35388
rect 32952 35328 33016 35332
rect 33032 35388 33096 35392
rect 33032 35332 33036 35388
rect 33036 35332 33092 35388
rect 33092 35332 33096 35388
rect 33032 35328 33096 35332
rect 33112 35388 33176 35392
rect 33112 35332 33116 35388
rect 33116 35332 33172 35388
rect 33172 35332 33176 35388
rect 33112 35328 33176 35332
rect 33192 35388 33256 35392
rect 33192 35332 33196 35388
rect 33196 35332 33252 35388
rect 33252 35332 33256 35388
rect 33192 35328 33256 35332
rect 42952 35388 43016 35392
rect 42952 35332 42956 35388
rect 42956 35332 43012 35388
rect 43012 35332 43016 35388
rect 42952 35328 43016 35332
rect 43032 35388 43096 35392
rect 43032 35332 43036 35388
rect 43036 35332 43092 35388
rect 43092 35332 43096 35388
rect 43032 35328 43096 35332
rect 43112 35388 43176 35392
rect 43112 35332 43116 35388
rect 43116 35332 43172 35388
rect 43172 35332 43176 35388
rect 43112 35328 43176 35332
rect 43192 35388 43256 35392
rect 43192 35332 43196 35388
rect 43196 35332 43252 35388
rect 43252 35332 43256 35388
rect 43192 35328 43256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 27952 34844 28016 34848
rect 27952 34788 27956 34844
rect 27956 34788 28012 34844
rect 28012 34788 28016 34844
rect 27952 34784 28016 34788
rect 28032 34844 28096 34848
rect 28032 34788 28036 34844
rect 28036 34788 28092 34844
rect 28092 34788 28096 34844
rect 28032 34784 28096 34788
rect 28112 34844 28176 34848
rect 28112 34788 28116 34844
rect 28116 34788 28172 34844
rect 28172 34788 28176 34844
rect 28112 34784 28176 34788
rect 28192 34844 28256 34848
rect 28192 34788 28196 34844
rect 28196 34788 28252 34844
rect 28252 34788 28256 34844
rect 28192 34784 28256 34788
rect 37952 34844 38016 34848
rect 37952 34788 37956 34844
rect 37956 34788 38012 34844
rect 38012 34788 38016 34844
rect 37952 34784 38016 34788
rect 38032 34844 38096 34848
rect 38032 34788 38036 34844
rect 38036 34788 38092 34844
rect 38092 34788 38096 34844
rect 38032 34784 38096 34788
rect 38112 34844 38176 34848
rect 38112 34788 38116 34844
rect 38116 34788 38172 34844
rect 38172 34788 38176 34844
rect 38112 34784 38176 34788
rect 38192 34844 38256 34848
rect 38192 34788 38196 34844
rect 38196 34788 38252 34844
rect 38252 34788 38256 34844
rect 38192 34784 38256 34788
rect 47952 34844 48016 34848
rect 47952 34788 47956 34844
rect 47956 34788 48012 34844
rect 48012 34788 48016 34844
rect 47952 34784 48016 34788
rect 48032 34844 48096 34848
rect 48032 34788 48036 34844
rect 48036 34788 48092 34844
rect 48092 34788 48096 34844
rect 48032 34784 48096 34788
rect 48112 34844 48176 34848
rect 48112 34788 48116 34844
rect 48116 34788 48172 34844
rect 48172 34788 48176 34844
rect 48112 34784 48176 34788
rect 48192 34844 48256 34848
rect 48192 34788 48196 34844
rect 48196 34788 48252 34844
rect 48252 34788 48256 34844
rect 48192 34784 48256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 32952 34300 33016 34304
rect 32952 34244 32956 34300
rect 32956 34244 33012 34300
rect 33012 34244 33016 34300
rect 32952 34240 33016 34244
rect 33032 34300 33096 34304
rect 33032 34244 33036 34300
rect 33036 34244 33092 34300
rect 33092 34244 33096 34300
rect 33032 34240 33096 34244
rect 33112 34300 33176 34304
rect 33112 34244 33116 34300
rect 33116 34244 33172 34300
rect 33172 34244 33176 34300
rect 33112 34240 33176 34244
rect 33192 34300 33256 34304
rect 33192 34244 33196 34300
rect 33196 34244 33252 34300
rect 33252 34244 33256 34300
rect 33192 34240 33256 34244
rect 42952 34300 43016 34304
rect 42952 34244 42956 34300
rect 42956 34244 43012 34300
rect 43012 34244 43016 34300
rect 42952 34240 43016 34244
rect 43032 34300 43096 34304
rect 43032 34244 43036 34300
rect 43036 34244 43092 34300
rect 43092 34244 43096 34300
rect 43032 34240 43096 34244
rect 43112 34300 43176 34304
rect 43112 34244 43116 34300
rect 43116 34244 43172 34300
rect 43172 34244 43176 34300
rect 43112 34240 43176 34244
rect 43192 34300 43256 34304
rect 43192 34244 43196 34300
rect 43196 34244 43252 34300
rect 43252 34244 43256 34300
rect 43192 34240 43256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 27952 33756 28016 33760
rect 27952 33700 27956 33756
rect 27956 33700 28012 33756
rect 28012 33700 28016 33756
rect 27952 33696 28016 33700
rect 28032 33756 28096 33760
rect 28032 33700 28036 33756
rect 28036 33700 28092 33756
rect 28092 33700 28096 33756
rect 28032 33696 28096 33700
rect 28112 33756 28176 33760
rect 28112 33700 28116 33756
rect 28116 33700 28172 33756
rect 28172 33700 28176 33756
rect 28112 33696 28176 33700
rect 28192 33756 28256 33760
rect 28192 33700 28196 33756
rect 28196 33700 28252 33756
rect 28252 33700 28256 33756
rect 28192 33696 28256 33700
rect 37952 33756 38016 33760
rect 37952 33700 37956 33756
rect 37956 33700 38012 33756
rect 38012 33700 38016 33756
rect 37952 33696 38016 33700
rect 38032 33756 38096 33760
rect 38032 33700 38036 33756
rect 38036 33700 38092 33756
rect 38092 33700 38096 33756
rect 38032 33696 38096 33700
rect 38112 33756 38176 33760
rect 38112 33700 38116 33756
rect 38116 33700 38172 33756
rect 38172 33700 38176 33756
rect 38112 33696 38176 33700
rect 38192 33756 38256 33760
rect 38192 33700 38196 33756
rect 38196 33700 38252 33756
rect 38252 33700 38256 33756
rect 38192 33696 38256 33700
rect 47952 33756 48016 33760
rect 47952 33700 47956 33756
rect 47956 33700 48012 33756
rect 48012 33700 48016 33756
rect 47952 33696 48016 33700
rect 48032 33756 48096 33760
rect 48032 33700 48036 33756
rect 48036 33700 48092 33756
rect 48092 33700 48096 33756
rect 48032 33696 48096 33700
rect 48112 33756 48176 33760
rect 48112 33700 48116 33756
rect 48116 33700 48172 33756
rect 48172 33700 48176 33756
rect 48112 33696 48176 33700
rect 48192 33756 48256 33760
rect 48192 33700 48196 33756
rect 48196 33700 48252 33756
rect 48252 33700 48256 33756
rect 48192 33696 48256 33700
rect 26188 33628 26252 33692
rect 28580 33220 28644 33284
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 32952 33212 33016 33216
rect 32952 33156 32956 33212
rect 32956 33156 33012 33212
rect 33012 33156 33016 33212
rect 32952 33152 33016 33156
rect 33032 33212 33096 33216
rect 33032 33156 33036 33212
rect 33036 33156 33092 33212
rect 33092 33156 33096 33212
rect 33032 33152 33096 33156
rect 33112 33212 33176 33216
rect 33112 33156 33116 33212
rect 33116 33156 33172 33212
rect 33172 33156 33176 33212
rect 33112 33152 33176 33156
rect 33192 33212 33256 33216
rect 33192 33156 33196 33212
rect 33196 33156 33252 33212
rect 33252 33156 33256 33212
rect 33192 33152 33256 33156
rect 42952 33212 43016 33216
rect 42952 33156 42956 33212
rect 42956 33156 43012 33212
rect 43012 33156 43016 33212
rect 42952 33152 43016 33156
rect 43032 33212 43096 33216
rect 43032 33156 43036 33212
rect 43036 33156 43092 33212
rect 43092 33156 43096 33212
rect 43032 33152 43096 33156
rect 43112 33212 43176 33216
rect 43112 33156 43116 33212
rect 43116 33156 43172 33212
rect 43172 33156 43176 33212
rect 43112 33152 43176 33156
rect 43192 33212 43256 33216
rect 43192 33156 43196 33212
rect 43196 33156 43252 33212
rect 43252 33156 43256 33212
rect 43192 33152 43256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 27952 32668 28016 32672
rect 27952 32612 27956 32668
rect 27956 32612 28012 32668
rect 28012 32612 28016 32668
rect 27952 32608 28016 32612
rect 28032 32668 28096 32672
rect 28032 32612 28036 32668
rect 28036 32612 28092 32668
rect 28092 32612 28096 32668
rect 28032 32608 28096 32612
rect 28112 32668 28176 32672
rect 28112 32612 28116 32668
rect 28116 32612 28172 32668
rect 28172 32612 28176 32668
rect 28112 32608 28176 32612
rect 28192 32668 28256 32672
rect 28192 32612 28196 32668
rect 28196 32612 28252 32668
rect 28252 32612 28256 32668
rect 28192 32608 28256 32612
rect 37952 32668 38016 32672
rect 37952 32612 37956 32668
rect 37956 32612 38012 32668
rect 38012 32612 38016 32668
rect 37952 32608 38016 32612
rect 38032 32668 38096 32672
rect 38032 32612 38036 32668
rect 38036 32612 38092 32668
rect 38092 32612 38096 32668
rect 38032 32608 38096 32612
rect 38112 32668 38176 32672
rect 38112 32612 38116 32668
rect 38116 32612 38172 32668
rect 38172 32612 38176 32668
rect 38112 32608 38176 32612
rect 38192 32668 38256 32672
rect 38192 32612 38196 32668
rect 38196 32612 38252 32668
rect 38252 32612 38256 32668
rect 38192 32608 38256 32612
rect 47952 32668 48016 32672
rect 47952 32612 47956 32668
rect 47956 32612 48012 32668
rect 48012 32612 48016 32668
rect 47952 32608 48016 32612
rect 48032 32668 48096 32672
rect 48032 32612 48036 32668
rect 48036 32612 48092 32668
rect 48092 32612 48096 32668
rect 48032 32608 48096 32612
rect 48112 32668 48176 32672
rect 48112 32612 48116 32668
rect 48116 32612 48172 32668
rect 48172 32612 48176 32668
rect 48112 32608 48176 32612
rect 48192 32668 48256 32672
rect 48192 32612 48196 32668
rect 48196 32612 48252 32668
rect 48252 32612 48256 32668
rect 48192 32608 48256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 32952 32124 33016 32128
rect 32952 32068 32956 32124
rect 32956 32068 33012 32124
rect 33012 32068 33016 32124
rect 32952 32064 33016 32068
rect 33032 32124 33096 32128
rect 33032 32068 33036 32124
rect 33036 32068 33092 32124
rect 33092 32068 33096 32124
rect 33032 32064 33096 32068
rect 33112 32124 33176 32128
rect 33112 32068 33116 32124
rect 33116 32068 33172 32124
rect 33172 32068 33176 32124
rect 33112 32064 33176 32068
rect 33192 32124 33256 32128
rect 33192 32068 33196 32124
rect 33196 32068 33252 32124
rect 33252 32068 33256 32124
rect 33192 32064 33256 32068
rect 42952 32124 43016 32128
rect 42952 32068 42956 32124
rect 42956 32068 43012 32124
rect 43012 32068 43016 32124
rect 42952 32064 43016 32068
rect 43032 32124 43096 32128
rect 43032 32068 43036 32124
rect 43036 32068 43092 32124
rect 43092 32068 43096 32124
rect 43032 32064 43096 32068
rect 43112 32124 43176 32128
rect 43112 32068 43116 32124
rect 43116 32068 43172 32124
rect 43172 32068 43176 32124
rect 43112 32064 43176 32068
rect 43192 32124 43256 32128
rect 43192 32068 43196 32124
rect 43196 32068 43252 32124
rect 43252 32068 43256 32124
rect 43192 32064 43256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 27952 31580 28016 31584
rect 27952 31524 27956 31580
rect 27956 31524 28012 31580
rect 28012 31524 28016 31580
rect 27952 31520 28016 31524
rect 28032 31580 28096 31584
rect 28032 31524 28036 31580
rect 28036 31524 28092 31580
rect 28092 31524 28096 31580
rect 28032 31520 28096 31524
rect 28112 31580 28176 31584
rect 28112 31524 28116 31580
rect 28116 31524 28172 31580
rect 28172 31524 28176 31580
rect 28112 31520 28176 31524
rect 28192 31580 28256 31584
rect 28192 31524 28196 31580
rect 28196 31524 28252 31580
rect 28252 31524 28256 31580
rect 28192 31520 28256 31524
rect 37952 31580 38016 31584
rect 37952 31524 37956 31580
rect 37956 31524 38012 31580
rect 38012 31524 38016 31580
rect 37952 31520 38016 31524
rect 38032 31580 38096 31584
rect 38032 31524 38036 31580
rect 38036 31524 38092 31580
rect 38092 31524 38096 31580
rect 38032 31520 38096 31524
rect 38112 31580 38176 31584
rect 38112 31524 38116 31580
rect 38116 31524 38172 31580
rect 38172 31524 38176 31580
rect 38112 31520 38176 31524
rect 38192 31580 38256 31584
rect 38192 31524 38196 31580
rect 38196 31524 38252 31580
rect 38252 31524 38256 31580
rect 38192 31520 38256 31524
rect 47952 31580 48016 31584
rect 47952 31524 47956 31580
rect 47956 31524 48012 31580
rect 48012 31524 48016 31580
rect 47952 31520 48016 31524
rect 48032 31580 48096 31584
rect 48032 31524 48036 31580
rect 48036 31524 48092 31580
rect 48092 31524 48096 31580
rect 48032 31520 48096 31524
rect 48112 31580 48176 31584
rect 48112 31524 48116 31580
rect 48116 31524 48172 31580
rect 48172 31524 48176 31580
rect 48112 31520 48176 31524
rect 48192 31580 48256 31584
rect 48192 31524 48196 31580
rect 48196 31524 48252 31580
rect 48252 31524 48256 31580
rect 48192 31520 48256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 32952 31036 33016 31040
rect 32952 30980 32956 31036
rect 32956 30980 33012 31036
rect 33012 30980 33016 31036
rect 32952 30976 33016 30980
rect 33032 31036 33096 31040
rect 33032 30980 33036 31036
rect 33036 30980 33092 31036
rect 33092 30980 33096 31036
rect 33032 30976 33096 30980
rect 33112 31036 33176 31040
rect 33112 30980 33116 31036
rect 33116 30980 33172 31036
rect 33172 30980 33176 31036
rect 33112 30976 33176 30980
rect 33192 31036 33256 31040
rect 33192 30980 33196 31036
rect 33196 30980 33252 31036
rect 33252 30980 33256 31036
rect 33192 30976 33256 30980
rect 42952 31036 43016 31040
rect 42952 30980 42956 31036
rect 42956 30980 43012 31036
rect 43012 30980 43016 31036
rect 42952 30976 43016 30980
rect 43032 31036 43096 31040
rect 43032 30980 43036 31036
rect 43036 30980 43092 31036
rect 43092 30980 43096 31036
rect 43032 30976 43096 30980
rect 43112 31036 43176 31040
rect 43112 30980 43116 31036
rect 43116 30980 43172 31036
rect 43172 30980 43176 31036
rect 43112 30976 43176 30980
rect 43192 31036 43256 31040
rect 43192 30980 43196 31036
rect 43196 30980 43252 31036
rect 43252 30980 43256 31036
rect 43192 30976 43256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 27952 30492 28016 30496
rect 27952 30436 27956 30492
rect 27956 30436 28012 30492
rect 28012 30436 28016 30492
rect 27952 30432 28016 30436
rect 28032 30492 28096 30496
rect 28032 30436 28036 30492
rect 28036 30436 28092 30492
rect 28092 30436 28096 30492
rect 28032 30432 28096 30436
rect 28112 30492 28176 30496
rect 28112 30436 28116 30492
rect 28116 30436 28172 30492
rect 28172 30436 28176 30492
rect 28112 30432 28176 30436
rect 28192 30492 28256 30496
rect 28192 30436 28196 30492
rect 28196 30436 28252 30492
rect 28252 30436 28256 30492
rect 28192 30432 28256 30436
rect 37952 30492 38016 30496
rect 37952 30436 37956 30492
rect 37956 30436 38012 30492
rect 38012 30436 38016 30492
rect 37952 30432 38016 30436
rect 38032 30492 38096 30496
rect 38032 30436 38036 30492
rect 38036 30436 38092 30492
rect 38092 30436 38096 30492
rect 38032 30432 38096 30436
rect 38112 30492 38176 30496
rect 38112 30436 38116 30492
rect 38116 30436 38172 30492
rect 38172 30436 38176 30492
rect 38112 30432 38176 30436
rect 38192 30492 38256 30496
rect 38192 30436 38196 30492
rect 38196 30436 38252 30492
rect 38252 30436 38256 30492
rect 38192 30432 38256 30436
rect 47952 30492 48016 30496
rect 47952 30436 47956 30492
rect 47956 30436 48012 30492
rect 48012 30436 48016 30492
rect 47952 30432 48016 30436
rect 48032 30492 48096 30496
rect 48032 30436 48036 30492
rect 48036 30436 48092 30492
rect 48092 30436 48096 30492
rect 48032 30432 48096 30436
rect 48112 30492 48176 30496
rect 48112 30436 48116 30492
rect 48116 30436 48172 30492
rect 48172 30436 48176 30492
rect 48112 30432 48176 30436
rect 48192 30492 48256 30496
rect 48192 30436 48196 30492
rect 48196 30436 48252 30492
rect 48252 30436 48256 30492
rect 48192 30432 48256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 32952 29948 33016 29952
rect 32952 29892 32956 29948
rect 32956 29892 33012 29948
rect 33012 29892 33016 29948
rect 32952 29888 33016 29892
rect 33032 29948 33096 29952
rect 33032 29892 33036 29948
rect 33036 29892 33092 29948
rect 33092 29892 33096 29948
rect 33032 29888 33096 29892
rect 33112 29948 33176 29952
rect 33112 29892 33116 29948
rect 33116 29892 33172 29948
rect 33172 29892 33176 29948
rect 33112 29888 33176 29892
rect 33192 29948 33256 29952
rect 33192 29892 33196 29948
rect 33196 29892 33252 29948
rect 33252 29892 33256 29948
rect 33192 29888 33256 29892
rect 42952 29948 43016 29952
rect 42952 29892 42956 29948
rect 42956 29892 43012 29948
rect 43012 29892 43016 29948
rect 42952 29888 43016 29892
rect 43032 29948 43096 29952
rect 43032 29892 43036 29948
rect 43036 29892 43092 29948
rect 43092 29892 43096 29948
rect 43032 29888 43096 29892
rect 43112 29948 43176 29952
rect 43112 29892 43116 29948
rect 43116 29892 43172 29948
rect 43172 29892 43176 29948
rect 43112 29888 43176 29892
rect 43192 29948 43256 29952
rect 43192 29892 43196 29948
rect 43196 29892 43252 29948
rect 43252 29892 43256 29948
rect 43192 29888 43256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 27952 29404 28016 29408
rect 27952 29348 27956 29404
rect 27956 29348 28012 29404
rect 28012 29348 28016 29404
rect 27952 29344 28016 29348
rect 28032 29404 28096 29408
rect 28032 29348 28036 29404
rect 28036 29348 28092 29404
rect 28092 29348 28096 29404
rect 28032 29344 28096 29348
rect 28112 29404 28176 29408
rect 28112 29348 28116 29404
rect 28116 29348 28172 29404
rect 28172 29348 28176 29404
rect 28112 29344 28176 29348
rect 28192 29404 28256 29408
rect 28192 29348 28196 29404
rect 28196 29348 28252 29404
rect 28252 29348 28256 29404
rect 28192 29344 28256 29348
rect 37952 29404 38016 29408
rect 37952 29348 37956 29404
rect 37956 29348 38012 29404
rect 38012 29348 38016 29404
rect 37952 29344 38016 29348
rect 38032 29404 38096 29408
rect 38032 29348 38036 29404
rect 38036 29348 38092 29404
rect 38092 29348 38096 29404
rect 38032 29344 38096 29348
rect 38112 29404 38176 29408
rect 38112 29348 38116 29404
rect 38116 29348 38172 29404
rect 38172 29348 38176 29404
rect 38112 29344 38176 29348
rect 38192 29404 38256 29408
rect 38192 29348 38196 29404
rect 38196 29348 38252 29404
rect 38252 29348 38256 29404
rect 38192 29344 38256 29348
rect 47952 29404 48016 29408
rect 47952 29348 47956 29404
rect 47956 29348 48012 29404
rect 48012 29348 48016 29404
rect 47952 29344 48016 29348
rect 48032 29404 48096 29408
rect 48032 29348 48036 29404
rect 48036 29348 48092 29404
rect 48092 29348 48096 29404
rect 48032 29344 48096 29348
rect 48112 29404 48176 29408
rect 48112 29348 48116 29404
rect 48116 29348 48172 29404
rect 48172 29348 48176 29404
rect 48112 29344 48176 29348
rect 48192 29404 48256 29408
rect 48192 29348 48196 29404
rect 48196 29348 48252 29404
rect 48252 29348 48256 29404
rect 48192 29344 48256 29348
rect 35388 29004 35452 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 32952 28860 33016 28864
rect 32952 28804 32956 28860
rect 32956 28804 33012 28860
rect 33012 28804 33016 28860
rect 32952 28800 33016 28804
rect 33032 28860 33096 28864
rect 33032 28804 33036 28860
rect 33036 28804 33092 28860
rect 33092 28804 33096 28860
rect 33032 28800 33096 28804
rect 33112 28860 33176 28864
rect 33112 28804 33116 28860
rect 33116 28804 33172 28860
rect 33172 28804 33176 28860
rect 33112 28800 33176 28804
rect 33192 28860 33256 28864
rect 33192 28804 33196 28860
rect 33196 28804 33252 28860
rect 33252 28804 33256 28860
rect 33192 28800 33256 28804
rect 42952 28860 43016 28864
rect 42952 28804 42956 28860
rect 42956 28804 43012 28860
rect 43012 28804 43016 28860
rect 42952 28800 43016 28804
rect 43032 28860 43096 28864
rect 43032 28804 43036 28860
rect 43036 28804 43092 28860
rect 43092 28804 43096 28860
rect 43032 28800 43096 28804
rect 43112 28860 43176 28864
rect 43112 28804 43116 28860
rect 43116 28804 43172 28860
rect 43172 28804 43176 28860
rect 43112 28800 43176 28804
rect 43192 28860 43256 28864
rect 43192 28804 43196 28860
rect 43196 28804 43252 28860
rect 43252 28804 43256 28860
rect 43192 28800 43256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 27952 28316 28016 28320
rect 27952 28260 27956 28316
rect 27956 28260 28012 28316
rect 28012 28260 28016 28316
rect 27952 28256 28016 28260
rect 28032 28316 28096 28320
rect 28032 28260 28036 28316
rect 28036 28260 28092 28316
rect 28092 28260 28096 28316
rect 28032 28256 28096 28260
rect 28112 28316 28176 28320
rect 28112 28260 28116 28316
rect 28116 28260 28172 28316
rect 28172 28260 28176 28316
rect 28112 28256 28176 28260
rect 28192 28316 28256 28320
rect 28192 28260 28196 28316
rect 28196 28260 28252 28316
rect 28252 28260 28256 28316
rect 28192 28256 28256 28260
rect 37952 28316 38016 28320
rect 37952 28260 37956 28316
rect 37956 28260 38012 28316
rect 38012 28260 38016 28316
rect 37952 28256 38016 28260
rect 38032 28316 38096 28320
rect 38032 28260 38036 28316
rect 38036 28260 38092 28316
rect 38092 28260 38096 28316
rect 38032 28256 38096 28260
rect 38112 28316 38176 28320
rect 38112 28260 38116 28316
rect 38116 28260 38172 28316
rect 38172 28260 38176 28316
rect 38112 28256 38176 28260
rect 38192 28316 38256 28320
rect 38192 28260 38196 28316
rect 38196 28260 38252 28316
rect 38252 28260 38256 28316
rect 38192 28256 38256 28260
rect 47952 28316 48016 28320
rect 47952 28260 47956 28316
rect 47956 28260 48012 28316
rect 48012 28260 48016 28316
rect 47952 28256 48016 28260
rect 48032 28316 48096 28320
rect 48032 28260 48036 28316
rect 48036 28260 48092 28316
rect 48092 28260 48096 28316
rect 48032 28256 48096 28260
rect 48112 28316 48176 28320
rect 48112 28260 48116 28316
rect 48116 28260 48172 28316
rect 48172 28260 48176 28316
rect 48112 28256 48176 28260
rect 48192 28316 48256 28320
rect 48192 28260 48196 28316
rect 48196 28260 48252 28316
rect 48252 28260 48256 28316
rect 48192 28256 48256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 32952 27772 33016 27776
rect 32952 27716 32956 27772
rect 32956 27716 33012 27772
rect 33012 27716 33016 27772
rect 32952 27712 33016 27716
rect 33032 27772 33096 27776
rect 33032 27716 33036 27772
rect 33036 27716 33092 27772
rect 33092 27716 33096 27772
rect 33032 27712 33096 27716
rect 33112 27772 33176 27776
rect 33112 27716 33116 27772
rect 33116 27716 33172 27772
rect 33172 27716 33176 27772
rect 33112 27712 33176 27716
rect 33192 27772 33256 27776
rect 33192 27716 33196 27772
rect 33196 27716 33252 27772
rect 33252 27716 33256 27772
rect 33192 27712 33256 27716
rect 42952 27772 43016 27776
rect 42952 27716 42956 27772
rect 42956 27716 43012 27772
rect 43012 27716 43016 27772
rect 42952 27712 43016 27716
rect 43032 27772 43096 27776
rect 43032 27716 43036 27772
rect 43036 27716 43092 27772
rect 43092 27716 43096 27772
rect 43032 27712 43096 27716
rect 43112 27772 43176 27776
rect 43112 27716 43116 27772
rect 43116 27716 43172 27772
rect 43172 27716 43176 27772
rect 43112 27712 43176 27716
rect 43192 27772 43256 27776
rect 43192 27716 43196 27772
rect 43196 27716 43252 27772
rect 43252 27716 43256 27772
rect 43192 27712 43256 27716
rect 36124 27236 36188 27300
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 27952 27228 28016 27232
rect 27952 27172 27956 27228
rect 27956 27172 28012 27228
rect 28012 27172 28016 27228
rect 27952 27168 28016 27172
rect 28032 27228 28096 27232
rect 28032 27172 28036 27228
rect 28036 27172 28092 27228
rect 28092 27172 28096 27228
rect 28032 27168 28096 27172
rect 28112 27228 28176 27232
rect 28112 27172 28116 27228
rect 28116 27172 28172 27228
rect 28172 27172 28176 27228
rect 28112 27168 28176 27172
rect 28192 27228 28256 27232
rect 28192 27172 28196 27228
rect 28196 27172 28252 27228
rect 28252 27172 28256 27228
rect 28192 27168 28256 27172
rect 37952 27228 38016 27232
rect 37952 27172 37956 27228
rect 37956 27172 38012 27228
rect 38012 27172 38016 27228
rect 37952 27168 38016 27172
rect 38032 27228 38096 27232
rect 38032 27172 38036 27228
rect 38036 27172 38092 27228
rect 38092 27172 38096 27228
rect 38032 27168 38096 27172
rect 38112 27228 38176 27232
rect 38112 27172 38116 27228
rect 38116 27172 38172 27228
rect 38172 27172 38176 27228
rect 38112 27168 38176 27172
rect 38192 27228 38256 27232
rect 38192 27172 38196 27228
rect 38196 27172 38252 27228
rect 38252 27172 38256 27228
rect 38192 27168 38256 27172
rect 47952 27228 48016 27232
rect 47952 27172 47956 27228
rect 47956 27172 48012 27228
rect 48012 27172 48016 27228
rect 47952 27168 48016 27172
rect 48032 27228 48096 27232
rect 48032 27172 48036 27228
rect 48036 27172 48092 27228
rect 48092 27172 48096 27228
rect 48032 27168 48096 27172
rect 48112 27228 48176 27232
rect 48112 27172 48116 27228
rect 48116 27172 48172 27228
rect 48172 27172 48176 27228
rect 48112 27168 48176 27172
rect 48192 27228 48256 27232
rect 48192 27172 48196 27228
rect 48196 27172 48252 27228
rect 48252 27172 48256 27228
rect 48192 27168 48256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 32952 26684 33016 26688
rect 32952 26628 32956 26684
rect 32956 26628 33012 26684
rect 33012 26628 33016 26684
rect 32952 26624 33016 26628
rect 33032 26684 33096 26688
rect 33032 26628 33036 26684
rect 33036 26628 33092 26684
rect 33092 26628 33096 26684
rect 33032 26624 33096 26628
rect 33112 26684 33176 26688
rect 33112 26628 33116 26684
rect 33116 26628 33172 26684
rect 33172 26628 33176 26684
rect 33112 26624 33176 26628
rect 33192 26684 33256 26688
rect 33192 26628 33196 26684
rect 33196 26628 33252 26684
rect 33252 26628 33256 26684
rect 33192 26624 33256 26628
rect 42952 26684 43016 26688
rect 42952 26628 42956 26684
rect 42956 26628 43012 26684
rect 43012 26628 43016 26684
rect 42952 26624 43016 26628
rect 43032 26684 43096 26688
rect 43032 26628 43036 26684
rect 43036 26628 43092 26684
rect 43092 26628 43096 26684
rect 43032 26624 43096 26628
rect 43112 26684 43176 26688
rect 43112 26628 43116 26684
rect 43116 26628 43172 26684
rect 43172 26628 43176 26684
rect 43112 26624 43176 26628
rect 43192 26684 43256 26688
rect 43192 26628 43196 26684
rect 43196 26628 43252 26684
rect 43252 26628 43256 26684
rect 43192 26624 43256 26628
rect 35388 26284 35452 26348
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 27952 26140 28016 26144
rect 27952 26084 27956 26140
rect 27956 26084 28012 26140
rect 28012 26084 28016 26140
rect 27952 26080 28016 26084
rect 28032 26140 28096 26144
rect 28032 26084 28036 26140
rect 28036 26084 28092 26140
rect 28092 26084 28096 26140
rect 28032 26080 28096 26084
rect 28112 26140 28176 26144
rect 28112 26084 28116 26140
rect 28116 26084 28172 26140
rect 28172 26084 28176 26140
rect 28112 26080 28176 26084
rect 28192 26140 28256 26144
rect 28192 26084 28196 26140
rect 28196 26084 28252 26140
rect 28252 26084 28256 26140
rect 28192 26080 28256 26084
rect 37952 26140 38016 26144
rect 37952 26084 37956 26140
rect 37956 26084 38012 26140
rect 38012 26084 38016 26140
rect 37952 26080 38016 26084
rect 38032 26140 38096 26144
rect 38032 26084 38036 26140
rect 38036 26084 38092 26140
rect 38092 26084 38096 26140
rect 38032 26080 38096 26084
rect 38112 26140 38176 26144
rect 38112 26084 38116 26140
rect 38116 26084 38172 26140
rect 38172 26084 38176 26140
rect 38112 26080 38176 26084
rect 38192 26140 38256 26144
rect 38192 26084 38196 26140
rect 38196 26084 38252 26140
rect 38252 26084 38256 26140
rect 38192 26080 38256 26084
rect 47952 26140 48016 26144
rect 47952 26084 47956 26140
rect 47956 26084 48012 26140
rect 48012 26084 48016 26140
rect 47952 26080 48016 26084
rect 48032 26140 48096 26144
rect 48032 26084 48036 26140
rect 48036 26084 48092 26140
rect 48092 26084 48096 26140
rect 48032 26080 48096 26084
rect 48112 26140 48176 26144
rect 48112 26084 48116 26140
rect 48116 26084 48172 26140
rect 48172 26084 48176 26140
rect 48112 26080 48176 26084
rect 48192 26140 48256 26144
rect 48192 26084 48196 26140
rect 48196 26084 48252 26140
rect 48252 26084 48256 26140
rect 48192 26080 48256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 32952 25596 33016 25600
rect 32952 25540 32956 25596
rect 32956 25540 33012 25596
rect 33012 25540 33016 25596
rect 32952 25536 33016 25540
rect 33032 25596 33096 25600
rect 33032 25540 33036 25596
rect 33036 25540 33092 25596
rect 33092 25540 33096 25596
rect 33032 25536 33096 25540
rect 33112 25596 33176 25600
rect 33112 25540 33116 25596
rect 33116 25540 33172 25596
rect 33172 25540 33176 25596
rect 33112 25536 33176 25540
rect 33192 25596 33256 25600
rect 33192 25540 33196 25596
rect 33196 25540 33252 25596
rect 33252 25540 33256 25596
rect 33192 25536 33256 25540
rect 42952 25596 43016 25600
rect 42952 25540 42956 25596
rect 42956 25540 43012 25596
rect 43012 25540 43016 25596
rect 42952 25536 43016 25540
rect 43032 25596 43096 25600
rect 43032 25540 43036 25596
rect 43036 25540 43092 25596
rect 43092 25540 43096 25596
rect 43032 25536 43096 25540
rect 43112 25596 43176 25600
rect 43112 25540 43116 25596
rect 43116 25540 43172 25596
rect 43172 25540 43176 25596
rect 43112 25536 43176 25540
rect 43192 25596 43256 25600
rect 43192 25540 43196 25596
rect 43196 25540 43252 25596
rect 43252 25540 43256 25596
rect 43192 25536 43256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 27952 25052 28016 25056
rect 27952 24996 27956 25052
rect 27956 24996 28012 25052
rect 28012 24996 28016 25052
rect 27952 24992 28016 24996
rect 28032 25052 28096 25056
rect 28032 24996 28036 25052
rect 28036 24996 28092 25052
rect 28092 24996 28096 25052
rect 28032 24992 28096 24996
rect 28112 25052 28176 25056
rect 28112 24996 28116 25052
rect 28116 24996 28172 25052
rect 28172 24996 28176 25052
rect 28112 24992 28176 24996
rect 28192 25052 28256 25056
rect 28192 24996 28196 25052
rect 28196 24996 28252 25052
rect 28252 24996 28256 25052
rect 28192 24992 28256 24996
rect 37952 25052 38016 25056
rect 37952 24996 37956 25052
rect 37956 24996 38012 25052
rect 38012 24996 38016 25052
rect 37952 24992 38016 24996
rect 38032 25052 38096 25056
rect 38032 24996 38036 25052
rect 38036 24996 38092 25052
rect 38092 24996 38096 25052
rect 38032 24992 38096 24996
rect 38112 25052 38176 25056
rect 38112 24996 38116 25052
rect 38116 24996 38172 25052
rect 38172 24996 38176 25052
rect 38112 24992 38176 24996
rect 38192 25052 38256 25056
rect 38192 24996 38196 25052
rect 38196 24996 38252 25052
rect 38252 24996 38256 25052
rect 38192 24992 38256 24996
rect 47952 25052 48016 25056
rect 47952 24996 47956 25052
rect 47956 24996 48012 25052
rect 48012 24996 48016 25052
rect 47952 24992 48016 24996
rect 48032 25052 48096 25056
rect 48032 24996 48036 25052
rect 48036 24996 48092 25052
rect 48092 24996 48096 25052
rect 48032 24992 48096 24996
rect 48112 25052 48176 25056
rect 48112 24996 48116 25052
rect 48116 24996 48172 25052
rect 48172 24996 48176 25052
rect 48112 24992 48176 24996
rect 48192 25052 48256 25056
rect 48192 24996 48196 25052
rect 48196 24996 48252 25052
rect 48252 24996 48256 25052
rect 48192 24992 48256 24996
rect 31892 24984 31956 24988
rect 31892 24928 31906 24984
rect 31906 24928 31956 24984
rect 31892 24924 31956 24928
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 37596 23564 37660 23628
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 31892 17580 31956 17644
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 27660 14724 27724 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 32444 11052 32508 11116
rect 36124 11052 36188 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 35388 10644 35452 10708
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 26188 6700 26252 6764
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 37596 5068 37660 5132
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 28580 4116 28644 4180
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 32444 3572 32508 3636
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 27660 2348 27724 2412
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 27944 54432 28264 54448
rect 27944 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28264 54432
rect 27944 53344 28264 54368
rect 27944 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28264 53344
rect 27944 52256 28264 53280
rect 27944 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28264 52256
rect 27944 51168 28264 52192
rect 27944 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28264 51168
rect 27944 50080 28264 51104
rect 27944 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28264 50080
rect 27944 48992 28264 50016
rect 27944 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28264 48992
rect 27944 47904 28264 48928
rect 27944 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28264 47904
rect 27944 46816 28264 47840
rect 27944 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28264 46816
rect 27944 45728 28264 46752
rect 27944 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28264 45728
rect 27944 44640 28264 45664
rect 27944 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28264 44640
rect 27944 43552 28264 44576
rect 27944 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28264 43552
rect 27944 42464 28264 43488
rect 27944 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28264 42464
rect 27944 41376 28264 42400
rect 27944 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28264 41376
rect 27944 40288 28264 41312
rect 27944 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28264 40288
rect 27944 39200 28264 40224
rect 27944 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28264 39200
rect 27944 38112 28264 39136
rect 27944 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28264 38112
rect 27944 37024 28264 38048
rect 27944 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28264 37024
rect 27944 35936 28264 36960
rect 27944 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28264 35936
rect 27944 34848 28264 35872
rect 27944 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28264 34848
rect 27944 33760 28264 34784
rect 27944 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28264 33760
rect 26187 33692 26253 33693
rect 26187 33690 26188 33692
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 26006 33630 26188 33690
rect 26006 22110 26066 33630
rect 26187 33628 26188 33630
rect 26252 33628 26253 33692
rect 26187 33627 26253 33628
rect 27944 32672 28264 33696
rect 32944 53888 33264 54448
rect 32944 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33264 53888
rect 32944 52800 33264 53824
rect 32944 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33264 52800
rect 32944 51712 33264 52736
rect 32944 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33264 51712
rect 32944 50624 33264 51648
rect 32944 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33264 50624
rect 32944 49536 33264 50560
rect 32944 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33264 49536
rect 32944 48448 33264 49472
rect 32944 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33264 48448
rect 32944 47360 33264 48384
rect 32944 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33264 47360
rect 32944 46272 33264 47296
rect 32944 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33264 46272
rect 32944 45184 33264 46208
rect 32944 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33264 45184
rect 32944 44096 33264 45120
rect 32944 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33264 44096
rect 32944 43008 33264 44032
rect 32944 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33264 43008
rect 32944 41920 33264 42944
rect 32944 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33264 41920
rect 32944 40832 33264 41856
rect 32944 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33264 40832
rect 32944 39744 33264 40768
rect 32944 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33264 39744
rect 32944 38656 33264 39680
rect 32944 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33264 38656
rect 32944 37568 33264 38592
rect 32944 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33264 37568
rect 32944 36480 33264 37504
rect 32944 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33264 36480
rect 32944 35392 33264 36416
rect 32944 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33264 35392
rect 32944 34304 33264 35328
rect 32944 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33264 34304
rect 28579 33284 28645 33285
rect 28579 33220 28580 33284
rect 28644 33220 28645 33284
rect 28579 33219 28645 33220
rect 27944 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28264 32672
rect 27944 31584 28264 32608
rect 27944 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28264 31584
rect 27944 30496 28264 31520
rect 27944 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28264 30496
rect 27944 29408 28264 30432
rect 27944 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28264 29408
rect 27944 28320 28264 29344
rect 27944 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28264 28320
rect 27944 27232 28264 28256
rect 27944 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28264 27232
rect 27944 26144 28264 27168
rect 27944 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28264 26144
rect 27944 25056 28264 26080
rect 27944 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28264 25056
rect 27944 23968 28264 24992
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 26006 22050 26250 22110
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 26190 6765 26250 22050
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27659 14788 27725 14789
rect 27659 14724 27660 14788
rect 27724 14724 27725 14788
rect 27659 14723 27725 14724
rect 26187 6764 26253 6765
rect 26187 6700 26188 6764
rect 26252 6700 26253 6764
rect 26187 6699 26253 6700
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27662 2413 27722 14723
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 28582 4181 28642 33219
rect 32944 33216 33264 34240
rect 32944 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33264 33216
rect 32944 32128 33264 33152
rect 32944 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33264 32128
rect 32944 31040 33264 32064
rect 32944 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33264 31040
rect 32944 29952 33264 30976
rect 32944 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33264 29952
rect 32944 28864 33264 29888
rect 37944 54432 38264 54448
rect 37944 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38264 54432
rect 37944 53344 38264 54368
rect 37944 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38264 53344
rect 37944 52256 38264 53280
rect 37944 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38264 52256
rect 37944 51168 38264 52192
rect 37944 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38264 51168
rect 37944 50080 38264 51104
rect 37944 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38264 50080
rect 37944 48992 38264 50016
rect 37944 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38264 48992
rect 37944 47904 38264 48928
rect 37944 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38264 47904
rect 37944 46816 38264 47840
rect 37944 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38264 46816
rect 37944 45728 38264 46752
rect 37944 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38264 45728
rect 37944 44640 38264 45664
rect 37944 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38264 44640
rect 37944 43552 38264 44576
rect 37944 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38264 43552
rect 37944 42464 38264 43488
rect 37944 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38264 42464
rect 37944 41376 38264 42400
rect 37944 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38264 41376
rect 37944 40288 38264 41312
rect 37944 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38264 40288
rect 37944 39200 38264 40224
rect 37944 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38264 39200
rect 37944 38112 38264 39136
rect 37944 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38264 38112
rect 37944 37024 38264 38048
rect 37944 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38264 37024
rect 37944 35936 38264 36960
rect 37944 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38264 35936
rect 37944 34848 38264 35872
rect 37944 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38264 34848
rect 37944 33760 38264 34784
rect 37944 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38264 33760
rect 37944 32672 38264 33696
rect 37944 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38264 32672
rect 37944 31584 38264 32608
rect 37944 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38264 31584
rect 37944 30496 38264 31520
rect 37944 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38264 30496
rect 37944 29408 38264 30432
rect 37944 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38264 29408
rect 35387 29068 35453 29069
rect 35387 29004 35388 29068
rect 35452 29004 35453 29068
rect 35387 29003 35453 29004
rect 32944 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33264 28864
rect 32944 27776 33264 28800
rect 32944 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33264 27776
rect 32944 26688 33264 27712
rect 32944 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33264 26688
rect 32944 25600 33264 26624
rect 35390 26349 35450 29003
rect 37944 28320 38264 29344
rect 37944 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38264 28320
rect 36123 27300 36189 27301
rect 36123 27236 36124 27300
rect 36188 27236 36189 27300
rect 36123 27235 36189 27236
rect 35387 26348 35453 26349
rect 35387 26284 35388 26348
rect 35452 26284 35453 26348
rect 35387 26283 35453 26284
rect 32944 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33264 25600
rect 31891 24988 31957 24989
rect 31891 24924 31892 24988
rect 31956 24924 31957 24988
rect 31891 24923 31957 24924
rect 31894 17645 31954 24923
rect 32944 24512 33264 25536
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 31891 17644 31957 17645
rect 31891 17580 31892 17644
rect 31956 17580 31957 17644
rect 31891 17579 31957 17580
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32443 11116 32509 11117
rect 32443 11052 32444 11116
rect 32508 11052 32509 11116
rect 32443 11051 32509 11052
rect 28579 4180 28645 4181
rect 28579 4116 28580 4180
rect 28644 4116 28645 4180
rect 28579 4115 28645 4116
rect 32446 3637 32506 11051
rect 32944 10368 33264 11392
rect 35390 10709 35450 26283
rect 36126 11117 36186 27235
rect 37944 27232 38264 28256
rect 37944 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38264 27232
rect 37944 26144 38264 27168
rect 37944 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38264 26144
rect 37944 25056 38264 26080
rect 37944 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38264 25056
rect 37944 23968 38264 24992
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37595 23628 37661 23629
rect 37595 23564 37596 23628
rect 37660 23564 37661 23628
rect 37595 23563 37661 23564
rect 36123 11116 36189 11117
rect 36123 11052 36124 11116
rect 36188 11052 36189 11116
rect 36123 11051 36189 11052
rect 35387 10708 35453 10709
rect 35387 10644 35388 10708
rect 35452 10644 35453 10708
rect 35387 10643 35453 10644
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 37598 5133 37658 23563
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37595 5132 37661 5133
rect 37595 5068 37596 5132
rect 37660 5068 37661 5132
rect 37595 5067 37661 5068
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32443 3636 32509 3637
rect 32443 3572 32444 3636
rect 32508 3572 32509 3636
rect 32443 3571 32509 3572
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27659 2412 27725 2413
rect 27659 2348 27660 2412
rect 27724 2348 27725 2412
rect 27659 2347 27725 2348
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 53888 43264 54448
rect 42944 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43264 53888
rect 42944 52800 43264 53824
rect 42944 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43264 52800
rect 42944 51712 43264 52736
rect 42944 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43264 51712
rect 42944 50624 43264 51648
rect 42944 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43264 50624
rect 42944 49536 43264 50560
rect 42944 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43264 49536
rect 42944 48448 43264 49472
rect 42944 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43264 48448
rect 42944 47360 43264 48384
rect 42944 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43264 47360
rect 42944 46272 43264 47296
rect 42944 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43264 46272
rect 42944 45184 43264 46208
rect 42944 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43264 45184
rect 42944 44096 43264 45120
rect 42944 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43264 44096
rect 42944 43008 43264 44032
rect 42944 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43264 43008
rect 42944 41920 43264 42944
rect 42944 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43264 41920
rect 42944 40832 43264 41856
rect 42944 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43264 40832
rect 42944 39744 43264 40768
rect 42944 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43264 39744
rect 42944 38656 43264 39680
rect 42944 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43264 38656
rect 42944 37568 43264 38592
rect 42944 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43264 37568
rect 42944 36480 43264 37504
rect 42944 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43264 36480
rect 42944 35392 43264 36416
rect 42944 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43264 35392
rect 42944 34304 43264 35328
rect 42944 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43264 34304
rect 42944 33216 43264 34240
rect 42944 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43264 33216
rect 42944 32128 43264 33152
rect 42944 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43264 32128
rect 42944 31040 43264 32064
rect 42944 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43264 31040
rect 42944 29952 43264 30976
rect 42944 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43264 29952
rect 42944 28864 43264 29888
rect 42944 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43264 28864
rect 42944 27776 43264 28800
rect 42944 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43264 27776
rect 42944 26688 43264 27712
rect 42944 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43264 26688
rect 42944 25600 43264 26624
rect 42944 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43264 25600
rect 42944 24512 43264 25536
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 54432 48264 54448
rect 47944 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48264 54432
rect 47944 53344 48264 54368
rect 47944 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48264 53344
rect 47944 52256 48264 53280
rect 47944 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48264 52256
rect 47944 51168 48264 52192
rect 47944 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48264 51168
rect 47944 50080 48264 51104
rect 47944 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48264 50080
rect 47944 48992 48264 50016
rect 47944 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48264 48992
rect 47944 47904 48264 48928
rect 47944 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48264 47904
rect 47944 46816 48264 47840
rect 47944 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48264 46816
rect 47944 45728 48264 46752
rect 47944 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48264 45728
rect 47944 44640 48264 45664
rect 47944 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48264 44640
rect 47944 43552 48264 44576
rect 47944 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48264 43552
rect 47944 42464 48264 43488
rect 47944 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48264 42464
rect 47944 41376 48264 42400
rect 47944 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48264 41376
rect 47944 40288 48264 41312
rect 47944 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48264 40288
rect 47944 39200 48264 40224
rect 47944 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48264 39200
rect 47944 38112 48264 39136
rect 47944 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48264 38112
rect 47944 37024 48264 38048
rect 47944 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48264 37024
rect 47944 35936 48264 36960
rect 47944 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48264 35936
rect 47944 34848 48264 35872
rect 47944 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48264 34848
rect 47944 33760 48264 34784
rect 47944 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48264 33760
rect 47944 32672 48264 33696
rect 47944 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48264 32672
rect 47944 31584 48264 32608
rect 47944 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48264 31584
rect 47944 30496 48264 31520
rect 47944 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48264 30496
rect 47944 29408 48264 30432
rect 47944 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48264 29408
rect 47944 28320 48264 29344
rect 47944 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48264 28320
rect 47944 27232 48264 28256
rect 47944 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48264 27232
rect 47944 26144 48264 27168
rect 47944 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48264 26144
rect 47944 25056 48264 26080
rect 47944 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48264 25056
rect 47944 23968 48264 24992
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_1  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1676037725
transform 1 0 46000 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1676037725
transform 1 0 46276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _107_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 46736 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1676037725
transform 1 0 46920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 46552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 46736 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 46000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1676037725
transform 1 0 46276 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1676037725
transform 1 0 46644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform 1 0 45908 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 45172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 44528 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 45632 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 45816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 45448 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1676037725
transform 1 0 45632 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 44160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 43240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 44160 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1676037725
transform 1 0 44988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 44896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1676037725
transform 1 0 45172 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 43792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform 1 0 42780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 45172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 45908 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1676037725
transform 1 0 46368 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 43884 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1676037725
transform 1 0 43424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 37628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 29716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 28520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 32292 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 33120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 34868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 35604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 35236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 35972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 36064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 36616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 32384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 34868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 39008 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 38548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 44068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 45172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 35696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 38088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 39376 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 40020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 40756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 40756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 39836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _165_
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 14812 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1676037725
transform 1 0 17020 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 19412 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 20792 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 22816 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 43792 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 43332 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 40388 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 42688 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 31556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 30452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 30268 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 27324 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 32292 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 30360 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 22172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 25852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 22172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 36064 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 33672 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 36064 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 34500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 34040 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 33856 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 28244 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 26680 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 27600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 31004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11408 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23736 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25300 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24104 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 23368 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 27416 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 26128 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29256 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29532 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 30452 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 30360 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27416 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__194 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 25852 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 25576 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 23552 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22908 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 31924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 30912 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 31556 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 28796 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28796 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__195
timestamp 1676037725
transform 1 0 28428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 28336 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 26588 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 24932 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22264 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 30728 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 28152 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 29072 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28428 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 25116 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__196
timestamp 1676037725
transform 1 0 34040 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 32844 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 28612 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 25944 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29900 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28336 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 27232 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 27876 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27784 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 26680 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 23368 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__197
timestamp 1676037725
transform 1 0 32292 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 30912 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 25576 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 23644 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20240 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29532 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22356 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 27324 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 21160 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 20792 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21528 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 25668 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22264 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 19320 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 23184 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 20240 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 17112 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14352 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31372 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25668 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 27416 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 27324 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 29900 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 33396 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 36248 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 34868 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 37260 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 32476 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 32752 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 35420 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 41124 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 43240 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 41952 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 42780 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1676037725
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120
timestamp 1676037725
transform 1 0 12144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1676037725
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1676037725
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_217
timestamp 1676037725
transform 1 0 21068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_236
timestamp 1676037725
transform 1 0 22816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1676037725
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1676037725
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1676037725
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1676037725
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1676037725
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_467
timestamp 1676037725
transform 1 0 44068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_495
timestamp 1676037725
transform 1 0 46644 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1676037725
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_523
timestamp 1676037725
transform 1 0 49220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_23
timestamp 1676037725
transform 1 0 3220 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1676037725
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp 1676037725
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1676037725
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_64
timestamp 1676037725
transform 1 0 6992 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_76
timestamp 1676037725
transform 1 0 8096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_84
timestamp 1676037725
transform 1 0 8832 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1676037725
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_118
timestamp 1676037725
transform 1 0 11960 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_124
timestamp 1676037725
transform 1 0 12512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_135
timestamp 1676037725
transform 1 0 13524 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_151
timestamp 1676037725
transform 1 0 14996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1676037725
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_191
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_251
timestamp 1676037725
transform 1 0 24196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_259
timestamp 1676037725
transform 1 0 24932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1676037725
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1676037725
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_321
timestamp 1676037725
transform 1 0 30636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1676037725
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_355
timestamp 1676037725
transform 1 0 33764 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_375
timestamp 1676037725
transform 1 0 35604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1676037725
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_411
timestamp 1676037725
transform 1 0 38916 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_431
timestamp 1676037725
transform 1 0 40756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1676037725
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_467
timestamp 1676037725
transform 1 0 44068 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_487
timestamp 1676037725
transform 1 0 45908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_499
timestamp 1676037725
transform 1 0 47012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_176
timestamp 1676037725
transform 1 0 17296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1676037725
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_227
timestamp 1676037725
transform 1 0 21988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_239
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_271
timestamp 1676037725
transform 1 0 26036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_283
timestamp 1676037725
transform 1 0 27140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_295
timestamp 1676037725
transform 1 0 28244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_327
timestamp 1676037725
transform 1 0 31188 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_347
timestamp 1676037725
transform 1 0 33028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1676037725
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1676037725
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1676037725
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1676037725
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_439
timestamp 1676037725
transform 1 0 41492 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_459
timestamp 1676037725
transform 1 0 43332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_471
timestamp 1676037725
transform 1 0 44436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_495
timestamp 1676037725
transform 1 0 46644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_521
timestamp 1676037725
transform 1 0 49036 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_494
timestamp 1676037725
transform 1 0 46552 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1676037725
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1676037725
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1676037725
transform 1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_425
timestamp 1676037725
transform 1 0 40204 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_435
timestamp 1676037725
transform 1 0 41124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_491
timestamp 1676037725
transform 1 0 46276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_315
timestamp 1676037725
transform 1 0 30084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_327
timestamp 1676037725
transform 1 0 31188 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_335
timestamp 1676037725
transform 1 0 31924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_406
timestamp 1676037725
transform 1 0 38456 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_414
timestamp 1676037725
transform 1 0 39192 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_427
timestamp 1676037725
transform 1 0 40388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_435
timestamp 1676037725
transform 1 0 41124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_443
timestamp 1676037725
transform 1 0 41860 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_448
timestamp 1676037725
transform 1 0 42320 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_460
timestamp 1676037725
transform 1 0 43424 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_472
timestamp 1676037725
transform 1 0 44528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_482
timestamp 1676037725
transform 1 0 45448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_494
timestamp 1676037725
transform 1 0 46552 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_500
timestamp 1676037725
transform 1 0 47104 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_508
timestamp 1676037725
transform 1 0 47840 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_359
timestamp 1676037725
transform 1 0 34132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_371
timestamp 1676037725
transform 1 0 35236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_383
timestamp 1676037725
transform 1 0 36340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_399
timestamp 1676037725
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_407
timestamp 1676037725
transform 1 0 38548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_415
timestamp 1676037725
transform 1 0 39284 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_420
timestamp 1676037725
transform 1 0 39744 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_432
timestamp 1676037725
transform 1 0 40848 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_444
timestamp 1676037725
transform 1 0 41952 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_331
timestamp 1676037725
transform 1 0 31556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1676037725
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_371
timestamp 1676037725
transform 1 0 35236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_375
timestamp 1676037725
transform 1 0 35604 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_380
timestamp 1676037725
transform 1 0 36064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_404
timestamp 1676037725
transform 1 0 38272 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_417
timestamp 1676037725
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_442
timestamp 1676037725
transform 1 0 41768 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_454
timestamp 1676037725
transform 1 0 42872 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_466
timestamp 1676037725
transform 1 0 43976 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_474
timestamp 1676037725
transform 1 0 44712 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_297
timestamp 1676037725
transform 1 0 28428 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_302
timestamp 1676037725
transform 1 0 28888 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_314
timestamp 1676037725
transform 1 0 29992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_326
timestamp 1676037725
transform 1 0 31096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1676037725
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_344
timestamp 1676037725
transform 1 0 32752 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_368
timestamp 1676037725
transform 1 0 34960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_381
timestamp 1676037725
transform 1 0 36156 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1676037725
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_401
timestamp 1676037725
transform 1 0 37996 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_407
timestamp 1676037725
transform 1 0 38548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_419
timestamp 1676037725
transform 1 0 39652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_431
timestamp 1676037725
transform 1 0 40756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_443
timestamp 1676037725
transform 1 0 41860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_455
timestamp 1676037725
transform 1 0 42964 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_459
timestamp 1676037725
transform 1 0 43332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_471
timestamp 1676037725
transform 1 0 44436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_483
timestamp 1676037725
transform 1 0 45540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_495
timestamp 1676037725
transform 1 0 46644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1676037725
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_291
timestamp 1676037725
transform 1 0 27876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1676037725
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_340
timestamp 1676037725
transform 1 0 32384 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_347
timestamp 1676037725
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_359
timestamp 1676037725
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_372
timestamp 1676037725
transform 1 0 35328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_376
timestamp 1676037725
transform 1 0 35696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_397
timestamp 1676037725
transform 1 0 37628 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_408
timestamp 1676037725
transform 1 0 38640 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_426
timestamp 1676037725
transform 1 0 40296 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_438
timestamp 1676037725
transform 1 0 41400 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_450
timestamp 1676037725
transform 1 0 42504 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_462
timestamp 1676037725
transform 1 0 43608 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_474
timestamp 1676037725
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1676037725
transform 1 0 23092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_252
timestamp 1676037725
transform 1 0 24288 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_265
timestamp 1676037725
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_287
timestamp 1676037725
transform 1 0 27508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_308
timestamp 1676037725
transform 1 0 29440 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_320
timestamp 1676037725
transform 1 0 30544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1676037725
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_348
timestamp 1676037725
transform 1 0 33120 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_356
timestamp 1676037725
transform 1 0 33856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_378
timestamp 1676037725
transform 1 0 35880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1676037725
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_397
timestamp 1676037725
transform 1 0 37628 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_418
timestamp 1676037725
transform 1 0 39560 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_431
timestamp 1676037725
transform 1 0 40756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_443
timestamp 1676037725
transform 1 0 41860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_493
timestamp 1676037725
transform 1 0 46460 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_498
timestamp 1676037725
transform 1 0 46920 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1676037725
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1676037725
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_261
timestamp 1676037725
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_283
timestamp 1676037725
transform 1 0 27140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_295
timestamp 1676037725
transform 1 0 28244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_331
timestamp 1676037725
transform 1 0 31556 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_344
timestamp 1676037725
transform 1 0 32752 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_352
timestamp 1676037725
transform 1 0 33488 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_387
timestamp 1676037725
transform 1 0 36708 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_400
timestamp 1676037725
transform 1 0 37904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_426
timestamp 1676037725
transform 1 0 40296 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_434
timestamp 1676037725
transform 1 0 41032 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_439
timestamp 1676037725
transform 1 0 41492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_451
timestamp 1676037725
transform 1 0 42596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_463
timestamp 1676037725
transform 1 0 43700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_483
timestamp 1676037725
transform 1 0 45540 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_490
timestamp 1676037725
transform 1 0 46184 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_494
timestamp 1676037725
transform 1 0 46552 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_498
timestamp 1676037725
transform 1 0 46920 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_506
timestamp 1676037725
transform 1 0 47656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_242
timestamp 1676037725
transform 1 0 23368 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_254
timestamp 1676037725
transform 1 0 24472 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_266
timestamp 1676037725
transform 1 0 25576 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_272
timestamp 1676037725
transform 1 0 26128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1676037725
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_302
timestamp 1676037725
transform 1 0 28888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_315
timestamp 1676037725
transform 1 0 30084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_328
timestamp 1676037725
transform 1 0 31280 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_343
timestamp 1676037725
transform 1 0 32660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_353
timestamp 1676037725
transform 1 0 33580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_379
timestamp 1676037725
transform 1 0 35972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_384
timestamp 1676037725
transform 1 0 36432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_398
timestamp 1676037725
transform 1 0 37720 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_426
timestamp 1676037725
transform 1 0 40296 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_438
timestamp 1676037725
transform 1 0 41400 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_446
timestamp 1676037725
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_464
timestamp 1676037725
transform 1 0 43792 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_476
timestamp 1676037725
transform 1 0 44896 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_488
timestamp 1676037725
transform 1 0 46000 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_494
timestamp 1676037725
transform 1 0 46552 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_502
timestamp 1676037725
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_288
timestamp 1676037725
transform 1 0 27600 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_300
timestamp 1676037725
transform 1 0 28704 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_341
timestamp 1676037725
transform 1 0 32476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_354
timestamp 1676037725
transform 1 0 33672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1676037725
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_371
timestamp 1676037725
transform 1 0 35236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_392
timestamp 1676037725
transform 1 0 37168 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_399
timestamp 1676037725
transform 1 0 37812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_410
timestamp 1676037725
transform 1 0 38824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_418
timestamp 1676037725
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_485
timestamp 1676037725
transform 1 0 45724 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_492
timestamp 1676037725
transform 1 0 46368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_500
timestamp 1676037725
transform 1 0 47104 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_508
timestamp 1676037725
transform 1 0 47840 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_318
timestamp 1676037725
transform 1 0 30360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_331
timestamp 1676037725
transform 1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_343
timestamp 1676037725
transform 1 0 32660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_347
timestamp 1676037725
transform 1 0 33028 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_369
timestamp 1676037725
transform 1 0 35052 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 1676037725
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_431
timestamp 1676037725
transform 1 0 40756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_443
timestamp 1676037725
transform 1 0 41860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_454
timestamp 1676037725
transform 1 0 42872 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_466
timestamp 1676037725
transform 1 0 43976 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_478
timestamp 1676037725
transform 1 0 45080 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_490
timestamp 1676037725
transform 1 0 46184 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_502
timestamp 1676037725
transform 1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_261
timestamp 1676037725
transform 1 0 25116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_284
timestamp 1676037725
transform 1 0 27232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_290
timestamp 1676037725
transform 1 0 27784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1676037725
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_320
timestamp 1676037725
transform 1 0 30544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_333
timestamp 1676037725
transform 1 0 31740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_346
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_350
timestamp 1676037725
transform 1 0 33304 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_376
timestamp 1676037725
transform 1 0 35696 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_393
timestamp 1676037725
transform 1 0 37260 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_400
timestamp 1676037725
transform 1 0 37904 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1676037725
transform 1 0 38456 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_411
timestamp 1676037725
transform 1 0 38916 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1676037725
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_245
timestamp 1676037725
transform 1 0 23644 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_267
timestamp 1676037725
transform 1 0 25668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1676037725
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_322
timestamp 1676037725
transform 1 0 30728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1676037725
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_376
timestamp 1676037725
transform 1 0 35696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_383
timestamp 1676037725
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_408
timestamp 1676037725
transform 1 0 38640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_416
timestamp 1676037725
transform 1 0 39376 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_433
timestamp 1676037725
transform 1 0 40940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_440
timestamp 1676037725
transform 1 0 41584 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_454
timestamp 1676037725
transform 1 0 42872 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_466
timestamp 1676037725
transform 1 0 43976 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_475
timestamp 1676037725
transform 1 0 44804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_487
timestamp 1676037725
transform 1 0 45908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_499
timestamp 1676037725
transform 1 0 47012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_264
timestamp 1676037725
transform 1 0 25392 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_276
timestamp 1676037725
transform 1 0 26496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 1676037725
transform 1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_293
timestamp 1676037725
transform 1 0 28060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1676037725
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_320
timestamp 1676037725
transform 1 0 30544 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_332
timestamp 1676037725
transform 1 0 31648 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_344
timestamp 1676037725
transform 1 0 32752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_376
timestamp 1676037725
transform 1 0 35696 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1676037725
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_409
timestamp 1676037725
transform 1 0 38732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1676037725
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_426
timestamp 1676037725
transform 1 0 40296 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_438
timestamp 1676037725
transform 1 0 41400 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_450
timestamp 1676037725
transform 1 0 42504 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_462
timestamp 1676037725
transform 1 0 43608 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1676037725
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_246
timestamp 1676037725
transform 1 0 23736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1676037725
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1676037725
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_295
timestamp 1676037725
transform 1 0 28244 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_310
timestamp 1676037725
transform 1 0 29624 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_348
timestamp 1676037725
transform 1 0 33120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_355
timestamp 1676037725
transform 1 0 33764 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_363
timestamp 1676037725
transform 1 0 34500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_367
timestamp 1676037725
transform 1 0 34868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_375
timestamp 1676037725
transform 1 0 35604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_383
timestamp 1676037725
transform 1 0 36340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1676037725
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_399
timestamp 1676037725
transform 1 0 37812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_411
timestamp 1676037725
transform 1 0 38916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_434
timestamp 1676037725
transform 1 0 41032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_438
timestamp 1676037725
transform 1 0 41400 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_442
timestamp 1676037725
transform 1 0 41768 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1676037725
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1676037725
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1676037725
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_211
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_225
timestamp 1676037725
transform 1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_234
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_268
timestamp 1676037725
transform 1 0 25760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1676037725
transform 1 0 26496 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_286
timestamp 1676037725
transform 1 0 27416 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1676037725
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_317
timestamp 1676037725
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_327
timestamp 1676037725
transform 1 0 31188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_342
timestamp 1676037725
transform 1 0 32568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_353
timestamp 1676037725
transform 1 0 33580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1676037725
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_371
timestamp 1676037725
transform 1 0 35236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_379
timestamp 1676037725
transform 1 0 35972 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_383
timestamp 1676037725
transform 1 0 36340 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_404
timestamp 1676037725
transform 1 0 38272 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_412
timestamp 1676037725
transform 1 0 39008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_418
timestamp 1676037725
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_426
timestamp 1676037725
transform 1 0 40296 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_438
timestamp 1676037725
transform 1 0 41400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_446
timestamp 1676037725
transform 1 0 42136 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_450
timestamp 1676037725
transform 1 0 42504 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_462
timestamp 1676037725
transform 1 0 43608 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_472
timestamp 1676037725
transform 1 0 44528 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_209
timestamp 1676037725
transform 1 0 20332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1676037725
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_233
timestamp 1676037725
transform 1 0 22540 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_268
timestamp 1676037725
transform 1 0 25760 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_309
timestamp 1676037725
transform 1 0 29532 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_326
timestamp 1676037725
transform 1 0 31096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_330
timestamp 1676037725
transform 1 0 31464 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_365
timestamp 1676037725
transform 1 0 34684 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_378
timestamp 1676037725
transform 1 0 35880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_404
timestamp 1676037725
transform 1 0 38272 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_432
timestamp 1676037725
transform 1 0 40848 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_444
timestamp 1676037725
transform 1 0 41952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_457
timestamp 1676037725
transform 1 0 43148 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_462
timestamp 1676037725
transform 1 0 43608 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_474
timestamp 1676037725
transform 1 0 44712 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_482
timestamp 1676037725
transform 1 0 45448 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_488
timestamp 1676037725
transform 1 0 46000 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_500
timestamp 1676037725
transform 1 0 47104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1676037725
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_262
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_275
timestamp 1676037725
transform 1 0 26404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_317
timestamp 1676037725
transform 1 0 30268 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_327
timestamp 1676037725
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_340
timestamp 1676037725
transform 1 0 32384 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_352
timestamp 1676037725
transform 1 0 33488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_369
timestamp 1676037725
transform 1 0 35052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_379
timestamp 1676037725
transform 1 0 35972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_386
timestamp 1676037725
transform 1 0 36616 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_392
timestamp 1676037725
transform 1 0 37168 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_404
timestamp 1676037725
transform 1 0 38272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_408
timestamp 1676037725
transform 1 0 38640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_430
timestamp 1676037725
transform 1 0 40664 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_437
timestamp 1676037725
transform 1 0 41308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_449
timestamp 1676037725
transform 1 0 42412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_461
timestamp 1676037725
transform 1 0 43516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1676037725
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_483
timestamp 1676037725
transform 1 0 45540 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_487
timestamp 1676037725
transform 1 0 45908 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_499
timestamp 1676037725
transform 1 0 47012 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_511
timestamp 1676037725
transform 1 0 48116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_523
timestamp 1676037725
transform 1 0 49220 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_241
timestamp 1676037725
transform 1 0 23276 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_262
timestamp 1676037725
transform 1 0 25208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_266
timestamp 1676037725
transform 1 0 25576 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_291
timestamp 1676037725
transform 1 0 27876 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_297
timestamp 1676037725
transform 1 0 28428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_310
timestamp 1676037725
transform 1 0 29624 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_314
timestamp 1676037725
transform 1 0 29992 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_324
timestamp 1676037725
transform 1 0 30912 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_359
timestamp 1676037725
transform 1 0 34132 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_378
timestamp 1676037725
transform 1 0 35880 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_386
timestamp 1676037725
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_400
timestamp 1676037725
transform 1 0 37904 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_408
timestamp 1676037725
transform 1 0 38640 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1676037725
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_489
timestamp 1676037725
transform 1 0 46092 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_501
timestamp 1676037725
transform 1 0 47196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_285
timestamp 1676037725
transform 1 0 27324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1676037725
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_317
timestamp 1676037725
transform 1 0 30268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_322
timestamp 1676037725
transform 1 0 30728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_335
timestamp 1676037725
transform 1 0 31924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_342
timestamp 1676037725
transform 1 0 32568 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_350
timestamp 1676037725
transform 1 0 33304 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1676037725
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_373
timestamp 1676037725
transform 1 0 35420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_395
timestamp 1676037725
transform 1 0 37444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_408
timestamp 1676037725
transform 1 0 38640 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1676037725
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_465
timestamp 1676037725
transform 1 0 43884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_472
timestamp 1676037725
transform 1 0 44528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_481
timestamp 1676037725
transform 1 0 45356 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_486
timestamp 1676037725
transform 1 0 45816 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_498
timestamp 1676037725
transform 1 0 46920 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_506
timestamp 1676037725
transform 1 0 47656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_253
timestamp 1676037725
transform 1 0 24380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1676037725
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_316
timestamp 1676037725
transform 1 0 30176 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_328
timestamp 1676037725
transform 1 0 31280 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1676037725
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_372
timestamp 1676037725
transform 1 0 35328 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1676037725
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_398
timestamp 1676037725
transform 1 0 37720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_406
timestamp 1676037725
transform 1 0 38456 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_412
timestamp 1676037725
transform 1 0 39008 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_424
timestamp 1676037725
transform 1 0 40112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_428
timestamp 1676037725
transform 1 0 40480 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_432
timestamp 1676037725
transform 1 0 40848 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_444
timestamp 1676037725
transform 1 0 41952 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1676037725
transform 1 0 20700 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_217
timestamp 1676037725
transform 1 0 21068 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_229
timestamp 1676037725
transform 1 0 22172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_270
timestamp 1676037725
transform 1 0 25944 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_287
timestamp 1676037725
transform 1 0 27508 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_293
timestamp 1676037725
transform 1 0 28060 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1676037725
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_331
timestamp 1676037725
transform 1 0 31556 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_355
timestamp 1676037725
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_371
timestamp 1676037725
transform 1 0 35236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_375
timestamp 1676037725
transform 1 0 35604 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_381
timestamp 1676037725
transform 1 0 36156 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_386
timestamp 1676037725
transform 1 0 36616 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_398
timestamp 1676037725
transform 1 0 37720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_410
timestamp 1676037725
transform 1 0 38824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1676037725
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_426
timestamp 1676037725
transform 1 0 40296 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_438
timestamp 1676037725
transform 1 0 41400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_446
timestamp 1676037725
transform 1 0 42136 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_456
timestamp 1676037725
transform 1 0 43056 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_468
timestamp 1676037725
transform 1 0 44160 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1676037725
transform 1 0 19596 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_249
timestamp 1676037725
transform 1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_257
timestamp 1676037725
transform 1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1676037725
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1676037725
transform 1 0 27508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_300
timestamp 1676037725
transform 1 0 28704 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_313
timestamp 1676037725
transform 1 0 29900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_328
timestamp 1676037725
transform 1 0 31280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_343
timestamp 1676037725
transform 1 0 32660 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_356
timestamp 1676037725
transform 1 0 33856 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_368
timestamp 1676037725
transform 1 0 34960 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_380
timestamp 1676037725
transform 1 0 36064 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_415
timestamp 1676037725
transform 1 0 39284 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_439
timestamp 1676037725
transform 1 0 41492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1676037725
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_460
timestamp 1676037725
transform 1 0 43424 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_487
timestamp 1676037725
transform 1 0 45908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_499
timestamp 1676037725
transform 1 0 47012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1676037725
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_261
timestamp 1676037725
transform 1 0 25116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_287
timestamp 1676037725
transform 1 0 27508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_300
timestamp 1676037725
transform 1 0 28704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_314
timestamp 1676037725
transform 1 0 29992 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_326
timestamp 1676037725
transform 1 0 31096 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_338
timestamp 1676037725
transform 1 0 32200 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_350
timestamp 1676037725
transform 1 0 33304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_355
timestamp 1676037725
transform 1 0 33764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1676037725
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_393
timestamp 1676037725
transform 1 0 37260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_405
timestamp 1676037725
transform 1 0 38364 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_413
timestamp 1676037725
transform 1 0 39100 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_417
timestamp 1676037725
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_425
timestamp 1676037725
transform 1 0 40204 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_429
timestamp 1676037725
transform 1 0 40572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_437
timestamp 1676037725
transform 1 0 41308 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_449
timestamp 1676037725
transform 1 0 42412 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_455
timestamp 1676037725
transform 1 0 42964 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_471
timestamp 1676037725
transform 1 0 44436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1676037725
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_483
timestamp 1676037725
transform 1 0 45540 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_495
timestamp 1676037725
transform 1 0 46644 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_507
timestamp 1676037725
transform 1 0 47748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_519
timestamp 1676037725
transform 1 0 48852 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_241
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_251
timestamp 1676037725
transform 1 0 24196 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_263
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_267
timestamp 1676037725
transform 1 0 25668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1676037725
transform 1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1676037725
transform 1 0 28520 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_308
timestamp 1676037725
transform 1 0 29440 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1676037725
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_365
timestamp 1676037725
transform 1 0 34684 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_378
timestamp 1676037725
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1676037725
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_415
timestamp 1676037725
transform 1 0 39284 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_422
timestamp 1676037725
transform 1 0 39928 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_434
timestamp 1676037725
transform 1 0 41032 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_442
timestamp 1676037725
transform 1 0 41768 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1676037725
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_471
timestamp 1676037725
transform 1 0 44436 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_480
timestamp 1676037725
transform 1 0 45264 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_492
timestamp 1676037725
transform 1 0 46368 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1676037725
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_276
timestamp 1676037725
transform 1 0 26496 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_282
timestamp 1676037725
transform 1 0 27048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_292
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1676037725
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1676037725
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_324
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_336
timestamp 1676037725
transform 1 0 32016 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1676037725
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_376
timestamp 1676037725
transform 1 0 35696 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_383
timestamp 1676037725
transform 1 0 36340 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_390
timestamp 1676037725
transform 1 0 36984 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_402
timestamp 1676037725
transform 1 0 38088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_414
timestamp 1676037725
transform 1 0 39192 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_427
timestamp 1676037725
transform 1 0 40388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_437
timestamp 1676037725
transform 1 0 41308 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_461
timestamp 1676037725
transform 1 0 43516 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_473
timestamp 1676037725
transform 1 0 44620 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1676037725
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_237
timestamp 1676037725
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_253
timestamp 1676037725
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_265
timestamp 1676037725
transform 1 0 25484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1676037725
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_296
timestamp 1676037725
transform 1 0 28336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_300
timestamp 1676037725
transform 1 0 28704 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_310
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_344
timestamp 1676037725
transform 1 0 32752 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_374
timestamp 1676037725
transform 1 0 35512 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_386
timestamp 1676037725
transform 1 0 36616 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_409
timestamp 1676037725
transform 1 0 38732 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_413
timestamp 1676037725
transform 1 0 39100 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_425
timestamp 1676037725
transform 1 0 40204 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_437
timestamp 1676037725
transform 1 0 41308 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1676037725
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_460
timestamp 1676037725
transform 1 0 43424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_468
timestamp 1676037725
transform 1 0 44160 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_479
timestamp 1676037725
transform 1 0 45172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_491
timestamp 1676037725
transform 1 0 46276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1676037725
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1676037725
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_275
timestamp 1676037725
transform 1 0 26404 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_283
timestamp 1676037725
transform 1 0 27140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_341
timestamp 1676037725
transform 1 0 32476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_370
timestamp 1676037725
transform 1 0 35144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_382
timestamp 1676037725
transform 1 0 36248 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_387
timestamp 1676037725
transform 1 0 36708 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_399
timestamp 1676037725
transform 1 0 37812 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_405
timestamp 1676037725
transform 1 0 38364 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_415
timestamp 1676037725
transform 1 0 39284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_443
timestamp 1676037725
transform 1 0 41860 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_467
timestamp 1676037725
transform 1 0 44068 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_482
timestamp 1676037725
transform 1 0 45448 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_494
timestamp 1676037725
transform 1 0 46552 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_506
timestamp 1676037725
transform 1 0 47656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_245
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_266
timestamp 1676037725
transform 1 0 25576 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1676037725
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_303
timestamp 1676037725
transform 1 0 28980 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_311
timestamp 1676037725
transform 1 0 29716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_377
timestamp 1676037725
transform 1 0 35788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1676037725
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_425
timestamp 1676037725
transform 1 0 40204 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_437
timestamp 1676037725
transform 1 0 41308 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_445
timestamp 1676037725
transform 1 0 42044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_457
timestamp 1676037725
transform 1 0 43148 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_474
timestamp 1676037725
transform 1 0 44712 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_481
timestamp 1676037725
transform 1 0 45356 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_493
timestamp 1676037725
transform 1 0 46460 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_501
timestamp 1676037725
transform 1 0 47196 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1676037725
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1676037725
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_342
timestamp 1676037725
transform 1 0 32568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_355
timestamp 1676037725
transform 1 0 33764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1676037725
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_388
timestamp 1676037725
transform 1 0 36800 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_396
timestamp 1676037725
transform 1 0 37536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_402
timestamp 1676037725
transform 1 0 38088 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_411
timestamp 1676037725
transform 1 0 38916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_453
timestamp 1676037725
transform 1 0 42780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_463
timestamp 1676037725
transform 1 0 43700 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_470
timestamp 1676037725
transform 1 0 44344 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1676037725
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1676037725
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_249
timestamp 1676037725
transform 1 0 24012 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_260
timestamp 1676037725
transform 1 0 25024 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_264
timestamp 1676037725
transform 1 0 25392 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_274
timestamp 1676037725
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1676037725
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_296
timestamp 1676037725
transform 1 0 28336 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1676037725
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1676037725
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_351
timestamp 1676037725
transform 1 0 33396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_363
timestamp 1676037725
transform 1 0 34500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_386
timestamp 1676037725
transform 1 0 36616 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_404
timestamp 1676037725
transform 1 0 38272 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1676037725
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1676037725
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_462
timestamp 1676037725
transform 1 0 43608 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_486
timestamp 1676037725
transform 1 0 45816 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_498
timestamp 1676037725
transform 1 0 46920 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1676037725
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1676037725
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1676037725
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1676037725
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1676037725
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_392
timestamp 1676037725
transform 1 0 37168 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_399
timestamp 1676037725
transform 1 0 37812 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_407
timestamp 1676037725
transform 1 0 38548 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1676037725
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_468
timestamp 1676037725
transform 1 0 44160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_499
timestamp 1676037725
transform 1 0 47012 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_507
timestamp 1676037725
transform 1 0 47748 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1676037725
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1676037725
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1676037725
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1676037725
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1676037725
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_360
timestamp 1676037725
transform 1 0 34224 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_372
timestamp 1676037725
transform 1 0 35328 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_384
timestamp 1676037725
transform 1 0 36432 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_404
timestamp 1676037725
transform 1 0 38272 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_432
timestamp 1676037725
transform 1 0 40848 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_445
timestamp 1676037725
transform 1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_460
timestamp 1676037725
transform 1 0 43424 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_464
timestamp 1676037725
transform 1 0 43792 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_469
timestamp 1676037725
transform 1 0 44252 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_475
timestamp 1676037725
transform 1 0 44804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_496
timestamp 1676037725
transform 1 0 46736 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1676037725
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1676037725
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_275
timestamp 1676037725
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_287
timestamp 1676037725
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_299
timestamp 1676037725
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_320
timestamp 1676037725
transform 1 0 30544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_333
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_341
timestamp 1676037725
transform 1 0 32476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_354
timestamp 1676037725
transform 1 0 33672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_411
timestamp 1676037725
transform 1 0 38916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1676037725
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_427
timestamp 1676037725
transform 1 0 40388 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_448
timestamp 1676037725
transform 1 0 42320 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_455
timestamp 1676037725
transform 1 0 42964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_459
timestamp 1676037725
transform 1 0 43332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1676037725
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_483
timestamp 1676037725
transform 1 0 45540 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_490
timestamp 1676037725
transform 1 0 46184 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_502
timestamp 1676037725
transform 1 0 47288 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_508
timestamp 1676037725
transform 1 0 47840 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_261
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_265
timestamp 1676037725
transform 1 0 25484 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1676037725
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_304
timestamp 1676037725
transform 1 0 29072 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_328
timestamp 1676037725
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_359
timestamp 1676037725
transform 1 0 34132 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_367
timestamp 1676037725
transform 1 0 34868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_377
timestamp 1676037725
transform 1 0 35788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1676037725
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_400
timestamp 1676037725
transform 1 0 37904 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_413
timestamp 1676037725
transform 1 0 39100 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_421
timestamp 1676037725
transform 1 0 39836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_431
timestamp 1676037725
transform 1 0 40756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1676037725
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_457
timestamp 1676037725
transform 1 0 43148 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_469
timestamp 1676037725
transform 1 0 44252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_493
timestamp 1676037725
transform 1 0 46460 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_501
timestamp 1676037725
transform 1 0 47196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1676037725
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_269
timestamp 1676037725
transform 1 0 25852 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_279
timestamp 1676037725
transform 1 0 26772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_291
timestamp 1676037725
transform 1 0 27876 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1676037725
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_331
timestamp 1676037725
transform 1 0 31556 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_355
timestamp 1676037725
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1676037725
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_376
timestamp 1676037725
transform 1 0 35696 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_383
timestamp 1676037725
transform 1 0 36340 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_395
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_407
timestamp 1676037725
transform 1 0 38548 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_412
timestamp 1676037725
transform 1 0 39008 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_442
timestamp 1676037725
transform 1 0 41768 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_454
timestamp 1676037725
transform 1 0 42872 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_460
timestamp 1676037725
transform 1 0 43424 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_470
timestamp 1676037725
transform 1 0 44344 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_488
timestamp 1676037725
transform 1 0 46000 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_495
timestamp 1676037725
transform 1 0 46644 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_507
timestamp 1676037725
transform 1 0 47748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_519
timestamp 1676037725
transform 1 0 48852 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_317
timestamp 1676037725
transform 1 0 30268 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1676037725
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_348
timestamp 1676037725
transform 1 0 33120 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_352
timestamp 1676037725
transform 1 0 33488 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_373
timestamp 1676037725
transform 1 0 35420 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1676037725
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_401
timestamp 1676037725
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_408
timestamp 1676037725
transform 1 0 38640 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_420
timestamp 1676037725
transform 1 0 39744 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_432
timestamp 1676037725
transform 1 0 40848 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1676037725
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_460
timestamp 1676037725
transform 1 0 43424 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_488
timestamp 1676037725
transform 1 0 46000 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1676037725
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_525
timestamp 1676037725
transform 1 0 49404 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1676037725
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1676037725
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_315
timestamp 1676037725
transform 1 0 30084 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1676037725
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_349
timestamp 1676037725
transform 1 0 33212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1676037725
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_376
timestamp 1676037725
transform 1 0 35696 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_384
timestamp 1676037725
transform 1 0 36432 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_390
timestamp 1676037725
transform 1 0 36984 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_403
timestamp 1676037725
transform 1 0 38180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_415
timestamp 1676037725
transform 1 0 39284 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1676037725
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_443
timestamp 1676037725
transform 1 0 41860 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_467
timestamp 1676037725
transform 1 0 44068 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1676037725
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_488
timestamp 1676037725
transform 1 0 46000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_500
timestamp 1676037725
transform 1 0 47104 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_508
timestamp 1676037725
transform 1 0 47840 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_525
timestamp 1676037725
transform 1 0 49404 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_303
timestamp 1676037725
transform 1 0 28980 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_315
timestamp 1676037725
transform 1 0 30084 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_320
timestamp 1676037725
transform 1 0 30544 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1676037725
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_342
timestamp 1676037725
transform 1 0 32568 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_368
timestamp 1676037725
transform 1 0 34960 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_381
timestamp 1676037725
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 1676037725
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_397
timestamp 1676037725
transform 1 0 37628 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_401
timestamp 1676037725
transform 1 0 37996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_426
timestamp 1676037725
transform 1 0 40296 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_434
timestamp 1676037725
transform 1 0 41032 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_446
timestamp 1676037725
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_471
timestamp 1676037725
transform 1 0 44436 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_495
timestamp 1676037725
transform 1 0 46644 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1676037725
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_525
timestamp 1676037725
transform 1 0 49404 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1676037725
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1676037725
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_277
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_285
timestamp 1676037725
transform 1 0 27324 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1676037725
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_317
timestamp 1676037725
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_340
timestamp 1676037725
transform 1 0 32384 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_352
timestamp 1676037725
transform 1 0 33488 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_376
timestamp 1676037725
transform 1 0 35696 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_388
timestamp 1676037725
transform 1 0 36800 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_399
timestamp 1676037725
transform 1 0 37812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_412
timestamp 1676037725
transform 1 0 39008 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_444
timestamp 1676037725
transform 1 0 41952 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_451
timestamp 1676037725
transform 1 0 42596 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_459
timestamp 1676037725
transform 1 0 43332 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_464
timestamp 1676037725
transform 1 0 43792 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_501
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_511
timestamp 1676037725
transform 1 0 48116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1676037725
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1676037725
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1676037725
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_317
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1676037725
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_343
timestamp 1676037725
transform 1 0 32660 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_353
timestamp 1676037725
transform 1 0 33580 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_365
timestamp 1676037725
transform 1 0 34684 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_376
timestamp 1676037725
transform 1 0 35696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1676037725
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_397
timestamp 1676037725
transform 1 0 37628 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_418
timestamp 1676037725
transform 1 0 39560 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_430
timestamp 1676037725
transform 1 0 40664 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_436
timestamp 1676037725
transform 1 0 41216 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_446
timestamp 1676037725
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_478
timestamp 1676037725
transform 1 0 45080 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_490
timestamp 1676037725
transform 1 0 46184 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_502
timestamp 1676037725
transform 1 0 47288 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_517
timestamp 1676037725
transform 1 0 48668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_521
timestamp 1676037725
transform 1 0 49036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_525
timestamp 1676037725
transform 1 0 49404 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_275
timestamp 1676037725
transform 1 0 26404 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_287
timestamp 1676037725
transform 1 0 27508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1676037725
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_321
timestamp 1676037725
transform 1 0 30636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_342
timestamp 1676037725
transform 1 0 32568 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1676037725
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_373
timestamp 1676037725
transform 1 0 35420 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_383
timestamp 1676037725
transform 1 0 36340 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_391
timestamp 1676037725
transform 1 0 37076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_402
timestamp 1676037725
transform 1 0 38088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_409
timestamp 1676037725
transform 1 0 38732 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 1676037725
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_428
timestamp 1676037725
transform 1 0 40480 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_436
timestamp 1676037725
transform 1 0 41216 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_440
timestamp 1676037725
transform 1 0 41584 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_455
timestamp 1676037725
transform 1 0 42964 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_468
timestamp 1676037725
transform 1 0 44160 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1676037725
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1676037725
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_237
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_254
timestamp 1676037725
transform 1 0 24472 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_266
timestamp 1676037725
transform 1 0 25576 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1676037725
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_297
timestamp 1676037725
transform 1 0 28428 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_318
timestamp 1676037725
transform 1 0 30360 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_324
timestamp 1676037725
transform 1 0 30912 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1676037725
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_369
timestamp 1676037725
transform 1 0 35052 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1676037725
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_410
timestamp 1676037725
transform 1 0 38824 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_418
timestamp 1676037725
transform 1 0 39560 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_446
timestamp 1676037725
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_470
timestamp 1676037725
transform 1 0 44344 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_482
timestamp 1676037725
transform 1 0 45448 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_494
timestamp 1676037725
transform 1 0 46552 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_502
timestamp 1676037725
transform 1 0 47288 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_517
timestamp 1676037725
transform 1 0 48668 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_521
timestamp 1676037725
transform 1 0 49036 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_525
timestamp 1676037725
transform 1 0 49404 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1676037725
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1676037725
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_337
timestamp 1676037725
transform 1 0 32108 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_352
timestamp 1676037725
transform 1 0 33488 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_376
timestamp 1676037725
transform 1 0 35696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_382
timestamp 1676037725
transform 1 0 36248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_410
timestamp 1676037725
transform 1 0 38824 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_417
timestamp 1676037725
transform 1 0 39468 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_443
timestamp 1676037725
transform 1 0 41860 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_467
timestamp 1676037725
transform 1 0 44068 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1676037725
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_521
timestamp 1676037725
transform 1 0 49036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1676037725
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1676037725
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1676037725
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1676037725
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1676037725
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1676037725
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_350
timestamp 1676037725
transform 1 0 33304 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_356
timestamp 1676037725
transform 1 0 33856 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_369
timestamp 1676037725
transform 1 0 35052 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1676037725
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_415
timestamp 1676037725
transform 1 0 39284 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_439
timestamp 1676037725
transform 1 0 41492 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_471
timestamp 1676037725
transform 1 0 44436 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_483
timestamp 1676037725
transform 1 0 45540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_495
timestamp 1676037725
transform 1 0 46644 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_525
timestamp 1676037725
transform 1 0 49404 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1676037725
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1676037725
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1676037725
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1676037725
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_321
timestamp 1676037725
transform 1 0 30636 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_327
timestamp 1676037725
transform 1 0 31188 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_349
timestamp 1676037725
transform 1 0 33212 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_357
timestamp 1676037725
transform 1 0 33948 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1676037725
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_376
timestamp 1676037725
transform 1 0 35696 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_382
timestamp 1676037725
transform 1 0 36248 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_394
timestamp 1676037725
transform 1 0 37352 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_406
timestamp 1676037725
transform 1 0 38456 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_418
timestamp 1676037725
transform 1 0 39560 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_464
timestamp 1676037725
transform 1 0 43792 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_521
timestamp 1676037725
transform 1 0 49036 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1676037725
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1676037725
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1676037725
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1676037725
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1676037725
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1676037725
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1676037725
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_365
timestamp 1676037725
transform 1 0 34684 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_378
timestamp 1676037725
transform 1 0 35880 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 1676037725
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_401
timestamp 1676037725
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_422
timestamp 1676037725
transform 1 0 39928 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_430
timestamp 1676037725
transform 1 0 40664 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_440
timestamp 1676037725
transform 1 0 41584 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_471
timestamp 1676037725
transform 1 0 44436 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_483
timestamp 1676037725
transform 1 0 45540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_495
timestamp 1676037725
transform 1 0 46644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_521
timestamp 1676037725
transform 1 0 49036 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_525
timestamp 1676037725
transform 1 0 49404 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_221
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_229
timestamp 1676037725
transform 1 0 22172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_240
timestamp 1676037725
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1676037725
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1676037725
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_333
timestamp 1676037725
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_341
timestamp 1676037725
transform 1 0 32476 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_355
timestamp 1676037725
transform 1 0 33764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_384
timestamp 1676037725
transform 1 0 36432 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_396
timestamp 1676037725
transform 1 0 37536 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_408
timestamp 1676037725
transform 1 0 38640 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_434
timestamp 1676037725
transform 1 0 41032 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_458
timestamp 1676037725
transform 1 0 43240 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_470
timestamp 1676037725
transform 1 0 44344 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1676037725
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_525
timestamp 1676037725
transform 1 0 49404 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1676037725
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1676037725
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_349
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_355
timestamp 1676037725
transform 1 0 33764 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_358
timestamp 1676037725
transform 1 0 34040 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_371
timestamp 1676037725
transform 1 0 35236 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_383
timestamp 1676037725
transform 1 0 36340 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1676037725
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_399
timestamp 1676037725
transform 1 0 37812 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_420
timestamp 1676037725
transform 1 0 39744 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_446
timestamp 1676037725
transform 1 0 42136 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_457
timestamp 1676037725
transform 1 0 43148 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_468
timestamp 1676037725
transform 1 0 44160 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_480
timestamp 1676037725
transform 1 0 45264 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_492
timestamp 1676037725
transform 1 0 46368 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_517
timestamp 1676037725
transform 1 0 48668 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_521
timestamp 1676037725
transform 1 0 49036 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_525
timestamp 1676037725
transform 1 0 49404 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1676037725
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1676037725
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1676037725
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1676037725
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1676037725
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1676037725
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1676037725
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1676037725
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1676037725
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_443
timestamp 1676037725
transform 1 0 41860 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_451
timestamp 1676037725
transform 1 0 42596 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_454
timestamp 1676037725
transform 1 0 42872 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_467
timestamp 1676037725
transform 1 0 44068 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1676037725
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_513
timestamp 1676037725
transform 1 0 48300 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_521
timestamp 1676037725
transform 1 0 49036 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1676037725
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1676037725
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1676037725
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1676037725
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1676037725
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1676037725
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1676037725
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1676037725
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_426
timestamp 1676037725
transform 1 0 40296 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_438
timestamp 1676037725
transform 1 0 41400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_446
timestamp 1676037725
transform 1 0 42136 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1676037725
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1676037725
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1676037725
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1676037725
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_517
timestamp 1676037725
transform 1 0 48668 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_525
timestamp 1676037725
transform 1 0 49404 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1676037725
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1676037725
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1676037725
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1676037725
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1676037725
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1676037725
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1676037725
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1676037725
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1676037725
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1676037725
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1676037725
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1676037725
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1676037725
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_521
timestamp 1676037725
transform 1 0 49036 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1676037725
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1676037725
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1676037725
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1676037725
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1676037725
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1676037725
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1676037725
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1676037725
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1676037725
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1676037725
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1676037725
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1676037725
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1676037725
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1676037725
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1676037725
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_460
timestamp 1676037725
transform 1 0 43424 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_466
timestamp 1676037725
transform 1 0 43976 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_478
timestamp 1676037725
transform 1 0 45080 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_490
timestamp 1676037725
transform 1 0 46184 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_502
timestamp 1676037725
transform 1 0 47288 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_521
timestamp 1676037725
transform 1 0 49036 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_525
timestamp 1676037725
transform 1 0 49404 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1676037725
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_233
timestamp 1676037725
transform 1 0 22540 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_239
timestamp 1676037725
transform 1 0 23092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1676037725
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1676037725
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1676037725
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1676037725
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1676037725
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1676037725
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1676037725
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1676037725
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1676037725
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1676037725
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1676037725
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1676037725
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_429
timestamp 1676037725
transform 1 0 40572 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_442
timestamp 1676037725
transform 1 0 41768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_455
timestamp 1676037725
transform 1 0 42964 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_461
timestamp 1676037725
transform 1 0 43516 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_473
timestamp 1676037725
transform 1 0 44620 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_257
timestamp 1676037725
transform 1 0 24748 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_269
timestamp 1676037725
transform 1 0 25852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1676037725
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1676037725
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1676037725
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1676037725
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1676037725
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1676037725
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1676037725
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1676037725
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1676037725
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1676037725
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1676037725
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1676037725
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1676037725
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1676037725
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1676037725
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1676037725
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1676037725
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_521
timestamp 1676037725
transform 1 0 49036 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_525
timestamp 1676037725
transform 1 0 49404 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1676037725
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1676037725
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1676037725
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1676037725
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1676037725
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1676037725
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1676037725
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1676037725
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1676037725
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1676037725
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1676037725
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1676037725
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1676037725
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1676037725
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1676037725
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1676037725
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1676037725
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_521
timestamp 1676037725
transform 1 0 49036 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1676037725
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1676037725
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1676037725
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1676037725
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1676037725
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1676037725
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1676037725
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1676037725
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1676037725
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1676037725
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1676037725
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1676037725
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1676037725
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1676037725
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1676037725
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1676037725
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1676037725
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1676037725
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1676037725
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1676037725
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1676037725
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1676037725
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1676037725
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1676037725
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1676037725
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1676037725
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1676037725
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_525
timestamp 1676037725
transform 1 0 49404 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1676037725
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1676037725
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1676037725
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1676037725
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1676037725
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1676037725
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1676037725
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1676037725
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1676037725
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1676037725
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1676037725
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1676037725
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1676037725
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1676037725
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1676037725
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1676037725
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1676037725
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_521
timestamp 1676037725
transform 1 0 49036 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1676037725
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1676037725
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1676037725
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1676037725
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1676037725
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1676037725
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1676037725
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1676037725
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1676037725
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1676037725
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1676037725
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1676037725
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1676037725
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1676037725
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1676037725
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1676037725
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1676037725
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1676037725
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1676037725
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1676037725
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_525
timestamp 1676037725
transform 1 0 49404 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_205
timestamp 1676037725
transform 1 0 19964 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_211
timestamp 1676037725
transform 1 0 20516 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_223
timestamp 1676037725
transform 1 0 21620 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_235
timestamp 1676037725
transform 1 0 22724 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1676037725
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1676037725
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1676037725
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1676037725
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1676037725
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1676037725
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1676037725
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1676037725
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1676037725
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1676037725
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1676037725
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1676037725
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1676037725
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1676037725
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1676037725
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1676037725
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1676037725
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1676037725
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1676037725
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1676037725
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1676037725
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1676037725
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1676037725
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1676037725
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1676037725
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1676037725
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1676037725
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1676037725
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1676037725
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1676037725
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1676037725
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1676037725
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1676037725
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1676037725
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1676037725
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_525
timestamp 1676037725
transform 1 0 49404 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1676037725
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1676037725
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1676037725
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1676037725
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1676037725
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1676037725
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1676037725
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1676037725
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1676037725
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1676037725
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1676037725
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1676037725
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1676037725
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1676037725
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1676037725
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1676037725
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1676037725
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1676037725
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_521
timestamp 1676037725
transform 1 0 49036 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1676037725
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1676037725
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1676037725
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1676037725
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1676037725
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1676037725
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1676037725
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1676037725
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1676037725
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1676037725
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1676037725
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1676037725
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1676037725
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_525
timestamp 1676037725
transform 1 0 49404 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1676037725
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1676037725
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1676037725
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1676037725
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1676037725
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1676037725
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1676037725
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1676037725
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1676037725
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1676037725
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1676037725
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1676037725
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1676037725
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1676037725
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1676037725
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1676037725
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1676037725
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_521
timestamp 1676037725
transform 1 0 49036 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1676037725
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1676037725
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1676037725
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1676037725
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1676037725
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1676037725
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1676037725
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1676037725
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1676037725
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1676037725
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1676037725
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1676037725
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1676037725
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1676037725
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_517
timestamp 1676037725
transform 1 0 48668 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_521
timestamp 1676037725
transform 1 0 49036 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_525
timestamp 1676037725
transform 1 0 49404 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1676037725
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1676037725
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1676037725
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1676037725
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1676037725
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1676037725
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1676037725
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1676037725
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1676037725
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1676037725
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1676037725
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1676037725
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1676037725
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1676037725
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1676037725
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1676037725
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1676037725
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1676037725
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1676037725
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1676037725
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1676037725
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1676037725
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1676037725
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1676037725
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1676037725
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1676037725
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1676037725
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1676037725
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1676037725
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1676037725
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1676037725
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1676037725
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1676037725
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1676037725
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_517
timestamp 1676037725
transform 1 0 48668 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_521
timestamp 1676037725
transform 1 0 49036 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_525
timestamp 1676037725
transform 1 0 49404 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_242
timestamp 1676037725
transform 1 0 23368 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1676037725
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1676037725
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1676037725
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1676037725
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1676037725
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1676037725
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1676037725
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1676037725
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1676037725
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1676037725
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1676037725
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1676037725
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1676037725
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1676037725
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1676037725
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_525
timestamp 1676037725
transform 1 0 49404 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1676037725
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1676037725
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_213
timestamp 1676037725
transform 1 0 20700 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1676037725
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_239
timestamp 1676037725
transform 1 0 23092 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_251
timestamp 1676037725
transform 1 0 24196 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_263
timestamp 1676037725
transform 1 0 25300 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_275
timestamp 1676037725
transform 1 0 26404 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1676037725
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1676037725
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1676037725
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1676037725
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1676037725
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1676037725
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1676037725
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1676037725
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1676037725
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1676037725
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1676037725
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1676037725
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1676037725
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1676037725
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1676037725
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_517
timestamp 1676037725
transform 1 0 48668 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_525
timestamp 1676037725
transform 1 0 49404 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1676037725
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1676037725
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1676037725
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1676037725
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1676037725
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1676037725
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1676037725
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1676037725
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1676037725
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1676037725
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1676037725
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1676037725
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1676037725
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1676037725
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1676037725
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1676037725
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1676037725
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1676037725
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1676037725
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1676037725
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1676037725
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1676037725
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1676037725
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1676037725
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1676037725
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1676037725
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1676037725
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1676037725
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1676037725
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1676037725
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1676037725
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1676037725
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1676037725
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1676037725
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1676037725
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1676037725
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1676037725
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1676037725
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1676037725
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1676037725
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1676037725
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_517
timestamp 1676037725
transform 1 0 48668 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_525
timestamp 1676037725
transform 1 0 49404 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1676037725
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1676037725
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1676037725
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1676037725
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1676037725
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1676037725
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1676037725
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1676037725
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1676037725
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1676037725
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1676037725
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1676037725
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1676037725
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1676037725
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1676037725
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_460
timestamp 1676037725
transform 1 0 43424 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_472
timestamp 1676037725
transform 1 0 44528 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1676037725
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1676037725
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1676037725
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_213
timestamp 1676037725
transform 1 0 20700 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_221
timestamp 1676037725
transform 1 0 21436 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_231
timestamp 1676037725
transform 1 0 22356 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_238
timestamp 1676037725
transform 1 0 23000 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_250
timestamp 1676037725
transform 1 0 24104 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_262
timestamp 1676037725
transform 1 0 25208 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_274
timestamp 1676037725
transform 1 0 26312 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1676037725
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1676037725
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1676037725
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1676037725
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1676037725
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1676037725
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1676037725
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1676037725
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1676037725
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1676037725
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1676037725
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1676037725
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1676037725
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1676037725
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_525
timestamp 1676037725
transform 1 0 49404 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_219
timestamp 1676037725
transform 1 0 21252 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_231
timestamp 1676037725
transform 1 0 22356 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_243
timestamp 1676037725
transform 1 0 23460 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1676037725
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1676037725
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1676037725
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1676037725
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1676037725
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1676037725
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1676037725
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1676037725
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1676037725
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1676037725
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1676037725
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1676037725
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1676037725
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1676037725
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_521
timestamp 1676037725
transform 1 0 49036 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_525
timestamp 1676037725
transform 1 0 49404 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1676037725
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1676037725
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_272
timestamp 1676037725
transform 1 0 26128 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1676037725
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_330
timestamp 1676037725
transform 1 0 31464 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1676037725
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1676037725
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1676037725
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1676037725
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1676037725
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1676037725
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1676037725
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1676037725
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1676037725
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1676037725
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_517
timestamp 1676037725
transform 1 0 48668 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_525
timestamp 1676037725
transform 1 0 49404 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_173
timestamp 1676037725
transform 1 0 17020 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_182
timestamp 1676037725
transform 1 0 17848 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1676037725
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_217
timestamp 1676037725
transform 1 0 21068 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_224
timestamp 1676037725
transform 1 0 21712 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_236
timestamp 1676037725
transform 1 0 22816 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1676037725
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_258
timestamp 1676037725
transform 1 0 24840 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_270
timestamp 1676037725
transform 1 0 25944 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_282
timestamp 1676037725
transform 1 0 27048 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1676037725
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1676037725
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1676037725
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1676037725
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1676037725
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1676037725
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1676037725
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1676037725
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1676037725
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1676037725
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_513
timestamp 1676037725
transform 1 0 48300 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_521
timestamp 1676037725
transform 1 0 49036 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1676037725
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1676037725
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1676037725
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1676037725
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1676037725
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1676037725
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1676037725
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1676037725
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1676037725
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1676037725
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1676037725
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1676037725
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1676037725
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1676037725
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_521
timestamp 1676037725
transform 1 0 49036 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_525
timestamp 1676037725
transform 1 0 49404 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1676037725
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_229
timestamp 1676037725
transform 1 0 22172 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_288
timestamp 1676037725
transform 1 0 27600 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1676037725
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1676037725
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1676037725
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1676037725
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1676037725
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1676037725
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1676037725
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_525
timestamp 1676037725
transform 1 0 49404 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_197
timestamp 1676037725
transform 1 0 19228 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_204
timestamp 1676037725
transform 1 0 19872 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_211
timestamp 1676037725
transform 1 0 20516 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1676037725
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1676037725
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1676037725
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1676037725
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1676037725
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1676037725
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1676037725
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1676037725
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1676037725
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1676037725
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1676037725
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1676037725
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1676037725
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1676037725
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1676037725
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1676037725
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_521
timestamp 1676037725
transform 1 0 49036 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_525
timestamp 1676037725
transform 1 0 49404 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1676037725
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1676037725
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1676037725
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1676037725
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1676037725
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1676037725
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1676037725
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1676037725
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1676037725
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1676037725
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1676037725
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1676037725
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1676037725
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1676037725
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_513
timestamp 1676037725
transform 1 0 48300 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_525
timestamp 1676037725
transform 1 0 49404 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1676037725
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1676037725
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1676037725
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1676037725
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1676037725
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1676037725
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1676037725
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1676037725
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_525
timestamp 1676037725
transform 1 0 49404 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1676037725
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_213
timestamp 1676037725
transform 1 0 20700 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_218
timestamp 1676037725
transform 1 0 21160 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_230
timestamp 1676037725
transform 1 0 22264 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_240
timestamp 1676037725
transform 1 0 23184 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1676037725
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1676037725
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1676037725
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1676037725
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1676037725
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1676037725
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1676037725
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1676037725
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1676037725
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1676037725
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1676037725
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1676037725
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1676037725
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1676037725
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1676037725
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1676037725
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1676037725
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1676037725
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1676037725
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1676037725
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1676037725
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1676037725
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1676037725
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1676037725
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1676037725
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1676037725
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1676037725
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1676037725
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1676037725
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1676037725
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1676037725
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1676037725
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1676037725
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1676037725
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_525
timestamp 1676037725
transform 1 0 49404 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1676037725
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1676037725
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_159
timestamp 1676037725
transform 1 0 15732 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_171
timestamp 1676037725
transform 1 0 16836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_183
timestamp 1676037725
transform 1 0 17940 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_203
timestamp 1676037725
transform 1 0 19780 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_215
timestamp 1676037725
transform 1 0 20884 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_227
timestamp 1676037725
transform 1 0 21988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_239
timestamp 1676037725
transform 1 0 23092 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1676037725
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1676037725
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1676037725
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1676037725
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1676037725
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_525
timestamp 1676037725
transform 1 0 49404 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1676037725
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1676037725
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1676037725
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1676037725
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1676037725
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1676037725
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1676037725
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1676037725
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1676037725
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1676037725
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1676037725
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1676037725
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1676037725
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1676037725
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1676037725
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_517
timestamp 1676037725
transform 1 0 48668 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_525
timestamp 1676037725
transform 1 0 49404 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1676037725
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1676037725
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1676037725
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_168
timestamp 1676037725
transform 1 0 16560 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_172
timestamp 1676037725
transform 1 0 16928 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1676037725
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1676037725
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1676037725
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1676037725
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1676037725
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1676037725
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1676037725
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1676037725
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1676037725
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1676037725
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1676037725
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1676037725
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_513
timestamp 1676037725
transform 1 0 48300 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_90_525
timestamp 1676037725
transform 1 0 49404 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1676037725
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1676037725
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1676037725
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1676037725
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1676037725
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1676037725
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_129
timestamp 1676037725
transform 1 0 12972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_141
timestamp 1676037725
transform 1 0 14076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_153
timestamp 1676037725
transform 1 0 15180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_165
timestamp 1676037725
transform 1 0 16284 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1676037725
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_517
timestamp 1676037725
transform 1 0 48668 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_525
timestamp 1676037725
transform 1 0 49404 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1676037725
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1676037725
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1676037725
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1676037725
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1676037725
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1676037725
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1676037725
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1676037725
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1676037725
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1676037725
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1676037725
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1676037725
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1676037725
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_513
timestamp 1676037725
transform 1 0 48300 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_92_525
timestamp 1676037725
transform 1 0 49404 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1676037725
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1676037725
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1676037725
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1676037725
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1676037725
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_97
timestamp 1676037725
transform 1 0 10028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_109
timestamp 1676037725
transform 1 0 11132 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1676037725
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1676037725
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1676037725
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1676037725
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1676037725
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1676037725
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_517
timestamp 1676037725
transform 1 0 48668 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_525
timestamp 1676037725
transform 1 0 49404 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1676037725
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1676037725
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1676037725
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1676037725
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1676037725
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1676037725
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1676037725
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1676037725
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1676037725
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1676037725
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1676037725
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1676037725
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1676037725
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1676037725
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1676037725
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1676037725
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1676037725
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1676037725
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1676037725
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1676037725
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1676037725
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1676037725
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1676037725
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1676037725
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1676037725
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1676037725
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1676037725
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1676037725
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1676037725
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_501
timestamp 1676037725
transform 1 0 47196 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_505
timestamp 1676037725
transform 1 0 47564 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_509
timestamp 1676037725
transform 1 0 47932 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_517
timestamp 1676037725
transform 1 0 48668 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_525
timestamp 1676037725
transform 1 0 49404 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_21
timestamp 1676037725
transform 1 0 3036 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_27
timestamp 1676037725
transform 1 0 3588 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_49
timestamp 1676037725
transform 1 0 5612 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1676037725
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_61
timestamp 1676037725
transform 1 0 6716 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_78
timestamp 1676037725
transform 1 0 8280 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_107
timestamp 1676037725
transform 1 0 10948 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1676037725
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_119
timestamp 1676037725
transform 1 0 12052 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_136
timestamp 1676037725
transform 1 0 13616 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_165
timestamp 1676037725
transform 1 0 16284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_177
timestamp 1676037725
transform 1 0 17388 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_194
timestamp 1676037725
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_222
timestamp 1676037725
transform 1 0 21528 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_233
timestamp 1676037725
transform 1 0 22540 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_268
timestamp 1676037725
transform 1 0 25760 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_293
timestamp 1676037725
transform 1 0 28060 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_297
timestamp 1676037725
transform 1 0 28428 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_305
timestamp 1676037725
transform 1 0 29164 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_309
timestamp 1676037725
transform 1 0 29532 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_321
timestamp 1676037725
transform 1 0 30636 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_326
timestamp 1676037725
transform 1 0 31096 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_334
timestamp 1676037725
transform 1 0 31832 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_349
timestamp 1676037725
transform 1 0 33212 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_355
timestamp 1676037725
transform 1 0 33764 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_363
timestamp 1676037725
transform 1 0 34500 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_365
timestamp 1676037725
transform 1 0 34684 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_377
timestamp 1676037725
transform 1 0 35788 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1676037725
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1676037725
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_405
timestamp 1676037725
transform 1 0 38364 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_409
timestamp 1676037725
transform 1 0 38732 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_414
timestamp 1676037725
transform 1 0 39192 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_421
timestamp 1676037725
transform 1 0 39836 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_433
timestamp 1676037725
transform 1 0 40940 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_443
timestamp 1676037725
transform 1 0 41860 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1676037725
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_461
timestamp 1676037725
transform 1 0 43516 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_467
timestamp 1676037725
transform 1 0 44068 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_472
timestamp 1676037725
transform 1 0 44528 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_477
timestamp 1676037725
transform 1 0 44988 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_489
timestamp 1676037725
transform 1 0 46092 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_495
timestamp 1676037725
transform 1 0 46644 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_502
timestamp 1676037725
transform 1 0 47288 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_517
timestamp 1676037725
transform 1 0 48668 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_525
timestamp 1676037725
transform 1 0 49404 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 47656 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 48484 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 49128 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 49128 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 49128 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 49036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 49036 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 49128 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 49128 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 49128 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 49128 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 49036 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 49128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 49036 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 49036 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 49036 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 49128 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 49128 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 49128 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 49128 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1676037725
transform 1 0 49036 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 49036 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1676037725
transform 1 0 49036 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 49128 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 49128 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 49128 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 49128 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 49128 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 49128 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 49128 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 49128 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1676037725
transform 1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1676037725
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1676037725
transform 1 0 19228 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 19964 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 21160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 22172 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 23184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1676037725
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 6716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1676037725
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 25484 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 28152 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 30820 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 33488 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 36156 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input68
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 48852 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1676037725
transform 1 0 48852 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1676037725
transform 1 0 48852 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 49036 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 49036 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 49036 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform 1 0 48300 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 38824 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 41492 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 44160 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1676037725
transform 1 0 46736 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 1564 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 47932 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 47932 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 47932 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 47932 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 47932 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 47932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 47932 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 47932 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 47932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 47932 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 47932 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 47932 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 34132 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 33948 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 34868 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 36708 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 39284 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 39100 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 40020 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 41860 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 42596 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 44436 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 45172 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 44252 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 47748 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 25208 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 27324 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 29716 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 31556 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 4140 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 6808 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 9476 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 12144 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 17480 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 20056 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 22632 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 49864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 49864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 49864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 49864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 49864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 49864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 49864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 49864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 49864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 49864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 49864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 49864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 49864 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 49864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 49864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 49864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 49864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 49864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 49864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 49864 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 49864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 49864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 49864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 49864 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 49864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 49864 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 49864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 49864 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 49864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 49864 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 49864 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 49864 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 49864 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 49864 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 49864 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 49864 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 49864 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 49864 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 49864 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 49864 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 49864 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 49864 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 49864 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 49864 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 49864 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 49864 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 49864 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 49864 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 49864 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 49864 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 49864 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 49864 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 49864 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 49864 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 49864 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35420 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 41676 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 42596 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 42228 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40204 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 39008 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40480 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 42320 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 43976 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 45172 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 44896 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 44160 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 44804 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 42596 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 42228 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38456 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37720 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 36984 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 39652 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 42228 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 42596 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 42596 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 41400 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40296 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38456 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37904 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38088 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40112 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 43976 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 41492 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 31280 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 27140 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28520 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28428 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 27416 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30268 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30728 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 30544 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33120 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33580 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 31924 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29440 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23736 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28428 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29900 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30728 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29992 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27692 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25300 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 26036 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27600 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32844 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33488 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32568 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33948 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34776 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34960 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32568 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31924 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29716 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31924 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33120 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34040 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35328 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 36248 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 36432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35604 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 39652 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38732 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 39008 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 39192 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 38916 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38456 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37720 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 36432 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33120 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 41216 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1__198
timestamp 1676037725
transform 1 0 37812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38456 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36248 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 42780 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 41860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 43424 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 41860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39284 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 37628 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38088 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38732 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36248 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 43516 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 41860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40020 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 45172 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0__199
timestamp 1676037725
transform 1 0 45080 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 43884 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40388 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 45172 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0__200
timestamp 1676037725
transform 1 0 44068 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 42872 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 44252 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0__201
timestamp 1676037725
transform 1 0 42688 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 43332 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0__202
timestamp 1676037725
transform 1 0 41492 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39928 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 41308 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 38732 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38272 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 35328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40756 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 37720 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37352 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 34132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40204 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 37536 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38180 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 34316 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 43332 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 42320 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 41308 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40020 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 43240 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 41308 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 41308 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 40204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39744 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 42136 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 39192 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37996 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36064 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 38456 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37260 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32384 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 42688 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 42228 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34408 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35052 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 31004 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 20332 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 28428 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36064 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32476 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 34224 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 31004 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30176 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 34868 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32936 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 28612 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38364 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 35604 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35512 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35328 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_6.mux_l2_in_1__192
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27876 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33396 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39284 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 34868 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 31004 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_8.mux_l2_in_1__193
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25024 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37536 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32752 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 22356 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20976 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28796 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36432 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 26404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27324 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32568 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28152 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32936 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30452 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_18.mux_l2_in_0__169
timestamp 1676037725
transform 1 0 33488 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33028 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39192 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28152 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 31556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32752 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37628 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23460 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 28612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28428 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24656 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30912 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 32108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37628 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 36340 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35144 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41032 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34960 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_28.mux_l1_in_1__175
timestamp 1676037725
transform 1 0 30452 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 30084 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40296 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 36156 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_30.mux_l1_in_1__176
timestamp 1676037725
transform 1 0 31556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36156 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41032 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 36156 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_32.mux_l1_in_1__177
timestamp 1676037725
transform 1 0 32292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 31096 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35052 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_34.mux_l1_in_1__178
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26036 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 31924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28244 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 32752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32016 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 35052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32752 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 37444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41216 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37812 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 42596 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 36340 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 33488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 33120 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37812 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 36248 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35052 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37996 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 42228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 38640 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 34592 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 34868 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38732 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 42596 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_50.mux_l2_in_0__187
timestamp 1676037725
transform 1 0 41308 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40112 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 35604 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_52.mux_l2_in_0__188
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39928 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 43056 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34592 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_54.mux_l2_in_0__189
timestamp 1676037725
transform 1 0 38272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38640 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_56.mux_l2_in_0__190
timestamp 1676037725
transform 1 0 37536 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38272 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_58.mux_l1_in_1__191
timestamp 1676037725
transform 1 0 23092 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22724 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38548 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 29440 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 34592 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 39744 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 44896 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 49422 56200 49478 57000 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 50200 688 51000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1398 56200 1454 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 50200 25984 51000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 50200 34144 51000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 50200 34960 51000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 50200 35776 51000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 50200 36592 51000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 50200 37408 51000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 50200 38224 51000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 50200 39040 51000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 50200 39856 51000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 50200 40672 51000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 50200 41488 51000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 50200 26800 51000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 50200 42304 51000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 50200 43120 51000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 50200 43936 51000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 50200 44752 51000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 50200 45568 51000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 50200 46384 51000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 50200 47200 51000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 50200 48016 51000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 50200 48832 51000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 50200 49648 51000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 50200 27616 51000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 50200 28432 51000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 50200 29248 51000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 50200 30064 51000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 50200 30880 51000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 50200 31696 51000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 50200 32512 51000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 50200 33328 51000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 50200 1504 51000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 50200 9664 51000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 50200 10480 51000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 50200 11296 51000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 50200 12112 51000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 50200 12928 51000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 50200 13744 51000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 50200 14560 51000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 50200 15376 51000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 50200 16192 51000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 50200 17008 51000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 50200 2320 51000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 50200 17824 51000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 50200 18640 51000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 50200 19456 51000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 50200 20272 51000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 50200 21088 51000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 50200 22720 51000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 50200 23536 51000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 50200 24352 51000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 50200 25168 51000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 50200 3136 51000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 50200 3952 51000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 50200 4768 51000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 50200 5584 51000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 50200 6400 51000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 50200 7216 51000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 50200 8032 51000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 50200 8848 51000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[0]
port 66 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[10]
port 67 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[11]
port 68 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[12]
port 69 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[13]
port 70 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[14]
port 71 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[15]
port 72 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[16]
port 73 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[17]
port 74 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[18]
port 75 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[19]
port 76 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[1]
port 77 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[20]
port 78 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[21]
port 79 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[22]
port 80 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[23]
port 81 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[24]
port 82 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[25]
port 83 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[26]
port 84 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[27]
port 85 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[28]
port 86 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[29]
port 87 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[2]
port 88 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[3]
port 89 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[4]
port 90 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[5]
port 91 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[6]
port 92 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[7]
port 93 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[8]
port 94 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[9]
port 95 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[0]
port 96 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[10]
port 97 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[11]
port 98 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[12]
port 99 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[13]
port 100 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[14]
port 101 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[15]
port 102 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[16]
port 103 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[17]
port 104 nsew signal tristate
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[18]
port 105 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[19]
port 106 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[1]
port 107 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[20]
port 108 nsew signal tristate
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[21]
port 109 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[22]
port 110 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[23]
port 111 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[24]
port 112 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[25]
port 113 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[26]
port 114 nsew signal tristate
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[27]
port 115 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[28]
port 116 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[29]
port 117 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[2]
port 118 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[3]
port 119 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[4]
port 120 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[5]
port 121 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[6]
port 122 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[7]
port 123 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[8]
port 124 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 4066 56200 4122 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 6734 56200 6790 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 9402 56200 9458 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 12070 56200 12126 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 25410 56200 25466 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 28078 56200 28134 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 30746 56200 30802 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 33414 56200 33470 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 14738 56200 14794 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 17406 56200 17462 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 20074 56200 20130 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 22742 56200 22798 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 36082 56200 36138 57000 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 prog_reset_bottom_in
port 140 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 reset_bottom_in
port 141 nsew signal input
flabel metal3 s 50200 50464 51000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 142 nsew signal input
flabel metal3 s 50200 51280 51000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 143 nsew signal input
flabel metal3 s 50200 52096 51000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 144 nsew signal input
flabel metal3 s 50200 52912 51000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 145 nsew signal input
flabel metal3 s 50200 53728 51000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 146 nsew signal input
flabel metal3 s 50200 54544 51000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 147 nsew signal input
flabel metal3 s 50200 55360 51000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 148 nsew signal input
flabel metal3 s 50200 56176 51000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 149 nsew signal input
flabel metal2 s 38750 56200 38806 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 150 nsew signal input
flabel metal2 s 41418 56200 41474 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 151 nsew signal input
flabel metal2 s 44086 56200 44142 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 152 nsew signal input
flabel metal2 s 46754 56200 46810 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 154 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 test_enable_bottom_in
port 158 nsew signal input
rlabel metal1 25484 54400 25484 54400 0 VGND
rlabel metal1 25484 53856 25484 53856 0 VPWR
rlabel metal2 24242 31178 24242 31178 0 cby_0__8_.cby_0__1_.ccff_tail
rlabel metal1 22540 42194 22540 42194 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 21574 30906 21574 30906 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 21436 34170 21436 34170 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 18722 37094 18722 37094 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 24104 16422 24104 16422 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal2 13478 4624 13478 4624 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal2 23506 13226 23506 13226 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal2 23874 16150 23874 16150 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal2 25530 17102 25530 17102 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal2 32614 9350 32614 9350 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 24610 12750 24610 12750 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal2 25530 14144 25530 14144 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 27094 24242 27094 24242 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal2 32798 10642 32798 10642 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal2 33442 22950 33442 22950 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 28520 22134 28520 22134 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal2 28566 15470 28566 15470 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal2 24886 24310 24886 24310 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal2 26174 23460 26174 23460 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal2 29302 10574 29302 10574 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23322 17510 23322 17510 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 23276 30702 23276 30702 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 29578 11288 29578 11288 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 29808 12852 29808 12852 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 29118 12954 29118 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23414 12716 23414 12716 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 26312 14246 26312 14246 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 27416 12954 27416 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 23184 12954 23184 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 25898 14688 25898 14688 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 25484 14586 25484 14586 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 31556 10098 31556 10098 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24978 16048 24978 16048 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 23552 18938 23552 18938 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 31970 10064 31970 10064 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29624 12818 29624 12818 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 29854 12886 29854 12886 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26956 14858 26956 14858 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 28980 13158 28980 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 27922 12682 27922 12682 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 25024 12410 25024 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 28106 12614 28106 12614 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 26496 13498 26496 13498 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 32798 10234 32798 10234 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27094 24106 27094 24106 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 24426 24378 24426 24378 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 32154 12682 32154 12682 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29854 10438 29854 10438 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28520 11322 28520 11322 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 25622 16660 25622 16660 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 30130 14042 30130 14042 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 28474 16422 28474 16422 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 25162 16456 25162 16456 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 29854 22134 29854 22134 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 27554 24038 27554 24038 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 29072 15334 29072 15334 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24840 28118 24840 28118 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 21528 37230 21528 37230 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 28888 15402 28888 15402 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27784 10778 27784 10778 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 27186 12410 27186 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26956 17306 26956 17306 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 27416 15674 27416 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 26726 18904 26726 18904 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 24748 18394 24748 18394 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 27094 24208 27094 24208 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 24840 28050 24840 28050 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 21850 41480 21850 41480 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 24397 45458 24397 45458 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 23184 42330 23184 42330 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 26128 45254 26128 45254 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 22448 41786 22448 41786 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal2 21666 48790 21666 48790 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 21206 49130 21206 49130 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 26151 45866 26151 45866 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 19550 47498 19550 47498 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 20010 44370 20010 44370 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 20102 50218 20102 50218 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 24173 46954 24173 46954 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 17342 48212 17342 48212 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 17526 48756 17526 48756 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 22724 46478 22724 46478 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 48668 53618 48668 53618 0 ccff_head
rlabel metal2 1518 1588 1518 1588 0 ccff_head_0
rlabel metal3 49504 748 49504 748 0 ccff_tail
rlabel metal1 1748 54094 1748 54094 0 ccff_tail_0
rlabel metal2 48530 26197 48530 26197 0 chanx_right_in[0]
rlabel metal2 49358 34391 49358 34391 0 chanx_right_in[10]
rlabel via2 49358 35037 49358 35037 0 chanx_right_in[11]
rlabel metal2 49358 35989 49358 35989 0 chanx_right_in[12]
rlabel metal2 49174 36703 49174 36703 0 chanx_right_in[13]
rlabel metal2 49174 37655 49174 37655 0 chanx_right_in[14]
rlabel via2 49358 38301 49358 38301 0 chanx_right_in[15]
rlabel metal2 49358 39253 49358 39253 0 chanx_right_in[16]
rlabel metal2 49358 39967 49358 39967 0 chanx_right_in[17]
rlabel metal2 49358 40919 49358 40919 0 chanx_right_in[18]
rlabel via2 49174 41531 49174 41531 0 chanx_right_in[19]
rlabel metal2 49358 26911 49358 26911 0 chanx_right_in[1]
rlabel metal2 49174 42483 49174 42483 0 chanx_right_in[20]
rlabel metal2 49174 43231 49174 43231 0 chanx_right_in[21]
rlabel metal2 49174 44183 49174 44183 0 chanx_right_in[22]
rlabel via2 49358 44829 49358 44829 0 chanx_right_in[23]
rlabel metal2 49358 45781 49358 45781 0 chanx_right_in[24]
rlabel metal2 49358 46495 49358 46495 0 chanx_right_in[25]
rlabel metal2 49358 47447 49358 47447 0 chanx_right_in[26]
rlabel via2 49174 48059 49174 48059 0 chanx_right_in[27]
rlabel metal2 49174 49011 49174 49011 0 chanx_right_in[28]
rlabel metal2 49174 49759 49174 49759 0 chanx_right_in[29]
rlabel metal2 49358 27863 49358 27863 0 chanx_right_in[2]
rlabel via2 49358 28509 49358 28509 0 chanx_right_in[3]
rlabel metal2 49358 29461 49358 29461 0 chanx_right_in[4]
rlabel metal2 49358 30175 49358 30175 0 chanx_right_in[5]
rlabel metal2 49358 31127 49358 31127 0 chanx_right_in[6]
rlabel via2 49358 31773 49358 31773 0 chanx_right_in[7]
rlabel metal2 49358 32725 49358 32725 0 chanx_right_in[8]
rlabel metal2 49358 33439 49358 33439 0 chanx_right_in[9]
rlabel metal3 49780 1564 49780 1564 0 chanx_right_out[0]
rlabel metal3 49734 9724 49734 9724 0 chanx_right_out[10]
rlabel via2 49174 10557 49174 10557 0 chanx_right_out[11]
rlabel metal2 49174 11509 49174 11509 0 chanx_right_out[12]
rlabel metal3 49734 12172 49734 12172 0 chanx_right_out[13]
rlabel metal3 49734 12988 49734 12988 0 chanx_right_out[14]
rlabel via2 49174 13821 49174 13821 0 chanx_right_out[15]
rlabel metal2 49174 14773 49174 14773 0 chanx_right_out[16]
rlabel metal3 49734 15436 49734 15436 0 chanx_right_out[17]
rlabel metal3 49734 16252 49734 16252 0 chanx_right_out[18]
rlabel via2 49174 17085 49174 17085 0 chanx_right_out[19]
rlabel metal3 49090 2380 49090 2380 0 chanx_right_out[1]
rlabel metal2 49174 18037 49174 18037 0 chanx_right_out[20]
rlabel metal3 49734 18700 49734 18700 0 chanx_right_out[21]
rlabel metal3 49734 19516 49734 19516 0 chanx_right_out[22]
rlabel via2 49174 20349 49174 20349 0 chanx_right_out[23]
rlabel metal2 49174 21301 49174 21301 0 chanx_right_out[24]
rlabel metal3 49734 21964 49734 21964 0 chanx_right_out[25]
rlabel metal3 49734 22780 49734 22780 0 chanx_right_out[26]
rlabel via2 49174 23613 49174 23613 0 chanx_right_out[27]
rlabel metal2 49174 24565 49174 24565 0 chanx_right_out[28]
rlabel metal3 49734 25228 49734 25228 0 chanx_right_out[29]
rlabel metal2 49174 3145 49174 3145 0 chanx_right_out[2]
rlabel via2 49174 4029 49174 4029 0 chanx_right_out[3]
rlabel metal2 49174 4981 49174 4981 0 chanx_right_out[4]
rlabel metal3 49734 5644 49734 5644 0 chanx_right_out[5]
rlabel metal3 49734 6460 49734 6460 0 chanx_right_out[6]
rlabel via2 49174 7293 49174 7293 0 chanx_right_out[7]
rlabel metal2 49174 8245 49174 8245 0 chanx_right_out[8]
rlabel metal3 49734 8908 49734 8908 0 chanx_right_out[9]
rlabel metal2 2254 1860 2254 1860 0 chany_bottom_in_0[0]
rlabel metal2 9614 1554 9614 1554 0 chany_bottom_in_0[10]
rlabel metal2 10350 1588 10350 1588 0 chany_bottom_in_0[11]
rlabel metal2 11086 1894 11086 1894 0 chany_bottom_in_0[12]
rlabel metal2 11822 1588 11822 1588 0 chany_bottom_in_0[13]
rlabel metal2 12558 1860 12558 1860 0 chany_bottom_in_0[14]
rlabel metal2 13294 1622 13294 1622 0 chany_bottom_in_0[15]
rlabel metal2 14030 1860 14030 1860 0 chany_bottom_in_0[16]
rlabel metal2 14766 1588 14766 1588 0 chany_bottom_in_0[17]
rlabel metal2 15502 1588 15502 1588 0 chany_bottom_in_0[18]
rlabel metal2 16238 823 16238 823 0 chany_bottom_in_0[19]
rlabel metal2 2990 1588 2990 1588 0 chany_bottom_in_0[1]
rlabel metal2 16974 2132 16974 2132 0 chany_bottom_in_0[20]
rlabel metal2 17710 1860 17710 1860 0 chany_bottom_in_0[21]
rlabel metal2 18446 1622 18446 1622 0 chany_bottom_in_0[22]
rlabel metal2 19182 1860 19182 1860 0 chany_bottom_in_0[23]
rlabel metal2 19918 2132 19918 2132 0 chany_bottom_in_0[24]
rlabel metal2 20654 1860 20654 1860 0 chany_bottom_in_0[25]
rlabel metal2 21390 1554 21390 1554 0 chany_bottom_in_0[26]
rlabel metal1 22172 2958 22172 2958 0 chany_bottom_in_0[27]
rlabel metal2 22862 1588 22862 1588 0 chany_bottom_in_0[28]
rlabel metal2 23598 1588 23598 1588 0 chany_bottom_in_0[29]
rlabel metal2 3726 1894 3726 1894 0 chany_bottom_in_0[2]
rlabel metal2 4462 1554 4462 1554 0 chany_bottom_in_0[3]
rlabel metal2 5198 1554 5198 1554 0 chany_bottom_in_0[4]
rlabel metal2 5934 1554 5934 1554 0 chany_bottom_in_0[5]
rlabel metal2 6670 1894 6670 1894 0 chany_bottom_in_0[6]
rlabel metal2 7406 1588 7406 1588 0 chany_bottom_in_0[7]
rlabel metal2 8142 1095 8142 1095 0 chany_bottom_in_0[8]
rlabel metal2 8878 1894 8878 1894 0 chany_bottom_in_0[9]
rlabel metal1 24702 3570 24702 3570 0 chany_bottom_out_0[0]
rlabel metal2 31694 1860 31694 1860 0 chany_bottom_out_0[10]
rlabel metal1 33534 2890 33534 2890 0 chany_bottom_out_0[11]
rlabel metal2 33166 1520 33166 1520 0 chany_bottom_out_0[12]
rlabel metal1 34178 4046 34178 4046 0 chany_bottom_out_0[13]
rlabel metal1 35006 3570 35006 3570 0 chany_bottom_out_0[14]
rlabel metal2 35374 1622 35374 1622 0 chany_bottom_out_0[15]
rlabel metal1 36662 3570 36662 3570 0 chany_bottom_out_0[16]
rlabel metal1 37398 2958 37398 2958 0 chany_bottom_out_0[17]
rlabel metal1 38686 2890 38686 2890 0 chany_bottom_out_0[18]
rlabel metal2 38318 1520 38318 1520 0 chany_bottom_out_0[19]
rlabel metal1 25346 2958 25346 2958 0 chany_bottom_out_0[1]
rlabel metal1 39330 4046 39330 4046 0 chany_bottom_out_0[20]
rlabel metal1 40158 3570 40158 3570 0 chany_bottom_out_0[21]
rlabel metal2 40526 1622 40526 1622 0 chany_bottom_out_0[22]
rlabel metal2 41262 2166 41262 2166 0 chany_bottom_out_0[23]
rlabel metal1 42550 2958 42550 2958 0 chany_bottom_out_0[24]
rlabel metal1 43838 2890 43838 2890 0 chany_bottom_out_0[25]
rlabel metal2 43470 1622 43470 1622 0 chany_bottom_out_0[26]
rlabel metal1 44482 4046 44482 4046 0 chany_bottom_out_0[27]
rlabel metal1 45310 3570 45310 3570 0 chany_bottom_out_0[28]
rlabel metal1 47012 2822 47012 2822 0 chany_bottom_out_0[29]
rlabel metal2 25806 1622 25806 1622 0 chany_bottom_out_0[2]
rlabel metal2 26542 1622 26542 1622 0 chany_bottom_out_0[3]
rlabel metal1 27554 2958 27554 2958 0 chany_bottom_out_0[4]
rlabel metal2 28014 823 28014 823 0 chany_bottom_out_0[5]
rlabel metal1 29210 2958 29210 2958 0 chany_bottom_out_0[6]
rlabel metal1 29854 3434 29854 3434 0 chany_bottom_out_0[7]
rlabel metal2 30222 1588 30222 1588 0 chany_bottom_out_0[8]
rlabel metal2 30958 2166 30958 2166 0 chany_bottom_out_0[9]
rlabel metal1 34454 14994 34454 14994 0 clknet_0_prog_clk
rlabel metal1 16560 4624 16560 4624 0 clknet_4_0_0_prog_clk
rlabel metal1 22218 41650 22218 41650 0 clknet_4_10_0_prog_clk
rlabel metal1 37950 31348 37950 31348 0 clknet_4_11_0_prog_clk
rlabel metal2 40066 20060 40066 20060 0 clknet_4_12_0_prog_clk
rlabel metal2 44022 20672 44022 20672 0 clknet_4_13_0_prog_clk
rlabel metal2 40158 26180 40158 26180 0 clknet_4_14_0_prog_clk
rlabel metal1 41492 43758 41492 43758 0 clknet_4_15_0_prog_clk
rlabel metal1 25944 7922 25944 7922 0 clknet_4_1_0_prog_clk
rlabel metal1 24702 22134 24702 22134 0 clknet_4_2_0_prog_clk
rlabel metal1 29486 23766 29486 23766 0 clknet_4_3_0_prog_clk
rlabel metal2 34086 9758 34086 9758 0 clknet_4_4_0_prog_clk
rlabel metal2 35834 7684 35834 7684 0 clknet_4_5_0_prog_clk
rlabel metal1 33994 20468 33994 20468 0 clknet_4_6_0_prog_clk
rlabel metal2 39698 17238 39698 17238 0 clknet_4_7_0_prog_clk
rlabel metal1 27324 25942 27324 25942 0 clknet_4_8_0_prog_clk
rlabel metal1 34316 20978 34316 20978 0 clknet_4_9_0_prog_clk
rlabel metal1 4370 54094 4370 54094 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 6762 55209 6762 55209 0 gfpga_pad_io_soc_dir[1]
rlabel metal1 9706 54094 9706 54094 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 12282 56236 12282 56236 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 25576 54162 25576 54162 0 gfpga_pad_io_soc_in[0]
rlabel metal2 28290 56236 28290 56236 0 gfpga_pad_io_soc_in[1]
rlabel metal1 30912 54162 30912 54162 0 gfpga_pad_io_soc_in[2]
rlabel metal1 33580 54162 33580 54162 0 gfpga_pad_io_soc_in[3]
rlabel metal1 15042 54094 15042 54094 0 gfpga_pad_io_soc_out[0]
rlabel metal2 17710 56236 17710 56236 0 gfpga_pad_io_soc_out[1]
rlabel metal2 20102 55711 20102 55711 0 gfpga_pad_io_soc_out[2]
rlabel metal1 22954 54094 22954 54094 0 gfpga_pad_io_soc_out[3]
rlabel metal1 36202 54230 36202 54230 0 isol_n
rlabel metal1 42642 43826 42642 43826 0 net1
rlabel metal1 48898 39270 48898 39270 0 net10
rlabel metal1 47380 21998 47380 21998 0 net100
rlabel metal1 47978 23018 47978 23018 0 net101
rlabel metal1 47196 23698 47196 23698 0 net102
rlabel metal1 44206 22712 44206 22712 0 net103
rlabel metal1 46736 25262 46736 25262 0 net104
rlabel metal1 47150 3026 47150 3026 0 net105
rlabel metal1 47518 4114 47518 4114 0 net106
rlabel metal1 47472 5202 47472 5202 0 net107
rlabel metal1 47978 5712 47978 5712 0 net108
rlabel metal1 47518 6766 47518 6766 0 net109
rlabel metal1 49128 40154 49128 40154 0 net11
rlabel metal1 47978 7412 47978 7412 0 net110
rlabel metal1 47932 8466 47932 8466 0 net111
rlabel metal1 47978 8874 47978 8874 0 net112
rlabel metal2 37674 8806 37674 8806 0 net113
rlabel metal1 34776 12750 34776 12750 0 net114
rlabel metal1 35650 12682 35650 12682 0 net115
rlabel metal1 35696 2414 35696 2414 0 net116
rlabel metal1 34776 4114 34776 4114 0 net117
rlabel metal1 34684 3502 34684 3502 0 net118
rlabel metal1 36938 2414 36938 2414 0 net119
rlabel metal1 46046 31790 46046 31790 0 net12
rlabel metal1 37766 3502 37766 3502 0 net120
rlabel metal1 38272 3026 38272 3026 0 net121
rlabel metal1 39514 3060 39514 3060 0 net122
rlabel metal1 40158 2516 40158 2516 0 net123
rlabel metal3 37743 23596 37743 23596 0 net124
rlabel metal1 39054 4114 39054 4114 0 net125
rlabel metal2 40066 4862 40066 4862 0 net126
rlabel metal1 41538 2414 41538 2414 0 net127
rlabel metal2 40158 4624 40158 4624 0 net128
rlabel metal2 42642 4556 42642 4556 0 net129
rlabel metal1 43056 41446 43056 41446 0 net13
rlabel metal2 43378 4420 43378 4420 0 net130
rlabel metal1 44206 2414 44206 2414 0 net131
rlabel metal2 42826 4862 42826 4862 0 net132
rlabel metal2 42734 4284 42734 4284 0 net133
rlabel metal1 43976 5134 43976 5134 0 net134
rlabel metal1 31878 17272 31878 17272 0 net135
rlabel metal1 28290 2414 28290 2414 0 net136
rlabel metal2 27554 4284 27554 4284 0 net137
rlabel metal1 29532 2414 29532 2414 0 net138
rlabel metal1 29486 3026 29486 3026 0 net139
rlabel metal1 41722 22508 41722 22508 0 net14
rlabel metal2 33350 5984 33350 5984 0 net140
rlabel metal1 33166 2414 33166 2414 0 net141
rlabel metal1 35972 13226 35972 13226 0 net142
rlabel metal1 4370 54196 4370 54196 0 net143
rlabel metal1 7038 54162 7038 54162 0 net144
rlabel metal2 9614 52700 9614 52700 0 net145
rlabel metal2 12282 52836 12282 52836 0 net146
rlabel metal1 15686 51578 15686 51578 0 net147
rlabel metal2 17710 52326 17710 52326 0 net148
rlabel metal2 20286 51782 20286 51782 0 net149
rlabel metal2 35374 13736 35374 13736 0 net15
rlabel metal2 22862 51782 22862 51782 0 net150
rlabel metal2 38686 23970 38686 23970 0 net151
rlabel metal2 37766 25466 37766 25466 0 net152
rlabel metal1 42550 17170 42550 17170 0 net153
rlabel metal1 38180 26350 38180 26350 0 net154
rlabel metal1 42136 26010 42136 26010 0 net155
rlabel metal2 41722 27268 41722 27268 0 net156
rlabel metal2 40434 27846 40434 27846 0 net157
rlabel metal1 38916 28186 38916 28186 0 net158
rlabel metal1 38180 27438 38180 27438 0 net159
rlabel metal1 49588 43146 49588 43146 0 net16
rlabel metal2 40894 18394 40894 18394 0 net160
rlabel metal1 42734 16490 42734 16490 0 net161
rlabel metal1 38134 23086 38134 23086 0 net162
rlabel metal1 42550 19278 42550 19278 0 net163
rlabel metal2 21022 16966 21022 16966 0 net164
rlabel metal2 20102 13498 20102 13498 0 net165
rlabel metal1 21988 13294 21988 13294 0 net166
rlabel metal1 27186 18258 27186 18258 0 net167
rlabel metal1 28796 16558 28796 16558 0 net168
rlabel metal2 33442 17476 33442 17476 0 net169
rlabel metal1 49542 44234 49542 44234 0 net17
rlabel metal2 24978 21114 24978 21114 0 net170
rlabel metal1 33304 13294 33304 13294 0 net171
rlabel metal2 28842 9146 28842 9146 0 net172
rlabel metal2 32338 8262 32338 8262 0 net173
rlabel metal1 36064 14382 36064 14382 0 net174
rlabel metal1 30590 15130 30590 15130 0 net175
rlabel metal1 32246 16218 32246 16218 0 net176
rlabel metal1 32016 15470 32016 15470 0 net177
rlabel metal2 26450 8908 26450 8908 0 net178
rlabel metal2 32430 6766 32430 6766 0 net179
rlabel metal1 48944 44710 48944 44710 0 net18
rlabel metal2 35742 7650 35742 7650 0 net180
rlabel metal1 28198 21114 28198 21114 0 net181
rlabel metal2 37490 9112 37490 9112 0 net182
rlabel metal1 38778 11866 38778 11866 0 net183
rlabel metal1 33626 12138 33626 12138 0 net184
rlabel metal1 35972 13906 35972 13906 0 net185
rlabel metal1 35052 11866 35052 11866 0 net186
rlabel metal1 41032 11730 41032 11730 0 net187
rlabel metal2 40342 8772 40342 8772 0 net188
rlabel metal2 39054 6970 39054 6970 0 net189
rlabel metal1 49542 45798 49542 45798 0 net19
rlabel metal2 38686 9486 38686 9486 0 net190
rlabel metal1 23230 8874 23230 8874 0 net191
rlabel metal1 28520 17646 28520 17646 0 net192
rlabel metal1 25530 17306 25530 17306 0 net193
rlabel metal2 26266 14212 26266 14212 0 net194
rlabel metal2 28750 12036 28750 12036 0 net195
rlabel metal1 33764 23086 33764 23086 0 net196
rlabel metal1 31924 25874 31924 25874 0 net197
rlabel metal1 37950 21114 37950 21114 0 net198
rlabel metal1 44804 20434 44804 20434 0 net199
rlabel metal2 11730 3570 11730 3570 0 net2
rlabel metal2 41262 40188 41262 40188 0 net20
rlabel metal1 43792 20910 43792 20910 0 net200
rlabel metal2 43010 22916 43010 22916 0 net201
rlabel metal2 40342 23970 40342 23970 0 net202
rlabel metal1 47702 47430 47702 47430 0 net21
rlabel metal2 33902 35880 33902 35880 0 net22
rlabel metal1 30958 25942 30958 25942 0 net23
rlabel metal1 49450 49742 49450 49742 0 net24
rlabel metal1 43608 21522 43608 21522 0 net25
rlabel metal1 43930 23188 43930 23188 0 net26
rlabel metal1 43240 24786 43240 24786 0 net27
rlabel metal1 45264 24174 45264 24174 0 net28
rlabel metal1 47012 24106 47012 24106 0 net29
rlabel metal1 37582 12920 37582 12920 0 net3
rlabel metal1 47426 31926 47426 31926 0 net30
rlabel metal1 48300 32742 48300 32742 0 net31
rlabel metal1 48024 33286 48024 33286 0 net32
rlabel metal2 2622 5916 2622 5916 0 net33
rlabel via2 9890 2363 9890 2363 0 net34
rlabel metal2 10626 3638 10626 3638 0 net35
rlabel metal2 22034 5746 22034 5746 0 net36
rlabel metal1 17434 1836 17434 1836 0 net37
rlabel metal1 13156 3026 13156 3026 0 net38
rlabel metal1 17986 2448 17986 2448 0 net39
rlabel metal1 46690 34714 46690 34714 0 net4
rlabel metal2 14398 3332 14398 3332 0 net40
rlabel metal1 22977 2618 22977 2618 0 net41
rlabel metal2 16146 2006 16146 2006 0 net42
rlabel metal1 17112 2278 17112 2278 0 net43
rlabel metal1 20378 17102 20378 17102 0 net44
rlabel metal1 30084 7854 30084 7854 0 net45
rlabel metal2 31142 6222 31142 6222 0 net46
rlabel metal2 22310 2040 22310 2040 0 net47
rlabel metal1 19550 2924 19550 2924 0 net48
rlabel via2 20286 3587 20286 3587 0 net49
rlabel metal1 47702 17646 47702 17646 0 net5
rlabel metal2 20930 3332 20930 3332 0 net50
rlabel metal1 24886 2346 24886 2346 0 net51
rlabel metal2 33350 9401 33350 9401 0 net52
rlabel metal1 24978 2414 24978 2414 0 net53
rlabel metal2 24610 2414 24610 2414 0 net54
rlabel metal2 4002 3298 4002 3298 0 net55
rlabel metal2 4738 2108 4738 2108 0 net56
rlabel metal2 5566 2108 5566 2108 0 net57
rlabel metal2 6762 1904 6762 1904 0 net58
rlabel metal1 19412 13226 19412 13226 0 net59
rlabel metal1 46966 17714 46966 17714 0 net6
rlabel metal2 21482 13158 21482 13158 0 net60
rlabel metal2 21206 2142 21206 2142 0 net61
rlabel metal1 16560 2856 16560 2856 0 net62
rlabel metal1 23230 46580 23230 46580 0 net63
rlabel metal2 25714 50524 25714 50524 0 net64
rlabel metal1 27370 46036 27370 46036 0 net65
rlabel metal1 31556 54298 31556 54298 0 net66
rlabel metal1 21528 46682 21528 46682 0 net67
rlabel metal1 23651 41582 23651 41582 0 net68
rlabel metal1 42412 50694 42412 50694 0 net69
rlabel metal1 38088 12818 38088 12818 0 net7
rlabel metal1 49496 51306 49496 51306 0 net70
rlabel metal1 49680 52462 49680 52462 0 net71
rlabel metal1 41998 52870 41998 52870 0 net72
rlabel metal1 31326 23188 31326 23188 0 net73
rlabel metal1 49726 53414 49726 53414 0 net74
rlabel metal1 35098 29274 35098 29274 0 net75
rlabel metal1 48484 53414 48484 53414 0 net76
rlabel metal1 31418 23188 31418 23188 0 net77
rlabel metal1 33764 29206 33764 29206 0 net78
rlabel metal1 39008 21590 39008 21590 0 net79
rlabel metal1 34822 14280 34822 14280 0 net8
rlabel metal1 34178 19414 34178 19414 0 net80
rlabel metal1 45954 16966 45954 16966 0 net81
rlabel metal1 2898 54162 2898 54162 0 net82
rlabel metal2 45218 6086 45218 6086 0 net83
rlabel metal1 46460 9146 46460 9146 0 net84
rlabel metal1 45494 9146 45494 9146 0 net85
rlabel metal1 46276 11594 46276 11594 0 net86
rlabel metal1 46966 12206 46966 12206 0 net87
rlabel metal1 47932 13294 47932 13294 0 net88
rlabel metal1 47886 13906 47886 13906 0 net89
rlabel metal1 41262 30090 41262 30090 0 net9
rlabel metal1 46828 14586 46828 14586 0 net90
rlabel metal1 44620 13362 44620 13362 0 net91
rlabel metal1 43976 14042 43976 14042 0 net92
rlabel metal1 45034 15606 45034 15606 0 net93
rlabel metal2 47978 4794 47978 4794 0 net94
rlabel metal1 46506 18122 46506 18122 0 net95
rlabel metal2 47978 19108 47978 19108 0 net96
rlabel metal1 47978 19754 47978 19754 0 net97
rlabel metal1 45540 19278 45540 19278 0 net98
rlabel metal1 45080 20502 45080 20502 0 net99
rlabel metal1 31372 25194 31372 25194 0 prog_clk
rlabel metal1 47196 3434 47196 3434 0 prog_reset_bottom_in
rlabel metal2 48990 50711 48990 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 48990 51323 48990 51323 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 48990 52275 48990 52275 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 49082 53023 49082 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 49082 53975 49082 53975 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 49128 53550 49128 53550 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 49274 55420 49274 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal3 49366 56236 49366 56236 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal1 38824 54162 38824 54162 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 41492 54162 41492 54162 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 44160 54162 44160 54162 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 46828 54230 46828 54230 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 2062 1836 2062 1836 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 41262 33609 41262 33609 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 40894 33898 40894 33898 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 2062 8772 2062 8772 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 34086 16252 34086 16252 0 sb_0__8_.mem_bottom_track_1.ccff_head
rlabel metal1 40240 20026 40240 20026 0 sb_0__8_.mem_bottom_track_1.ccff_tail
rlabel metal1 38732 20366 38732 20366 0 sb_0__8_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 44068 21590 44068 21590 0 sb_0__8_.mem_bottom_track_11.ccff_head
rlabel metal1 45770 21862 45770 21862 0 sb_0__8_.mem_bottom_track_11.ccff_tail
rlabel metal1 45540 22066 45540 22066 0 sb_0__8_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 43976 24718 43976 24718 0 sb_0__8_.mem_bottom_track_13.ccff_tail
rlabel metal1 45816 23630 45816 23630 0 sb_0__8_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 43700 25806 43700 25806 0 sb_0__8_.mem_bottom_track_15.ccff_tail
rlabel metal2 45126 25330 45126 25330 0 sb_0__8_.mem_bottom_track_15.mem_out\[0\]
rlabel metal1 40664 23630 40664 23630 0 sb_0__8_.mem_bottom_track_17.ccff_tail
rlabel metal1 44206 25670 44206 25670 0 sb_0__8_.mem_bottom_track_17.mem_out\[0\]
rlabel metal1 40112 25738 40112 25738 0 sb_0__8_.mem_bottom_track_19.ccff_tail
rlabel metal2 41814 26622 41814 26622 0 sb_0__8_.mem_bottom_track_19.mem_out\[0\]
rlabel metal1 38640 28594 38640 28594 0 sb_0__8_.mem_bottom_track_29.ccff_tail
rlabel metal2 39514 28594 39514 28594 0 sb_0__8_.mem_bottom_track_29.mem_out\[0\]
rlabel metal2 42918 18462 42918 18462 0 sb_0__8_.mem_bottom_track_3.ccff_tail
rlabel metal2 41814 20706 41814 20706 0 sb_0__8_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 39606 28458 39606 28458 0 sb_0__8_.mem_bottom_track_31.ccff_tail
rlabel metal2 39974 29920 39974 29920 0 sb_0__8_.mem_bottom_track_31.mem_out\[0\]
rlabel metal1 42678 28934 42678 28934 0 sb_0__8_.mem_bottom_track_33.ccff_tail
rlabel metal2 42550 29818 42550 29818 0 sb_0__8_.mem_bottom_track_33.mem_out\[0\]
rlabel metal2 41722 29903 41722 29903 0 sb_0__8_.mem_bottom_track_35.ccff_tail
rlabel metal1 43608 31858 43608 31858 0 sb_0__8_.mem_bottom_track_35.mem_out\[0\]
rlabel metal2 40342 29546 40342 29546 0 sb_0__8_.mem_bottom_track_45.ccff_tail
rlabel metal1 43424 33422 43424 33422 0 sb_0__8_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 39284 32198 39284 32198 0 sb_0__8_.mem_bottom_track_47.ccff_tail
rlabel metal1 41814 31892 41814 31892 0 sb_0__8_.mem_bottom_track_47.mem_out\[0\]
rlabel metal1 40112 26282 40112 26282 0 sb_0__8_.mem_bottom_track_49.ccff_tail
rlabel metal2 39698 30634 39698 30634 0 sb_0__8_.mem_bottom_track_49.mem_out\[0\]
rlabel metal2 40526 20264 40526 20264 0 sb_0__8_.mem_bottom_track_5.ccff_tail
rlabel metal1 43463 20026 43463 20026 0 sb_0__8_.mem_bottom_track_5.mem_out\[0\]
rlabel metal2 44114 27149 44114 27149 0 sb_0__8_.mem_bottom_track_51.mem_out\[0\]
rlabel metal1 40112 22542 40112 22542 0 sb_0__8_.mem_bottom_track_7.ccff_tail
rlabel metal2 39330 22338 39330 22338 0 sb_0__8_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 42550 23222 42550 23222 0 sb_0__8_.mem_bottom_track_9.mem_out\[0\]
rlabel metal1 28888 25670 28888 25670 0 sb_0__8_.mem_right_track_0.ccff_tail
rlabel metal1 39146 43622 39146 43622 0 sb_0__8_.mem_right_track_0.mem_out\[0\]
rlabel metal1 26956 25806 26956 25806 0 sb_0__8_.mem_right_track_0.mem_out\[1\]
rlabel metal2 31234 23936 31234 23936 0 sb_0__8_.mem_right_track_10.ccff_head
rlabel metal1 25898 20230 25898 20230 0 sb_0__8_.mem_right_track_10.ccff_tail
rlabel metal1 30452 24038 30452 24038 0 sb_0__8_.mem_right_track_10.mem_out\[0\]
rlabel metal1 24978 23290 24978 23290 0 sb_0__8_.mem_right_track_10.mem_out\[1\]
rlabel metal1 28842 20570 28842 20570 0 sb_0__8_.mem_right_track_12.ccff_tail
rlabel metal1 21666 13396 21666 13396 0 sb_0__8_.mem_right_track_12.mem_out\[0\]
rlabel metal1 33166 21420 33166 21420 0 sb_0__8_.mem_right_track_14.ccff_tail
rlabel metal2 34546 23766 34546 23766 0 sb_0__8_.mem_right_track_14.mem_out\[0\]
rlabel metal2 31786 20774 31786 20774 0 sb_0__8_.mem_right_track_16.ccff_tail
rlabel metal1 32614 21114 32614 21114 0 sb_0__8_.mem_right_track_16.mem_out\[0\]
rlabel metal1 31878 16558 31878 16558 0 sb_0__8_.mem_right_track_18.ccff_tail
rlabel metal1 30360 18326 30360 18326 0 sb_0__8_.mem_right_track_18.mem_out\[0\]
rlabel metal1 30636 25398 30636 25398 0 sb_0__8_.mem_right_track_2.ccff_tail
rlabel metal2 30314 27472 30314 27472 0 sb_0__8_.mem_right_track_2.mem_out\[0\]
rlabel metal1 29394 26758 29394 26758 0 sb_0__8_.mem_right_track_2.mem_out\[1\]
rlabel metal2 29486 11900 29486 11900 0 sb_0__8_.mem_right_track_20.ccff_tail
rlabel metal1 29624 13362 29624 13362 0 sb_0__8_.mem_right_track_20.mem_out\[0\]
rlabel metal1 27370 9078 27370 9078 0 sb_0__8_.mem_right_track_22.ccff_tail
rlabel metal1 26588 9010 26588 9010 0 sb_0__8_.mem_right_track_22.mem_out\[0\]
rlabel metal1 30452 8398 30452 8398 0 sb_0__8_.mem_right_track_24.ccff_tail
rlabel metal1 27774 8262 27774 8262 0 sb_0__8_.mem_right_track_24.mem_out\[0\]
rlabel metal1 34730 14042 34730 14042 0 sb_0__8_.mem_right_track_26.ccff_tail
rlabel metal2 32430 13532 32430 13532 0 sb_0__8_.mem_right_track_26.mem_out\[0\]
rlabel metal1 35006 19686 35006 19686 0 sb_0__8_.mem_right_track_28.ccff_tail
rlabel metal1 33849 20026 33849 20026 0 sb_0__8_.mem_right_track_28.mem_out\[0\]
rlabel metal2 36570 21148 36570 21148 0 sb_0__8_.mem_right_track_30.ccff_tail
rlabel metal1 35604 20230 35604 20230 0 sb_0__8_.mem_right_track_30.mem_out\[0\]
rlabel metal2 34362 17612 34362 17612 0 sb_0__8_.mem_right_track_32.ccff_tail
rlabel metal1 36892 21114 36892 21114 0 sb_0__8_.mem_right_track_32.mem_out\[0\]
rlabel metal2 31786 12517 31786 12517 0 sb_0__8_.mem_right_track_34.ccff_tail
rlabel metal1 33810 16422 33810 16422 0 sb_0__8_.mem_right_track_34.mem_out\[0\]
rlabel metal2 32246 6222 32246 6222 0 sb_0__8_.mem_right_track_36.ccff_tail
rlabel metal1 30767 6970 30767 6970 0 sb_0__8_.mem_right_track_36.mem_out\[0\]
rlabel metal1 33948 7310 33948 7310 0 sb_0__8_.mem_right_track_38.ccff_tail
rlabel metal2 32614 7140 32614 7140 0 sb_0__8_.mem_right_track_38.mem_out\[0\]
rlabel metal1 33258 26418 33258 26418 0 sb_0__8_.mem_right_track_4.ccff_tail
rlabel metal2 32062 28016 32062 28016 0 sb_0__8_.mem_right_track_4.mem_out\[0\]
rlabel metal1 30774 26418 30774 26418 0 sb_0__8_.mem_right_track_4.mem_out\[1\]
rlabel metal1 35788 8602 35788 8602 0 sb_0__8_.mem_right_track_40.ccff_tail
rlabel metal1 34454 8534 34454 8534 0 sb_0__8_.mem_right_track_40.mem_out\[0\]
rlabel metal1 37260 13158 37260 13158 0 sb_0__8_.mem_right_track_42.ccff_tail
rlabel metal1 36616 12138 36616 12138 0 sb_0__8_.mem_right_track_42.mem_out\[0\]
rlabel metal1 37582 15674 37582 15674 0 sb_0__8_.mem_right_track_44.ccff_tail
rlabel metal2 36064 15538 36064 15538 0 sb_0__8_.mem_right_track_44.mem_out\[0\]
rlabel metal2 39974 16864 39974 16864 0 sb_0__8_.mem_right_track_46.ccff_tail
rlabel metal1 37720 18326 37720 18326 0 sb_0__8_.mem_right_track_46.mem_out\[0\]
rlabel metal2 39422 14620 39422 14620 0 sb_0__8_.mem_right_track_48.ccff_tail
rlabel metal2 39054 18258 39054 18258 0 sb_0__8_.mem_right_track_48.mem_out\[0\]
rlabel metal1 40848 12614 40848 12614 0 sb_0__8_.mem_right_track_50.ccff_tail
rlabel metal1 40158 12750 40158 12750 0 sb_0__8_.mem_right_track_50.mem_out\[0\]
rlabel metal1 40526 8432 40526 8432 0 sb_0__8_.mem_right_track_52.ccff_tail
rlabel metal2 38778 10064 38778 10064 0 sb_0__8_.mem_right_track_52.mem_out\[0\]
rlabel metal1 37996 6834 37996 6834 0 sb_0__8_.mem_right_track_54.ccff_tail
rlabel metal1 36606 6970 36606 6970 0 sb_0__8_.mem_right_track_54.mem_out\[0\]
rlabel metal1 35052 8806 35052 8806 0 sb_0__8_.mem_right_track_56.ccff_tail
rlabel metal2 35190 8466 35190 8466 0 sb_0__8_.mem_right_track_56.mem_out\[0\]
rlabel metal1 33258 14926 33258 14926 0 sb_0__8_.mem_right_track_58.mem_out\[0\]
rlabel metal1 33994 23630 33994 23630 0 sb_0__8_.mem_right_track_6.ccff_tail
rlabel metal2 35006 26826 35006 26826 0 sb_0__8_.mem_right_track_6.mem_out\[0\]
rlabel metal1 32338 23766 32338 23766 0 sb_0__8_.mem_right_track_6.mem_out\[1\]
rlabel metal1 33902 24582 33902 24582 0 sb_0__8_.mem_right_track_8.mem_out\[0\]
rlabel metal1 29624 23630 29624 23630 0 sb_0__8_.mem_right_track_8.mem_out\[1\]
rlabel metal2 36570 9588 36570 9588 0 sb_0__8_.mux_bottom_track_1.out
rlabel metal1 39330 19822 39330 19822 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 38870 20604 38870 20604 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36478 15062 36478 15062 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40710 14246 40710 14246 0 sb_0__8_.mux_bottom_track_11.out
rlabel metal1 44804 20570 44804 20570 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 41170 14348 41170 14348 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37950 15402 37950 15402 0 sb_0__8_.mux_bottom_track_13.out
rlabel metal1 43746 20842 43746 20842 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 43654 18258 43654 18258 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38548 15878 38548 15878 0 sb_0__8_.mux_bottom_track_15.out
rlabel metal1 43378 22746 43378 22746 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 39468 19108 39468 19108 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37536 15878 37536 15878 0 sb_0__8_.mux_bottom_track_17.out
rlabel metal1 40480 23766 40480 23766 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37628 16082 37628 16082 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35466 16422 35466 16422 0 sb_0__8_.mux_bottom_track_19.out
rlabel metal1 39330 23766 39330 23766 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36248 16490 36248 16490 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34638 6766 34638 6766 0 sb_0__8_.mux_bottom_track_29.out
rlabel metal1 39238 25194 39238 25194 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36478 17714 36478 17714 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 40480 12070 40480 12070 0 sb_0__8_.mux_bottom_track_3.out
rlabel metal1 43010 17238 43010 17238 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40664 12206 40664 12206 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33580 18054 33580 18054 0 sb_0__8_.mux_bottom_track_31.out
rlabel metal1 38502 26418 38502 26418 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35374 18258 35374 18258 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38410 9486 38410 9486 0 sb_0__8_.mux_bottom_track_33.out
rlabel metal1 41814 25738 41814 25738 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40296 16558 40296 16558 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 39054 18394 39054 18394 0 sb_0__8_.mux_bottom_track_35.out
rlabel metal1 42596 31926 42596 31926 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40526 18258 40526 18258 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35006 18734 35006 18734 0 sb_0__8_.mux_bottom_track_45.out
rlabel metal2 40250 30736 40250 30736 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37628 18734 37628 18734 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35926 18598 35926 18598 0 sb_0__8_.mux_bottom_track_47.out
rlabel metal1 38456 28050 38456 28050 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36984 18802 36984 18802 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32154 19006 32154 19006 0 sb_0__8_.mux_bottom_track_49.out
rlabel metal1 39376 27370 39376 27370 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32384 22950 32384 22950 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 39284 13158 39284 13158 0 sb_0__8_.mux_bottom_track_5.out
rlabel metal1 40940 18802 40940 18802 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 39514 15946 39514 15946 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34822 12682 34822 12682 0 sb_0__8_.mux_bottom_track_51.out
rlabel metal1 42688 16626 42688 16626 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40250 14518 40250 14518 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36662 16626 36662 16626 0 sb_0__8_.mux_bottom_track_7.out
rlabel metal2 39238 23324 39238 23324 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38640 23222 38640 23222 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37996 21862 37996 21862 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40296 13158 40296 13158 0 sb_0__8_.mux_bottom_track_9.out
rlabel metal1 43240 19346 43240 19346 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40250 13328 40250 13328 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 43378 25160 43378 25160 0 sb_0__8_.mux_right_track_0.out
rlabel metal2 31510 29682 31510 29682 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33166 27948 33166 27948 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29394 27846 29394 27846 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20378 17272 20378 17272 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36294 24276 36294 24276 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37444 20026 37444 20026 0 sb_0__8_.mux_right_track_10.out
rlabel metal1 30682 23086 30682 23086 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30636 26826 30636 26826 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28520 22950 28520 22950 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20056 13498 20056 13498 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 35098 19380 35098 19380 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 36478 19720 36478 19720 0 sb_0__8_.mux_right_track_12.out
rlabel metal1 30544 22950 30544 22950 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 13362 21022 13362 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36662 19856 36662 19856 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 42826 20808 42826 20808 0 sb_0__8_.mux_right_track_14.out
rlabel metal1 32936 21658 32936 21658 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28934 18054 28934 18054 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38870 20978 38870 20978 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 41216 19482 41216 19482 0 sb_0__8_.mux_right_track_16.out
rlabel metal1 33626 20910 33626 20910 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32430 20808 32430 20808 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36754 19346 36754 19346 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43470 18020 43470 18020 0 sb_0__8_.mux_right_track_18.out
rlabel metal1 31234 17034 31234 17034 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33074 17272 33074 17272 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 36754 25024 36754 25024 0 sb_0__8_.mux_right_track_2.out
rlabel metal1 31556 27098 31556 27098 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 31418 28186 31418 28186 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30866 26758 30866 26758 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 26036 21114 26036 21114 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30222 25194 30222 25194 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38180 15130 38180 15130 0 sb_0__8_.mux_right_track_20.out
rlabel metal1 32798 13226 32798 13226 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34960 13498 34960 13498 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36984 11866 36984 11866 0 sb_0__8_.mux_right_track_22.out
rlabel metal2 23506 8704 23506 8704 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 36294 11747 36294 11747 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 44344 13294 44344 13294 0 sb_0__8_.mux_right_track_24.out
rlabel metal1 26956 8602 26956 8602 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33994 8466 33994 8466 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 43654 14280 43654 14280 0 sb_0__8_.mux_right_track_26.out
rlabel metal1 33718 13430 33718 13430 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 41262 14450 41262 14450 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 42550 16558 42550 16558 0 sb_0__8_.mux_right_track_28.out
rlabel metal1 35328 18802 35328 18802 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32338 16626 32338 16626 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 40480 17646 40480 17646 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43562 16252 43562 16252 0 sb_0__8_.mux_right_track_30.out
rlabel metal1 36432 24582 36432 24582 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33580 15878 33580 15878 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel viali 41262 17644 41262 17644 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 42734 14926 42734 14926 0 sb_0__8_.mux_right_track_32.out
rlabel metal1 35880 23494 35880 23494 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 31372 15674 31372 15674 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 40802 17136 40802 17136 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 38502 11934 38502 11934 0 sb_0__8_.mux_right_track_34.out
rlabel metal1 32890 19210 32890 19210 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26128 8262 26128 8262 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38686 12240 38686 12240 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 45310 8432 45310 8432 0 sb_0__8_.mux_right_track_36.out
rlabel metal2 30038 6800 30038 6800 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32752 5882 32752 5882 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 44206 8500 44206 8500 0 sb_0__8_.mux_right_track_38.out
rlabel metal1 35696 7378 35696 7378 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37812 7242 37812 7242 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 38410 24446 38410 24446 0 sb_0__8_.mux_right_track_4.out
rlabel metal1 34178 27302 34178 27302 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33396 27438 33396 27438 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33718 25330 33718 25330 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 30544 25194 30544 25194 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 38594 25092 38594 25092 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 46874 9010 46874 9010 0 sb_0__8_.mux_right_track_40.out
rlabel metal1 35190 9010 35190 9010 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 37306 8942 37306 8942 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 45310 9554 45310 9554 0 sb_0__8_.mux_right_track_42.out
rlabel metal2 38318 11934 38318 11934 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39606 11560 39606 11560 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 42872 12614 42872 12614 0 sb_0__8_.mux_right_track_44.out
rlabel metal1 36754 21862 36754 21862 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33672 15402 33672 15402 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 40894 14212 40894 14212 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 43470 13430 43470 13430 0 sb_0__8_.mux_right_track_46.out
rlabel metal1 37996 22406 37996 22406 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35098 13838 35098 13838 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 40526 14892 40526 14892 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 45954 8534 45954 8534 0 sb_0__8_.mux_right_track_48.out
rlabel metal2 39238 17884 39238 17884 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39008 14246 39008 14246 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 38778 14144 38778 14144 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 46322 7378 46322 7378 0 sb_0__8_.mux_right_track_50.out
rlabel metal2 40664 12716 40664 12716 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40779 11594 40779 11594 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 46184 5678 46184 5678 0 sb_0__8_.mux_right_track_52.out
rlabel metal1 40296 8534 40296 8534 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 41262 7854 41262 7854 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 46000 4114 46000 4114 0 sb_0__8_.mux_right_track_54.out
rlabel metal2 39146 8058 39146 8058 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40618 6154 40618 6154 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 45172 5202 45172 5202 0 sb_0__8_.mux_right_track_56.out
rlabel metal1 38870 8942 38870 8942 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40066 7922 40066 7922 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 40434 7820 40434 7820 0 sb_0__8_.mux_right_track_58.out
rlabel metal2 32798 16150 32798 16150 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32223 12818 32223 12818 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32292 11356 32292 11356 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 42182 22984 42182 22984 0 sb_0__8_.mux_right_track_6.out
rlabel metal2 35834 27506 35834 27506 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35650 26010 35650 26010 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34638 22746 34638 22746 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33350 17663 33350 17663 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 33488 22474 33488 22474 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37720 22066 37720 22066 0 sb_0__8_.mux_right_track_8.out
rlabel metal2 31510 25670 31510 25670 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32706 25874 32706 25874 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31096 21658 31096 21658 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25116 17306 25116 17306 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30774 21658 30774 21658 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
<< properties >>
string FIXED_BBOX 0 0 51000 57000
<< end >>
