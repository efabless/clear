magic
tech sky130A
magscale 1 2
timestamp 1679321909
<< viali >>
rect 31585 54281 31619 54315
rect 41521 54281 41555 54315
rect 3249 54213 3283 54247
rect 5825 54213 5859 54247
rect 8401 54213 8435 54247
rect 10977 54213 11011 54247
rect 13553 54213 13587 54247
rect 16129 54213 16163 54247
rect 18705 54213 18739 54247
rect 21005 54213 21039 54247
rect 24869 54213 24903 54247
rect 28733 54213 28767 54247
rect 32965 54213 32999 54247
rect 33701 54213 33735 54247
rect 37565 54213 37599 54247
rect 42717 54213 42751 54247
rect 2237 54145 2271 54179
rect 4169 54145 4203 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9781 54145 9815 54179
rect 12541 54145 12575 54179
rect 15117 54145 15151 54179
rect 17693 54145 17727 54179
rect 20269 54145 20303 54179
rect 22753 54145 22787 54179
rect 25513 54145 25547 54179
rect 26433 54145 26467 54179
rect 27169 54145 27203 54179
rect 27905 54145 27939 54179
rect 29929 54145 29963 54179
rect 30665 54145 30699 54179
rect 31401 54145 31435 54179
rect 34897 54145 34931 54179
rect 35817 54145 35851 54179
rect 36553 54145 36587 54179
rect 38761 54145 38795 54179
rect 40049 54145 40083 54179
rect 40785 54145 40819 54179
rect 41705 54145 41739 54179
rect 43729 54145 43763 54179
rect 44373 54145 44407 54179
rect 45385 54145 45419 54179
rect 47961 54145 47995 54179
rect 23029 54077 23063 54111
rect 42993 54077 43027 54111
rect 48421 54077 48455 54111
rect 25053 54009 25087 54043
rect 28917 54009 28951 54043
rect 33149 54009 33183 54043
rect 33885 54009 33919 54043
rect 44189 54009 44223 54043
rect 3985 53941 4019 53975
rect 25697 53941 25731 53975
rect 26249 53941 26283 53975
rect 27353 53941 27387 53975
rect 28089 53941 28123 53975
rect 30113 53941 30147 53975
rect 30849 53941 30883 53975
rect 35081 53941 35115 53975
rect 36001 53941 36035 53975
rect 36737 53941 36771 53975
rect 37657 53941 37691 53975
rect 38945 53941 38979 53975
rect 40233 53941 40267 53975
rect 40969 53941 41003 53975
rect 43545 53941 43579 53975
rect 45201 53941 45235 53975
rect 23673 53669 23707 53703
rect 2421 53601 2455 53635
rect 5733 53601 5767 53635
rect 7573 53601 7607 53635
rect 10885 53601 10919 53635
rect 12725 53601 12759 53635
rect 16129 53601 16163 53635
rect 18337 53601 18371 53635
rect 20453 53601 20487 53635
rect 22293 53601 22327 53635
rect 47317 53601 47351 53635
rect 2145 53533 2179 53567
rect 5457 53533 5491 53567
rect 7297 53533 7331 53567
rect 10425 53533 10459 53567
rect 12357 53533 12391 53567
rect 15853 53533 15887 53567
rect 17693 53533 17727 53567
rect 20177 53533 20211 53567
rect 22017 53533 22051 53567
rect 23857 53533 23891 53567
rect 24685 53533 24719 53567
rect 29929 53533 29963 53567
rect 32321 53533 32355 53567
rect 35265 53533 35299 53567
rect 38209 53533 38243 53567
rect 41889 53533 41923 53567
rect 46857 53533 46891 53567
rect 24869 53465 24903 53499
rect 29745 53397 29779 53431
rect 32137 53397 32171 53431
rect 35081 53397 35115 53431
rect 38025 53397 38059 53431
rect 41705 53397 41739 53431
rect 46213 53193 46247 53227
rect 49157 53125 49191 53159
rect 1685 53057 1719 53091
rect 2881 53057 2915 53091
rect 4813 53057 4847 53091
rect 8033 53057 8067 53091
rect 9781 53057 9815 53091
rect 13185 53057 13219 53091
rect 15025 53057 15059 53091
rect 17601 53057 17635 53091
rect 19625 53057 19659 53091
rect 46397 53057 46431 53091
rect 47961 53057 47995 53091
rect 3157 52989 3191 53023
rect 5089 52989 5123 53023
rect 8309 52989 8343 53023
rect 10241 52989 10275 53023
rect 13461 52989 13495 53023
rect 15393 52989 15427 53023
rect 17877 52989 17911 53023
rect 20085 52989 20119 53023
rect 1869 52921 1903 52955
rect 2053 52513 2087 52547
rect 4629 52513 4663 52547
rect 9781 52513 9815 52547
rect 14933 52513 14967 52547
rect 1777 52445 1811 52479
rect 4353 52445 4387 52479
rect 9505 52445 9539 52479
rect 14657 52445 14691 52479
rect 23581 52105 23615 52139
rect 2789 52037 2823 52071
rect 1593 51969 1627 52003
rect 23765 51969 23799 52003
rect 49065 51969 49099 52003
rect 49249 51765 49283 51799
rect 13093 51561 13127 51595
rect 14473 51561 14507 51595
rect 24685 51561 24719 51595
rect 24869 51357 24903 51391
rect 49065 51357 49099 51391
rect 13001 51289 13035 51323
rect 14381 51289 14415 51323
rect 49249 51221 49283 51255
rect 22201 51017 22235 51051
rect 23305 50949 23339 50983
rect 1685 50881 1719 50915
rect 22109 50881 22143 50915
rect 23121 50881 23155 50915
rect 48973 50881 49007 50915
rect 1777 50677 1811 50711
rect 49249 50677 49283 50711
rect 20269 50473 20303 50507
rect 49065 50269 49099 50303
rect 20177 50201 20211 50235
rect 49249 50133 49283 50167
rect 12357 49929 12391 49963
rect 14749 49929 14783 49963
rect 12265 49861 12299 49895
rect 14657 49793 14691 49827
rect 18153 49385 18187 49419
rect 20361 49385 20395 49419
rect 18061 49181 18095 49215
rect 49065 49181 49099 49215
rect 20269 49113 20303 49147
rect 49249 49045 49283 49079
rect 49065 48705 49099 48739
rect 49249 48501 49283 48535
rect 10149 48161 10183 48195
rect 49065 48093 49099 48127
rect 1685 48025 1719 48059
rect 1869 48025 1903 48059
rect 10425 48025 10459 48059
rect 12173 48025 12207 48059
rect 49249 47957 49283 47991
rect 24593 47753 24627 47787
rect 24777 47617 24811 47651
rect 49065 47617 49099 47651
rect 49249 47413 49283 47447
rect 18429 46121 18463 46155
rect 26709 46121 26743 46155
rect 18613 45917 18647 45951
rect 19717 45917 19751 45951
rect 26893 45917 26927 45951
rect 48145 45917 48179 45951
rect 1685 45849 1719 45883
rect 49157 45849 49191 45883
rect 1777 45781 1811 45815
rect 19533 45781 19567 45815
rect 48605 45577 48639 45611
rect 15117 45509 15151 45543
rect 33885 45509 33919 45543
rect 14933 45441 14967 45475
rect 32689 45441 32723 45475
rect 32781 45441 32815 45475
rect 48145 45441 48179 45475
rect 48789 45441 48823 45475
rect 32873 45373 32907 45407
rect 33977 45373 34011 45407
rect 34161 45373 34195 45407
rect 32321 45237 32355 45271
rect 33517 45237 33551 45271
rect 47961 45237 47995 45271
rect 22937 45033 22971 45067
rect 25053 45033 25087 45067
rect 34897 44965 34931 44999
rect 35357 44897 35391 44931
rect 35541 44897 35575 44931
rect 48789 44897 48823 44931
rect 23121 44829 23155 44863
rect 25237 44829 25271 44863
rect 48513 44829 48547 44863
rect 35265 44693 35299 44727
rect 14381 44489 14415 44523
rect 36645 44489 36679 44523
rect 39221 44489 39255 44523
rect 14289 44353 14323 44387
rect 36553 44353 36587 44387
rect 39129 44353 39163 44387
rect 36829 44285 36863 44319
rect 39313 44285 39347 44319
rect 36185 44149 36219 44183
rect 38761 44149 38795 44183
rect 13553 43945 13587 43979
rect 16221 43945 16255 43979
rect 16957 43945 16991 43979
rect 20453 43945 20487 43979
rect 21281 43945 21315 43979
rect 21833 43945 21867 43979
rect 28457 43945 28491 43979
rect 12357 43877 12391 43911
rect 22937 43877 22971 43911
rect 29009 43809 29043 43843
rect 30297 43809 30331 43843
rect 33977 43809 34011 43843
rect 37749 43809 37783 43843
rect 37933 43809 37967 43843
rect 48789 43809 48823 43843
rect 19809 43741 19843 43775
rect 20361 43741 20395 43775
rect 22017 43741 22051 43775
rect 30021 43741 30055 43775
rect 32229 43741 32263 43775
rect 48513 43741 48547 43775
rect 12173 43673 12207 43707
rect 13461 43673 13495 43707
rect 15577 43673 15611 43707
rect 16129 43673 16163 43707
rect 16865 43673 16899 43707
rect 21189 43673 21223 43707
rect 22753 43673 22787 43707
rect 28825 43673 28859 43707
rect 32505 43673 32539 43707
rect 37657 43673 37691 43707
rect 28917 43605 28951 43639
rect 31769 43605 31803 43639
rect 37289 43605 37323 43639
rect 16865 43401 16899 43435
rect 19165 43401 19199 43435
rect 20361 43401 20395 43435
rect 20913 43401 20947 43435
rect 25881 43401 25915 43435
rect 40325 43401 40359 43435
rect 34805 43333 34839 43367
rect 12081 43265 12115 43299
rect 17049 43265 17083 43299
rect 19073 43265 19107 43299
rect 20269 43265 20303 43299
rect 21097 43265 21131 43299
rect 26249 43265 26283 43299
rect 32321 43265 32355 43299
rect 34529 43265 34563 43299
rect 40233 43265 40267 43299
rect 48789 43265 48823 43299
rect 12265 43197 12299 43231
rect 26341 43197 26375 43231
rect 26525 43197 26559 43231
rect 28825 43197 28859 43231
rect 29101 43197 29135 43231
rect 40509 43197 40543 43231
rect 48513 43197 48547 43231
rect 30573 43061 30607 43095
rect 32584 43061 32618 43095
rect 34069 43061 34103 43095
rect 36277 43061 36311 43095
rect 39865 43061 39899 43095
rect 27353 42857 27387 42891
rect 9413 42721 9447 42755
rect 17417 42721 17451 42755
rect 35909 42721 35943 42755
rect 40693 42721 40727 42755
rect 25605 42653 25639 42687
rect 35633 42653 35667 42687
rect 40509 42653 40543 42687
rect 48513 42653 48547 42687
rect 48789 42653 48823 42687
rect 9229 42585 9263 42619
rect 17233 42585 17267 42619
rect 25881 42585 25915 42619
rect 37381 42517 37415 42551
rect 40049 42517 40083 42551
rect 40417 42517 40451 42551
rect 7205 42313 7239 42347
rect 20729 42313 20763 42347
rect 22109 42313 22143 42347
rect 40049 42313 40083 42347
rect 41705 42313 41739 42347
rect 8033 42245 8067 42279
rect 27997 42245 28031 42279
rect 30297 42245 30331 42279
rect 7113 42177 7147 42211
rect 7849 42177 7883 42211
rect 20913 42177 20947 42211
rect 22293 42177 22327 42211
rect 24133 42177 24167 42211
rect 33885 42177 33919 42211
rect 41613 42177 41647 42211
rect 24409 42109 24443 42143
rect 27721 42109 27755 42143
rect 30021 42109 30055 42143
rect 34161 42109 34195 42143
rect 38301 42109 38335 42143
rect 38577 42109 38611 42143
rect 41889 42109 41923 42143
rect 48513 42109 48547 42143
rect 48789 42109 48823 42143
rect 25881 41973 25915 42007
rect 29469 41973 29503 42007
rect 31769 41973 31803 42007
rect 35633 41973 35667 42007
rect 41245 41973 41279 42007
rect 26985 41769 27019 41803
rect 36645 41769 36679 41803
rect 38853 41769 38887 41803
rect 21649 41633 21683 41667
rect 23673 41633 23707 41667
rect 27445 41633 27479 41667
rect 27537 41633 27571 41667
rect 34897 41633 34931 41667
rect 37105 41633 37139 41667
rect 31401 41565 31435 41599
rect 1685 41497 1719 41531
rect 21189 41497 21223 41531
rect 21925 41497 21959 41531
rect 31677 41497 31711 41531
rect 35173 41497 35207 41531
rect 37381 41497 37415 41531
rect 1777 41429 1811 41463
rect 27353 41429 27387 41463
rect 33149 41429 33183 41463
rect 5825 41225 5859 41259
rect 9873 41225 9907 41259
rect 10793 41225 10827 41259
rect 22017 41225 22051 41259
rect 29469 41225 29503 41259
rect 21189 41157 21223 41191
rect 22385 41157 22419 41191
rect 29837 41157 29871 41191
rect 33425 41157 33459 41191
rect 5733 41089 5767 41123
rect 9781 41089 9815 41123
rect 10701 41089 10735 41123
rect 27261 41089 27295 41123
rect 29929 41089 29963 41123
rect 38209 41089 38243 41123
rect 22477 41021 22511 41055
rect 22661 41021 22695 41055
rect 24777 41021 24811 41055
rect 25053 41021 25087 41055
rect 27537 41021 27571 41055
rect 30021 41021 30055 41055
rect 33149 41021 33183 41055
rect 38485 41021 38519 41055
rect 48513 41021 48547 41055
rect 48789 41021 48823 41055
rect 26525 40953 26559 40987
rect 23305 40885 23339 40919
rect 29009 40885 29043 40919
rect 34897 40885 34931 40919
rect 39957 40885 39991 40919
rect 25513 40681 25547 40715
rect 23213 40613 23247 40647
rect 35265 40613 35299 40647
rect 23857 40545 23891 40579
rect 26157 40545 26191 40579
rect 27353 40545 27387 40579
rect 31493 40545 31527 40579
rect 32689 40545 32723 40579
rect 32781 40545 32815 40579
rect 34069 40545 34103 40579
rect 34161 40545 34195 40579
rect 35817 40545 35851 40579
rect 39221 40545 39255 40579
rect 39405 40545 39439 40579
rect 48789 40545 48823 40579
rect 23673 40477 23707 40511
rect 27077 40477 27111 40511
rect 27169 40477 27203 40511
rect 29745 40477 29779 40511
rect 32597 40477 32631 40511
rect 48513 40477 48547 40511
rect 25881 40409 25915 40443
rect 25973 40409 26007 40443
rect 30021 40409 30055 40443
rect 35633 40409 35667 40443
rect 23581 40341 23615 40375
rect 26709 40341 26743 40375
rect 32229 40341 32263 40375
rect 33609 40341 33643 40375
rect 33977 40341 34011 40375
rect 35725 40341 35759 40375
rect 38761 40341 38795 40375
rect 39129 40341 39163 40375
rect 24961 40137 24995 40171
rect 34069 40137 34103 40171
rect 36461 40137 36495 40171
rect 40325 40137 40359 40171
rect 40785 40137 40819 40171
rect 38853 40069 38887 40103
rect 41153 40069 41187 40103
rect 23213 40001 23247 40035
rect 34713 40001 34747 40035
rect 38577 40001 38611 40035
rect 41245 40001 41279 40035
rect 23489 39933 23523 39967
rect 28181 39933 28215 39967
rect 28457 39933 28491 39967
rect 32321 39933 32355 39967
rect 32597 39933 32631 39967
rect 34989 39933 35023 39967
rect 41429 39933 41463 39967
rect 48513 39933 48547 39967
rect 48789 39933 48823 39967
rect 29929 39797 29963 39831
rect 32689 39593 32723 39627
rect 38761 39593 38795 39627
rect 22017 39525 22051 39559
rect 31953 39525 31987 39559
rect 22569 39457 22603 39491
rect 24593 39457 24627 39491
rect 24869 39457 24903 39491
rect 30205 39457 30239 39491
rect 33241 39457 33275 39491
rect 34253 39457 34287 39491
rect 36277 39457 36311 39491
rect 39221 39457 39255 39491
rect 39313 39457 39347 39491
rect 41245 39457 41279 39491
rect 48789 39457 48823 39491
rect 22385 39389 22419 39423
rect 33057 39389 33091 39423
rect 36001 39389 36035 39423
rect 40969 39389 41003 39423
rect 48513 39389 48547 39423
rect 30481 39321 30515 39355
rect 34069 39321 34103 39355
rect 35357 39321 35391 39355
rect 21465 39253 21499 39287
rect 22477 39253 22511 39287
rect 26341 39253 26375 39287
rect 33149 39253 33183 39287
rect 33609 39253 33643 39287
rect 33977 39253 34011 39287
rect 37749 39253 37783 39287
rect 39129 39253 39163 39287
rect 42717 39253 42751 39287
rect 22385 39049 22419 39083
rect 23213 39049 23247 39083
rect 24501 39049 24535 39083
rect 25881 39049 25915 39083
rect 27353 39049 27387 39083
rect 28917 39049 28951 39083
rect 34161 39049 34195 39083
rect 35541 39049 35575 39083
rect 35909 39049 35943 39083
rect 36001 39049 36035 39083
rect 36369 39049 36403 39083
rect 37933 39049 37967 39083
rect 38485 39049 38519 39083
rect 39313 39049 39347 39083
rect 39773 39049 39807 39083
rect 23305 38981 23339 39015
rect 24961 38981 24995 39015
rect 27813 38981 27847 39015
rect 31585 38981 31619 39015
rect 32781 38981 32815 39015
rect 36737 38981 36771 39015
rect 1777 38913 1811 38947
rect 24869 38913 24903 38947
rect 26249 38913 26283 38947
rect 26341 38913 26375 38947
rect 27721 38913 27755 38947
rect 34069 38913 34103 38947
rect 36829 38913 36863 38947
rect 37841 38913 37875 38947
rect 38853 38913 38887 38947
rect 39681 38913 39715 38947
rect 23397 38845 23431 38879
rect 25053 38845 25087 38879
rect 26433 38845 26467 38879
rect 27905 38845 27939 38879
rect 29009 38845 29043 38879
rect 29101 38845 29135 38879
rect 31033 38845 31067 38879
rect 32873 38845 32907 38879
rect 32965 38845 32999 38879
rect 34253 38845 34287 38879
rect 36093 38845 36127 38879
rect 36921 38845 36955 38879
rect 38025 38845 38059 38879
rect 38945 38845 38979 38879
rect 39037 38845 39071 38879
rect 39865 38845 39899 38879
rect 40325 38845 40359 38879
rect 40601 38845 40635 38879
rect 33701 38777 33735 38811
rect 1593 38709 1627 38743
rect 22845 38709 22879 38743
rect 28549 38709 28583 38743
rect 32413 38709 32447 38743
rect 34989 38709 35023 38743
rect 37473 38709 37507 38743
rect 42073 38709 42107 38743
rect 23305 38505 23339 38539
rect 27077 38505 27111 38539
rect 36645 38505 36679 38539
rect 39221 38505 39255 38539
rect 40049 38505 40083 38539
rect 49157 38505 49191 38539
rect 22845 38437 22879 38471
rect 28457 38437 28491 38471
rect 33701 38437 33735 38471
rect 43269 38437 43303 38471
rect 21097 38369 21131 38403
rect 23857 38369 23891 38403
rect 27537 38369 27571 38403
rect 27629 38369 27663 38403
rect 28917 38369 28951 38403
rect 29009 38369 29043 38403
rect 32597 38369 32631 38403
rect 33425 38369 33459 38403
rect 34161 38369 34195 38403
rect 34253 38369 34287 38403
rect 34897 38369 34931 38403
rect 40693 38369 40727 38403
rect 29745 38301 29779 38335
rect 31861 38301 31895 38335
rect 33333 38301 33367 38335
rect 40417 38301 40451 38335
rect 41521 38301 41555 38335
rect 49341 38301 49375 38335
rect 21373 38233 21407 38267
rect 23673 38233 23707 38267
rect 26617 38233 26651 38267
rect 27445 38233 27479 38267
rect 28825 38233 28859 38267
rect 30021 38233 30055 38267
rect 31769 38233 31803 38267
rect 35173 38233 35207 38267
rect 37105 38233 37139 38267
rect 37933 38233 37967 38267
rect 41797 38233 41831 38267
rect 23765 38165 23799 38199
rect 32873 38165 32907 38199
rect 33241 38165 33275 38199
rect 34069 38165 34103 38199
rect 40509 38165 40543 38199
rect 41245 38165 41279 38199
rect 33517 37961 33551 37995
rect 33977 37961 34011 37995
rect 49157 37961 49191 37995
rect 29193 37893 29227 37927
rect 30665 37893 30699 37927
rect 36001 37893 36035 37927
rect 42993 37893 43027 37927
rect 31493 37825 31527 37859
rect 33057 37825 33091 37859
rect 33885 37825 33919 37859
rect 36737 37825 36771 37859
rect 41153 37825 41187 37859
rect 49341 37825 49375 37859
rect 23121 37757 23155 37791
rect 23397 37757 23431 37791
rect 27169 37757 27203 37791
rect 27445 37757 27479 37791
rect 34069 37757 34103 37791
rect 38577 37757 38611 37791
rect 38853 37757 38887 37791
rect 41245 37757 41279 37791
rect 41337 37757 41371 37791
rect 43085 37757 43119 37791
rect 43177 37757 43211 37791
rect 42625 37689 42659 37723
rect 22661 37621 22695 37655
rect 24869 37621 24903 37655
rect 30205 37621 30239 37655
rect 40325 37621 40359 37655
rect 40785 37621 40819 37655
rect 21557 37417 21591 37451
rect 28549 37417 28583 37451
rect 42428 37417 42462 37451
rect 38577 37349 38611 37383
rect 40049 37349 40083 37383
rect 22753 37281 22787 37315
rect 23949 37281 23983 37315
rect 26065 37281 26099 37315
rect 27077 37281 27111 37315
rect 30297 37281 30331 37315
rect 31493 37281 31527 37315
rect 32689 37281 32723 37315
rect 37473 37281 37507 37315
rect 37565 37281 37599 37315
rect 39221 37281 39255 37315
rect 40601 37281 40635 37315
rect 42165 37281 42199 37315
rect 48053 37281 48087 37315
rect 48513 37281 48547 37315
rect 22477 37213 22511 37247
rect 22569 37213 22603 37247
rect 23673 37213 23707 37247
rect 24777 37213 24811 37247
rect 25973 37213 26007 37247
rect 26801 37213 26835 37247
rect 29193 37213 29227 37247
rect 30113 37213 30147 37247
rect 31309 37213 31343 37247
rect 32597 37213 32631 37247
rect 37381 37213 37415 37247
rect 38945 37213 38979 37247
rect 40509 37213 40543 37247
rect 41429 37213 41463 37247
rect 48789 37213 48823 37247
rect 25881 37145 25915 37179
rect 40417 37145 40451 37179
rect 22109 37077 22143 37111
rect 23305 37077 23339 37111
rect 23765 37077 23799 37111
rect 25513 37077 25547 37111
rect 29745 37077 29779 37111
rect 30205 37077 30239 37111
rect 30941 37077 30975 37111
rect 31401 37077 31435 37111
rect 32137 37077 32171 37111
rect 32505 37077 32539 37111
rect 37013 37077 37047 37111
rect 39037 37077 39071 37111
rect 43913 37077 43947 37111
rect 19441 36873 19475 36907
rect 26249 36873 26283 36907
rect 32321 36873 32355 36907
rect 32781 36873 32815 36907
rect 37841 36873 37875 36907
rect 26341 36805 26375 36839
rect 32689 36805 32723 36839
rect 40049 36805 40083 36839
rect 43085 36805 43119 36839
rect 1777 36737 1811 36771
rect 19809 36737 19843 36771
rect 19901 36737 19935 36771
rect 23397 36737 23431 36771
rect 27537 36737 27571 36771
rect 30297 36737 30331 36771
rect 39221 36737 39255 36771
rect 42993 36737 43027 36771
rect 49341 36737 49375 36771
rect 20085 36669 20119 36703
rect 23673 36669 23707 36703
rect 25421 36669 25455 36703
rect 26433 36669 26467 36703
rect 27629 36669 27663 36703
rect 27813 36669 27847 36703
rect 30389 36669 30423 36703
rect 30573 36669 30607 36703
rect 31769 36669 31803 36703
rect 32873 36669 32907 36703
rect 34437 36669 34471 36703
rect 34713 36669 34747 36703
rect 37933 36669 37967 36703
rect 38117 36669 38151 36703
rect 39773 36669 39807 36703
rect 43269 36669 43303 36703
rect 29929 36601 29963 36635
rect 37473 36601 37507 36635
rect 1593 36533 1627 36567
rect 22937 36533 22971 36567
rect 25881 36533 25915 36567
rect 27169 36533 27203 36567
rect 36185 36533 36219 36567
rect 41521 36533 41555 36567
rect 42625 36533 42659 36567
rect 49157 36533 49191 36567
rect 22293 36329 22327 36363
rect 23305 36329 23339 36363
rect 27629 36329 27663 36363
rect 32045 36329 32079 36363
rect 37473 36329 37507 36363
rect 40141 36329 40175 36363
rect 35081 36261 35115 36295
rect 41889 36261 41923 36295
rect 20545 36193 20579 36227
rect 23949 36193 23983 36227
rect 28365 36193 28399 36227
rect 32597 36193 32631 36227
rect 35541 36193 35575 36227
rect 35725 36193 35759 36227
rect 36737 36193 36771 36227
rect 36829 36193 36863 36227
rect 37933 36193 37967 36227
rect 38025 36193 38059 36227
rect 40785 36193 40819 36227
rect 42349 36193 42383 36227
rect 42533 36193 42567 36227
rect 23673 36125 23707 36159
rect 27353 36125 27387 36159
rect 28181 36125 28215 36159
rect 28273 36125 28307 36159
rect 32413 36125 32447 36159
rect 32505 36125 32539 36159
rect 36645 36125 36679 36159
rect 40509 36125 40543 36159
rect 20821 36057 20855 36091
rect 35449 36057 35483 36091
rect 37841 36057 37875 36091
rect 22845 35989 22879 36023
rect 23765 35989 23799 36023
rect 27813 35989 27847 36023
rect 36277 35989 36311 36023
rect 40601 35989 40635 36023
rect 42257 35989 42291 36023
rect 21281 35785 21315 35819
rect 26433 35785 26467 35819
rect 35633 35785 35667 35819
rect 36001 35785 36035 35819
rect 39865 35785 39899 35819
rect 32781 35717 32815 35751
rect 33517 35717 33551 35751
rect 36093 35717 36127 35751
rect 42901 35717 42935 35751
rect 24685 35649 24719 35683
rect 29101 35649 29135 35683
rect 32689 35649 32723 35683
rect 33885 35649 33919 35683
rect 34805 35649 34839 35683
rect 38117 35649 38151 35683
rect 40693 35649 40727 35683
rect 42625 35649 42659 35683
rect 49341 35649 49375 35683
rect 19533 35581 19567 35615
rect 19809 35581 19843 35615
rect 24961 35581 24995 35615
rect 29377 35581 29411 35615
rect 32873 35581 32907 35615
rect 34897 35581 34931 35615
rect 35081 35581 35115 35615
rect 36185 35581 36219 35615
rect 38393 35581 38427 35615
rect 40785 35581 40819 35615
rect 40877 35581 40911 35615
rect 40325 35513 40359 35547
rect 49157 35513 49191 35547
rect 27353 35445 27387 35479
rect 30849 35445 30883 35479
rect 31769 35445 31803 35479
rect 32321 35445 32355 35479
rect 34437 35445 34471 35479
rect 44373 35445 44407 35479
rect 24593 35241 24627 35275
rect 26065 35241 26099 35275
rect 29009 35241 29043 35275
rect 33977 35241 34011 35275
rect 37381 35241 37415 35275
rect 29745 35173 29779 35207
rect 22017 35105 22051 35139
rect 25145 35105 25179 35139
rect 26709 35105 26743 35139
rect 27261 35105 27295 35139
rect 27537 35105 27571 35139
rect 30297 35105 30331 35139
rect 31493 35105 31527 35139
rect 31677 35105 31711 35139
rect 32229 35105 32263 35139
rect 32505 35105 32539 35139
rect 36645 35105 36679 35139
rect 37933 35105 37967 35139
rect 39129 35105 39163 35139
rect 42717 35105 42751 35139
rect 44465 35105 44499 35139
rect 21741 35037 21775 35071
rect 25053 35037 25087 35071
rect 26433 35037 26467 35071
rect 30113 35037 30147 35071
rect 31401 35037 31435 35071
rect 36461 35037 36495 35071
rect 37841 35037 37875 35071
rect 41981 35037 42015 35071
rect 49341 35037 49375 35071
rect 26525 34969 26559 35003
rect 37749 34969 37783 35003
rect 42993 34969 43027 35003
rect 23489 34901 23523 34935
rect 24961 34901 24995 34935
rect 30205 34901 30239 34935
rect 31033 34901 31067 34935
rect 36001 34901 36035 34935
rect 36369 34901 36403 34935
rect 38577 34901 38611 34935
rect 38945 34901 38979 34935
rect 39037 34901 39071 34935
rect 49157 34901 49191 34935
rect 1593 34697 1627 34731
rect 25329 34697 25363 34731
rect 31033 34697 31067 34731
rect 31401 34697 31435 34731
rect 32689 34697 32723 34731
rect 32781 34697 32815 34731
rect 33517 34697 33551 34731
rect 35817 34697 35851 34731
rect 38945 34697 38979 34731
rect 39405 34697 39439 34731
rect 40509 34697 40543 34731
rect 40601 34697 40635 34731
rect 41337 34697 41371 34731
rect 41705 34697 41739 34731
rect 43453 34697 43487 34731
rect 49157 34697 49191 34731
rect 25789 34629 25823 34663
rect 43361 34629 43395 34663
rect 1777 34561 1811 34595
rect 23029 34561 23063 34595
rect 25697 34561 25731 34595
rect 28273 34561 28307 34595
rect 31493 34561 31527 34595
rect 39313 34561 39347 34595
rect 49341 34561 49375 34595
rect 24777 34493 24811 34527
rect 25973 34493 26007 34527
rect 31585 34493 31619 34527
rect 32965 34493 32999 34527
rect 34069 34493 34103 34527
rect 39589 34493 39623 34527
rect 40785 34493 40819 34527
rect 41797 34493 41831 34527
rect 41981 34493 42015 34527
rect 43545 34493 43579 34527
rect 32321 34425 32355 34459
rect 40141 34425 40175 34459
rect 42993 34425 43027 34459
rect 23286 34357 23320 34391
rect 28530 34357 28564 34391
rect 30021 34357 30055 34391
rect 34332 34357 34366 34391
rect 23305 34153 23339 34187
rect 26512 34153 26546 34187
rect 36277 34153 36311 34187
rect 24593 34085 24627 34119
rect 30757 34085 30791 34119
rect 23949 34017 23983 34051
rect 25237 34017 25271 34051
rect 27997 34017 28031 34051
rect 31401 34017 31435 34051
rect 36737 34017 36771 34051
rect 36921 34017 36955 34051
rect 38761 34017 38795 34051
rect 42165 34017 42199 34051
rect 42257 34017 42291 34051
rect 26249 33949 26283 33983
rect 29929 33949 29963 33983
rect 31125 33949 31159 33983
rect 32137 33949 32171 33983
rect 38577 33949 38611 33983
rect 38669 33949 38703 33983
rect 42073 33949 42107 33983
rect 49341 33949 49375 33983
rect 23765 33881 23799 33915
rect 23673 33813 23707 33847
rect 24961 33813 24995 33847
rect 25053 33813 25087 33847
rect 31217 33813 31251 33847
rect 35725 33813 35759 33847
rect 36645 33813 36679 33847
rect 37657 33813 37691 33847
rect 38209 33813 38243 33847
rect 39405 33813 39439 33847
rect 41705 33813 41739 33847
rect 49157 33813 49191 33847
rect 25053 33609 25087 33643
rect 28733 33609 28767 33643
rect 29101 33609 29135 33643
rect 38853 33609 38887 33643
rect 39313 33609 39347 33643
rect 23121 33541 23155 33575
rect 34253 33541 34287 33575
rect 25421 33473 25455 33507
rect 25513 33473 25547 33507
rect 30297 33473 30331 33507
rect 33977 33473 34011 33507
rect 37841 33473 37875 33507
rect 38669 33473 38703 33507
rect 39221 33473 39255 33507
rect 22845 33405 22879 33439
rect 25605 33405 25639 33439
rect 29193 33405 29227 33439
rect 29377 33405 29411 33439
rect 30389 33405 30423 33439
rect 30481 33405 30515 33439
rect 35725 33405 35759 33439
rect 37933 33405 37967 33439
rect 38117 33405 38151 33439
rect 39405 33405 39439 33439
rect 40325 33405 40359 33439
rect 40601 33405 40635 33439
rect 37473 33337 37507 33371
rect 24593 33269 24627 33303
rect 29929 33269 29963 33303
rect 36185 33269 36219 33303
rect 42073 33269 42107 33303
rect 22845 33065 22879 33099
rect 28457 33065 28491 33099
rect 30941 33065 30975 33099
rect 36534 33065 36568 33099
rect 38393 33065 38427 33099
rect 34897 32997 34931 33031
rect 38025 32997 38059 33031
rect 21373 32929 21407 32963
rect 27077 32929 27111 32963
rect 27261 32929 27295 32963
rect 28917 32929 28951 32963
rect 29101 32929 29135 32963
rect 30389 32929 30423 32963
rect 31493 32929 31527 32963
rect 35541 32929 35575 32963
rect 38945 32929 38979 32963
rect 40877 32929 40911 32963
rect 41061 32929 41095 32963
rect 42073 32929 42107 32963
rect 42257 32929 42291 32963
rect 21097 32861 21131 32895
rect 26065 32861 26099 32895
rect 26985 32861 27019 32895
rect 28825 32861 28859 32895
rect 31401 32861 31435 32895
rect 34529 32861 34563 32895
rect 35265 32861 35299 32895
rect 36277 32861 36311 32895
rect 38761 32861 38795 32895
rect 38853 32861 38887 32895
rect 40785 32861 40819 32895
rect 41981 32861 42015 32895
rect 43821 32861 43855 32895
rect 49341 32861 49375 32895
rect 30113 32793 30147 32827
rect 26617 32725 26651 32759
rect 29745 32725 29779 32759
rect 30205 32725 30239 32759
rect 31309 32725 31343 32759
rect 35357 32725 35391 32759
rect 36093 32725 36127 32759
rect 40417 32725 40451 32759
rect 41613 32725 41647 32759
rect 43637 32725 43671 32759
rect 49157 32725 49191 32759
rect 17233 32521 17267 32555
rect 17693 32521 17727 32555
rect 25605 32521 25639 32555
rect 27261 32521 27295 32555
rect 34253 32521 34287 32555
rect 35081 32521 35115 32555
rect 1777 32385 1811 32419
rect 17601 32385 17635 32419
rect 18613 32385 18647 32419
rect 23857 32385 23891 32419
rect 27629 32385 27663 32419
rect 28825 32385 28859 32419
rect 35173 32385 35207 32419
rect 39313 32385 39347 32419
rect 45017 32385 45051 32419
rect 48789 32385 48823 32419
rect 17877 32317 17911 32351
rect 24133 32317 24167 32351
rect 27721 32317 27755 32351
rect 27905 32317 27939 32351
rect 32505 32317 32539 32351
rect 32781 32317 32815 32351
rect 35265 32317 35299 32351
rect 39589 32317 39623 32351
rect 48513 32317 48547 32351
rect 1593 32181 1627 32215
rect 28457 32181 28491 32215
rect 34713 32181 34747 32215
rect 41061 32181 41095 32215
rect 42809 32181 42843 32215
rect 44833 32181 44867 32215
rect 24041 31977 24075 32011
rect 27537 31977 27571 32011
rect 28457 31977 28491 32011
rect 32321 31909 32355 31943
rect 37933 31909 37967 31943
rect 43637 31909 43671 31943
rect 22293 31841 22327 31875
rect 22569 31841 22603 31875
rect 25789 31841 25823 31875
rect 26065 31841 26099 31875
rect 28917 31841 28951 31875
rect 29009 31841 29043 31875
rect 32781 31841 32815 31875
rect 32965 31841 32999 31875
rect 35909 31841 35943 31875
rect 36093 31841 36127 31875
rect 38485 31841 38519 31875
rect 41889 31841 41923 31875
rect 42165 31841 42199 31875
rect 48789 31841 48823 31875
rect 24777 31773 24811 31807
rect 39497 31773 39531 31807
rect 48053 31773 48087 31807
rect 48513 31773 48547 31807
rect 32689 31705 32723 31739
rect 38393 31705 38427 31739
rect 28825 31637 28859 31671
rect 35449 31637 35483 31671
rect 35817 31637 35851 31671
rect 38301 31637 38335 31671
rect 39313 31637 39347 31671
rect 23857 31433 23891 31467
rect 26617 31433 26651 31467
rect 42993 31433 43027 31467
rect 47961 31433 47995 31467
rect 38669 31365 38703 31399
rect 43085 31365 43119 31399
rect 22385 31297 22419 31331
rect 23949 31297 23983 31331
rect 24869 31297 24903 31331
rect 33333 31297 33367 31331
rect 33425 31297 33459 31331
rect 34529 31297 34563 31331
rect 37749 31297 37783 31331
rect 38577 31297 38611 31331
rect 40877 31297 40911 31331
rect 45661 31297 45695 31331
rect 47869 31297 47903 31331
rect 48789 31297 48823 31331
rect 22477 31229 22511 31263
rect 22661 31229 22695 31263
rect 24133 31229 24167 31263
rect 25145 31229 25179 31263
rect 33609 31229 33643 31263
rect 34805 31229 34839 31263
rect 36277 31229 36311 31263
rect 38853 31229 38887 31263
rect 43177 31229 43211 31263
rect 48513 31229 48547 31263
rect 23489 31161 23523 31195
rect 40693 31161 40727 31195
rect 21465 31093 21499 31127
rect 22017 31093 22051 31127
rect 32965 31093 32999 31127
rect 37565 31093 37599 31127
rect 38209 31093 38243 31127
rect 42625 31093 42659 31127
rect 45477 31093 45511 31127
rect 23305 30889 23339 30923
rect 26617 30889 26651 30923
rect 48789 30889 48823 30923
rect 21465 30821 21499 30855
rect 22845 30821 22879 30855
rect 30941 30821 30975 30855
rect 36369 30821 36403 30855
rect 22109 30753 22143 30787
rect 23949 30753 23983 30787
rect 24869 30753 24903 30787
rect 27077 30753 27111 30787
rect 30297 30753 30331 30787
rect 35449 30753 35483 30787
rect 35633 30753 35667 30787
rect 36921 30753 36955 30787
rect 37933 30753 37967 30787
rect 39129 30753 39163 30787
rect 39221 30753 39255 30787
rect 40509 30753 40543 30787
rect 40601 30753 40635 30787
rect 21833 30685 21867 30719
rect 30205 30685 30239 30719
rect 31309 30685 31343 30719
rect 35357 30685 35391 30719
rect 36185 30685 36219 30719
rect 36829 30685 36863 30719
rect 39037 30685 39071 30719
rect 40417 30685 40451 30719
rect 41521 30685 41555 30719
rect 42165 30685 42199 30719
rect 43269 30685 43303 30719
rect 23765 30617 23799 30651
rect 25145 30617 25179 30651
rect 27353 30617 27387 30651
rect 30113 30617 30147 30651
rect 31585 30617 31619 30651
rect 37841 30617 37875 30651
rect 48697 30617 48731 30651
rect 20913 30549 20947 30583
rect 21925 30549 21959 30583
rect 23673 30549 23707 30583
rect 28825 30549 28859 30583
rect 29745 30549 29779 30583
rect 33057 30549 33091 30583
rect 34989 30549 35023 30583
rect 36737 30549 36771 30583
rect 37381 30549 37415 30583
rect 37749 30549 37783 30583
rect 38669 30549 38703 30583
rect 40049 30549 40083 30583
rect 41337 30549 41371 30583
rect 41981 30549 42015 30583
rect 43085 30549 43119 30583
rect 28733 30345 28767 30379
rect 41337 30345 41371 30379
rect 24501 30277 24535 30311
rect 26065 30277 26099 30311
rect 35909 30277 35943 30311
rect 37841 30277 37875 30311
rect 37933 30277 37967 30311
rect 39037 30277 39071 30311
rect 7389 30209 7423 30243
rect 23673 30209 23707 30243
rect 25973 30209 26007 30243
rect 30849 30209 30883 30243
rect 34069 30209 34103 30243
rect 34161 30209 34195 30243
rect 36001 30209 36035 30243
rect 49341 30209 49375 30243
rect 7573 30141 7607 30175
rect 9137 30141 9171 30175
rect 23581 30141 23615 30175
rect 25145 30141 25179 30175
rect 26157 30141 26191 30175
rect 28825 30141 28859 30175
rect 28917 30141 28951 30175
rect 29929 30141 29963 30175
rect 30941 30141 30975 30175
rect 31125 30141 31159 30175
rect 34253 30141 34287 30175
rect 36093 30141 36127 30175
rect 38025 30141 38059 30175
rect 38761 30141 38795 30175
rect 41429 30141 41463 30175
rect 41521 30141 41555 30175
rect 25605 30073 25639 30107
rect 28365 30073 28399 30107
rect 35541 30073 35575 30107
rect 40969 30073 41003 30107
rect 27813 30005 27847 30039
rect 30481 30005 30515 30039
rect 33701 30005 33735 30039
rect 37473 30005 37507 30039
rect 40509 30005 40543 30039
rect 49157 30005 49191 30039
rect 38761 29801 38795 29835
rect 42717 29801 42751 29835
rect 25329 29733 25363 29767
rect 2053 29665 2087 29699
rect 21925 29665 21959 29699
rect 25973 29665 26007 29699
rect 30297 29665 30331 29699
rect 32505 29665 32539 29699
rect 36461 29665 36495 29699
rect 36737 29665 36771 29699
rect 39405 29665 39439 29699
rect 40969 29665 41003 29699
rect 48789 29665 48823 29699
rect 1777 29597 1811 29631
rect 25697 29597 25731 29631
rect 26709 29597 26743 29631
rect 30113 29597 30147 29631
rect 32321 29597 32355 29631
rect 39129 29597 39163 29631
rect 48513 29597 48547 29631
rect 21189 29529 21223 29563
rect 41245 29529 41279 29563
rect 25789 29461 25823 29495
rect 29745 29461 29779 29495
rect 30205 29461 30239 29495
rect 31953 29461 31987 29495
rect 32413 29461 32447 29495
rect 38209 29461 38243 29495
rect 39221 29461 39255 29495
rect 22017 29257 22051 29291
rect 35725 29257 35759 29291
rect 41245 29257 41279 29291
rect 27997 29189 28031 29223
rect 30297 29189 30331 29223
rect 22385 29121 22419 29155
rect 22477 29121 22511 29155
rect 23305 29121 23339 29155
rect 27721 29121 27755 29155
rect 41153 29121 41187 29155
rect 49341 29121 49375 29155
rect 22661 29053 22695 29087
rect 30389 29053 30423 29087
rect 30481 29053 30515 29087
rect 33977 29053 34011 29087
rect 41429 29053 41463 29087
rect 21189 28985 21223 29019
rect 29929 28985 29963 29019
rect 40785 28985 40819 29019
rect 49157 28985 49191 29019
rect 29469 28917 29503 28951
rect 34240 28917 34274 28951
rect 36369 28917 36403 28951
rect 22201 28713 22235 28747
rect 49157 28645 49191 28679
rect 22661 28577 22695 28611
rect 22845 28577 22879 28611
rect 31309 28577 31343 28611
rect 34069 28577 34103 28611
rect 34161 28577 34195 28611
rect 35541 28577 35575 28611
rect 36645 28577 36679 28611
rect 37933 28577 37967 28611
rect 40693 28577 40727 28611
rect 26341 28509 26375 28543
rect 29929 28509 29963 28543
rect 31125 28509 31159 28543
rect 33977 28509 34011 28543
rect 36461 28509 36495 28543
rect 37657 28509 37691 28543
rect 38669 28509 38703 28543
rect 40417 28509 40451 28543
rect 49341 28509 49375 28543
rect 25513 28441 25547 28475
rect 27077 28441 27111 28475
rect 37749 28441 37783 28475
rect 40509 28441 40543 28475
rect 21649 28373 21683 28407
rect 22569 28373 22603 28407
rect 28365 28373 28399 28407
rect 30757 28373 30791 28407
rect 31217 28373 31251 28407
rect 33609 28373 33643 28407
rect 34897 28373 34931 28407
rect 35265 28373 35299 28407
rect 35357 28373 35391 28407
rect 36093 28373 36127 28407
rect 36553 28373 36587 28407
rect 37289 28373 37323 28407
rect 40049 28373 40083 28407
rect 4813 28169 4847 28203
rect 26433 28169 26467 28203
rect 36369 28169 36403 28203
rect 37473 28169 37507 28203
rect 37933 28169 37967 28203
rect 39037 28169 39071 28203
rect 20545 28101 20579 28135
rect 28273 28101 28307 28135
rect 32597 28101 32631 28135
rect 36461 28101 36495 28135
rect 48053 28101 48087 28135
rect 4997 28033 5031 28067
rect 7573 28033 7607 28067
rect 22477 28033 22511 28067
rect 24685 28033 24719 28067
rect 31217 28033 31251 28067
rect 37841 28033 37875 28067
rect 7757 27965 7791 27999
rect 9413 27965 9447 27999
rect 21373 27965 21407 27999
rect 22753 27965 22787 27999
rect 24961 27965 24995 27999
rect 27997 27965 28031 27999
rect 31309 27965 31343 27999
rect 31493 27965 31527 27999
rect 32321 27965 32355 27999
rect 36645 27965 36679 27999
rect 38025 27965 38059 27999
rect 39129 27965 39163 27999
rect 39313 27965 39347 27999
rect 30849 27897 30883 27931
rect 38669 27897 38703 27931
rect 24225 27829 24259 27863
rect 29745 27829 29779 27863
rect 34069 27829 34103 27863
rect 36001 27829 36035 27863
rect 48145 27829 48179 27863
rect 40312 27625 40346 27659
rect 7803 27557 7837 27591
rect 27629 27557 27663 27591
rect 41797 27557 41831 27591
rect 2053 27489 2087 27523
rect 24961 27489 24995 27523
rect 28273 27489 28307 27523
rect 30757 27489 30791 27523
rect 32321 27489 32355 27523
rect 35357 27489 35391 27523
rect 35541 27489 35575 27523
rect 40049 27489 40083 27523
rect 1777 27421 1811 27455
rect 7732 27421 7766 27455
rect 23397 27421 23431 27455
rect 27997 27421 28031 27455
rect 32965 27421 32999 27455
rect 35265 27421 35299 27455
rect 37013 27421 37047 27455
rect 44189 27421 44223 27455
rect 47225 27421 47259 27455
rect 48513 27421 48547 27455
rect 48789 27421 48823 27455
rect 25237 27353 25271 27387
rect 30573 27353 30607 27387
rect 32137 27353 32171 27387
rect 33793 27353 33827 27387
rect 37289 27353 37323 27387
rect 47409 27353 47443 27387
rect 26709 27285 26743 27319
rect 28089 27285 28123 27319
rect 30205 27285 30239 27319
rect 30665 27285 30699 27319
rect 31769 27285 31803 27319
rect 32229 27285 32263 27319
rect 34897 27285 34931 27319
rect 38761 27285 38795 27319
rect 44005 27285 44039 27319
rect 23121 27081 23155 27115
rect 31125 27081 31159 27115
rect 42073 27081 42107 27115
rect 23213 27013 23247 27047
rect 24133 27013 24167 27047
rect 34529 27013 34563 27047
rect 38577 27013 38611 27047
rect 47869 27013 47903 27047
rect 7849 26945 7883 26979
rect 33425 26945 33459 26979
rect 36921 26945 36955 26979
rect 37749 26945 37783 26979
rect 40332 26945 40366 26979
rect 47041 26945 47075 26979
rect 48789 26945 48823 26979
rect 8033 26877 8067 26911
rect 9597 26877 9631 26911
rect 23397 26877 23431 26911
rect 28549 26877 28583 26911
rect 28825 26877 28859 26911
rect 31217 26877 31251 26911
rect 31401 26877 31435 26911
rect 33517 26877 33551 26911
rect 33701 26877 33735 26911
rect 34260 26877 34294 26911
rect 40601 26877 40635 26911
rect 48513 26877 48547 26911
rect 22753 26809 22787 26843
rect 24225 26741 24259 26775
rect 27353 26741 27387 26775
rect 30297 26741 30331 26775
rect 30757 26741 30791 26775
rect 33057 26741 33091 26775
rect 36001 26741 36035 26775
rect 36737 26741 36771 26775
rect 46857 26741 46891 26775
rect 47961 26741 47995 26775
rect 7895 26537 7929 26571
rect 9689 26537 9723 26571
rect 30757 26537 30791 26571
rect 41797 26537 41831 26571
rect 23857 26469 23891 26503
rect 26617 26469 26651 26503
rect 38761 26469 38795 26503
rect 9137 26401 9171 26435
rect 22109 26401 22143 26435
rect 22385 26401 22419 26435
rect 25053 26401 25087 26435
rect 25145 26401 25179 26435
rect 27169 26401 27203 26435
rect 28365 26401 28399 26435
rect 31217 26401 31251 26435
rect 31309 26401 31343 26435
rect 32229 26401 32263 26435
rect 33977 26401 34011 26435
rect 39221 26401 39255 26435
rect 39405 26401 39439 26435
rect 40049 26401 40083 26435
rect 48789 26401 48823 26435
rect 7792 26333 7826 26367
rect 9321 26333 9355 26367
rect 26985 26333 27019 26367
rect 28181 26333 28215 26367
rect 28273 26333 28307 26367
rect 31125 26333 31159 26367
rect 34897 26333 34931 26367
rect 36921 26333 36955 26367
rect 39129 26333 39163 26367
rect 47409 26333 47443 26367
rect 48053 26333 48087 26367
rect 48513 26333 48547 26367
rect 24961 26265 24995 26299
rect 32505 26265 32539 26299
rect 35633 26265 35667 26299
rect 37657 26265 37691 26299
rect 40325 26265 40359 26299
rect 24593 26197 24627 26231
rect 27077 26197 27111 26231
rect 27813 26197 27847 26231
rect 47225 26197 47259 26231
rect 31493 25993 31527 26027
rect 32321 25993 32355 26027
rect 32689 25993 32723 26027
rect 37841 25993 37875 26027
rect 37933 25993 37967 26027
rect 39037 25993 39071 26027
rect 39129 25993 39163 26027
rect 42073 25993 42107 26027
rect 32781 25925 32815 25959
rect 35357 25925 35391 25959
rect 40601 25925 40635 25959
rect 46121 25925 46155 25959
rect 7573 25857 7607 25891
rect 24133 25857 24167 25891
rect 25145 25857 25179 25891
rect 31401 25857 31435 25891
rect 35265 25857 35299 25891
rect 40325 25857 40359 25891
rect 46857 25857 46891 25891
rect 49341 25857 49375 25891
rect 7757 25789 7791 25823
rect 9413 25789 9447 25823
rect 24225 25789 24259 25823
rect 24409 25789 24443 25823
rect 28457 25789 28491 25823
rect 28733 25789 28767 25823
rect 31677 25789 31711 25823
rect 32965 25789 32999 25823
rect 35541 25789 35575 25823
rect 38117 25789 38151 25823
rect 39221 25789 39255 25823
rect 46305 25721 46339 25755
rect 47041 25721 47075 25755
rect 23765 25653 23799 25687
rect 26065 25653 26099 25687
rect 30205 25653 30239 25687
rect 31033 25653 31067 25687
rect 34897 25653 34931 25687
rect 36921 25653 36955 25687
rect 37473 25653 37507 25687
rect 38669 25653 38703 25687
rect 49157 25653 49191 25687
rect 4997 25449 5031 25483
rect 10793 25449 10827 25483
rect 11069 25449 11103 25483
rect 27721 25449 27755 25483
rect 39497 25449 39531 25483
rect 14289 25381 14323 25415
rect 2053 25313 2087 25347
rect 22937 25313 22971 25347
rect 25145 25313 25179 25347
rect 28917 25313 28951 25347
rect 31401 25313 31435 25347
rect 32505 25313 32539 25347
rect 32597 25313 32631 25347
rect 33977 25313 34011 25347
rect 34069 25313 34103 25347
rect 35725 25313 35759 25347
rect 37013 25313 37047 25347
rect 37197 25313 37231 25347
rect 40509 25313 40543 25347
rect 40693 25313 40727 25347
rect 1777 25245 1811 25279
rect 5181 25245 5215 25279
rect 10609 25245 10643 25279
rect 14473 25245 14507 25279
rect 24041 25245 24075 25279
rect 24961 25245 24995 25279
rect 25973 25245 26007 25279
rect 28733 25245 28767 25279
rect 28825 25245 28859 25279
rect 29929 25245 29963 25279
rect 31309 25245 31343 25279
rect 32413 25245 32447 25279
rect 37749 25245 37783 25279
rect 45293 25245 45327 25279
rect 46029 25245 46063 25279
rect 22753 25177 22787 25211
rect 26249 25177 26283 25211
rect 31217 25177 31251 25211
rect 33885 25177 33919 25211
rect 35633 25177 35667 25211
rect 36921 25177 36955 25211
rect 38025 25177 38059 25211
rect 44465 25177 44499 25211
rect 44649 25177 44683 25211
rect 45477 25177 45511 25211
rect 46213 25177 46247 25211
rect 22293 25109 22327 25143
rect 22661 25109 22695 25143
rect 24593 25109 24627 25143
rect 25053 25109 25087 25143
rect 28365 25109 28399 25143
rect 30849 25109 30883 25143
rect 32045 25109 32079 25143
rect 33517 25109 33551 25143
rect 35173 25109 35207 25143
rect 35541 25109 35575 25143
rect 36553 25109 36587 25143
rect 40049 25109 40083 25143
rect 40417 25109 40451 25143
rect 32873 24905 32907 24939
rect 37841 24905 37875 24939
rect 25881 24837 25915 24871
rect 29653 24837 29687 24871
rect 8452 24769 8486 24803
rect 22937 24769 22971 24803
rect 27169 24769 27203 24803
rect 29377 24769 29411 24803
rect 32965 24769 32999 24803
rect 36921 24769 36955 24803
rect 37933 24769 37967 24803
rect 40233 24769 40267 24803
rect 47961 24769 47995 24803
rect 8539 24701 8573 24735
rect 19717 24701 19751 24735
rect 19993 24701 20027 24735
rect 25973 24701 26007 24735
rect 26157 24701 26191 24735
rect 31125 24701 31159 24735
rect 33149 24701 33183 24735
rect 33977 24701 34011 24735
rect 34253 24701 34287 24735
rect 36001 24701 36035 24735
rect 38117 24701 38151 24735
rect 49157 24701 49191 24735
rect 25513 24633 25547 24667
rect 36737 24633 36771 24667
rect 21465 24565 21499 24599
rect 27432 24565 27466 24599
rect 28917 24565 28951 24599
rect 32505 24565 32539 24599
rect 37473 24565 37507 24599
rect 10977 24361 11011 24395
rect 20821 24225 20855 24259
rect 25513 24225 25547 24259
rect 25605 24225 25639 24259
rect 26709 24225 26743 24259
rect 26893 24225 26927 24259
rect 28089 24225 28123 24259
rect 28273 24225 28307 24259
rect 30205 24225 30239 24259
rect 30297 24225 30331 24259
rect 34253 24225 34287 24259
rect 34989 24225 35023 24259
rect 35265 24225 35299 24259
rect 37749 24225 37783 24259
rect 40509 24225 40543 24259
rect 40693 24225 40727 24259
rect 10701 24157 10735 24191
rect 30113 24157 30147 24191
rect 33977 24157 34011 24191
rect 37657 24157 37691 24191
rect 40417 24157 40451 24191
rect 47961 24157 47995 24191
rect 21097 24089 21131 24123
rect 27997 24089 28031 24123
rect 37565 24089 37599 24123
rect 49157 24089 49191 24123
rect 11161 24021 11195 24055
rect 22569 24021 22603 24055
rect 25053 24021 25087 24055
rect 25421 24021 25455 24055
rect 26249 24021 26283 24055
rect 26617 24021 26651 24055
rect 27629 24021 27663 24055
rect 29745 24021 29779 24055
rect 33609 24021 33643 24055
rect 34069 24021 34103 24055
rect 36737 24021 36771 24055
rect 37197 24021 37231 24055
rect 40049 24021 40083 24055
rect 9505 23817 9539 23851
rect 16313 23817 16347 23851
rect 19349 23817 19383 23851
rect 19717 23817 19751 23851
rect 20729 23817 20763 23851
rect 21097 23817 21131 23851
rect 26249 23817 26283 23851
rect 27813 23817 27847 23851
rect 28641 23817 28675 23851
rect 34069 23817 34103 23851
rect 40509 23817 40543 23851
rect 12633 23749 12667 23783
rect 34989 23749 35023 23783
rect 39037 23749 39071 23783
rect 8861 23681 8895 23715
rect 12357 23681 12391 23715
rect 22017 23681 22051 23715
rect 25421 23681 25455 23715
rect 32321 23681 32355 23715
rect 34897 23681 34931 23715
rect 38761 23681 38795 23715
rect 47961 23681 47995 23715
rect 9045 23613 9079 23647
rect 14565 23613 14599 23647
rect 14841 23613 14875 23647
rect 19809 23613 19843 23647
rect 19993 23613 20027 23647
rect 21189 23613 21223 23647
rect 21281 23613 21315 23647
rect 22293 23613 22327 23647
rect 24041 23613 24075 23647
rect 26341 23613 26375 23647
rect 26433 23613 26467 23647
rect 28733 23613 28767 23647
rect 28825 23613 28859 23647
rect 35173 23613 35207 23647
rect 49157 23613 49191 23647
rect 14105 23545 14139 23579
rect 24777 23477 24811 23511
rect 25881 23477 25915 23511
rect 28273 23477 28307 23511
rect 32584 23477 32618 23511
rect 34529 23477 34563 23511
rect 5181 23273 5215 23307
rect 28917 23273 28951 23307
rect 31861 23273 31895 23307
rect 36645 23273 36679 23307
rect 34069 23205 34103 23239
rect 37473 23205 37507 23239
rect 2053 23137 2087 23171
rect 9275 23137 9309 23171
rect 17141 23137 17175 23171
rect 19441 23137 19475 23171
rect 23673 23137 23707 23171
rect 25237 23137 25271 23171
rect 27169 23137 27203 23171
rect 30113 23137 30147 23171
rect 34897 23137 34931 23171
rect 38853 23137 38887 23171
rect 1777 23069 1811 23103
rect 4169 23069 4203 23103
rect 9188 23069 9222 23103
rect 23397 23069 23431 23103
rect 24961 23069 24995 23103
rect 32321 23069 32355 23103
rect 37657 23069 37691 23103
rect 38577 23069 38611 23103
rect 40233 23069 40267 23103
rect 47961 23069 47995 23103
rect 5089 23001 5123 23035
rect 17417 23001 17451 23035
rect 19717 23001 19751 23035
rect 23489 23001 23523 23035
rect 27445 23001 27479 23035
rect 30389 23001 30423 23035
rect 32597 23001 32631 23035
rect 35173 23001 35207 23035
rect 38669 23001 38703 23035
rect 49157 23001 49191 23035
rect 4261 22933 4295 22967
rect 18889 22933 18923 22967
rect 21189 22933 21223 22967
rect 23029 22933 23063 22967
rect 24593 22933 24627 22967
rect 25053 22933 25087 22967
rect 38209 22933 38243 22967
rect 17785 22729 17819 22763
rect 19441 22729 19475 22763
rect 19809 22729 19843 22763
rect 30021 22729 30055 22763
rect 30113 22729 30147 22763
rect 31033 22729 31067 22763
rect 34069 22729 34103 22763
rect 21189 22661 21223 22695
rect 23765 22661 23799 22695
rect 31493 22661 31527 22695
rect 34161 22661 34195 22695
rect 44281 22661 44315 22695
rect 21097 22593 21131 22627
rect 23673 22593 23707 22627
rect 24961 22593 24995 22627
rect 25973 22593 26007 22627
rect 27169 22593 27203 22627
rect 31401 22593 31435 22627
rect 32505 22593 32539 22627
rect 37565 22593 37599 22627
rect 17877 22525 17911 22559
rect 17969 22525 18003 22559
rect 19901 22525 19935 22559
rect 19993 22525 20027 22559
rect 21281 22525 21315 22559
rect 23949 22525 23983 22559
rect 25053 22525 25087 22559
rect 25237 22525 25271 22559
rect 28917 22525 28951 22559
rect 30205 22525 30239 22559
rect 31677 22525 31711 22559
rect 34253 22525 34287 22559
rect 37841 22525 37875 22559
rect 39589 22525 39623 22559
rect 20729 22457 20763 22491
rect 24593 22457 24627 22491
rect 29653 22457 29687 22491
rect 44465 22457 44499 22491
rect 17417 22389 17451 22423
rect 23305 22389 23339 22423
rect 27432 22389 27466 22423
rect 33701 22389 33735 22423
rect 12909 22185 12943 22219
rect 15098 22185 15132 22219
rect 23305 22185 23339 22219
rect 35614 22185 35648 22219
rect 5549 22117 5583 22151
rect 25145 22117 25179 22151
rect 21465 22049 21499 22083
rect 22661 22049 22695 22083
rect 23949 22049 23983 22083
rect 26065 22049 26099 22083
rect 26249 22049 26283 22083
rect 29009 22049 29043 22083
rect 37105 22049 37139 22083
rect 12633 21981 12667 22015
rect 13737 21981 13771 22015
rect 14841 21981 14875 22015
rect 23765 21981 23799 22015
rect 25973 21981 26007 22015
rect 29929 21981 29963 22015
rect 35357 21981 35391 22015
rect 37841 21981 37875 22015
rect 47961 21981 47995 22015
rect 49157 21981 49191 22015
rect 5365 21913 5399 21947
rect 21281 21913 21315 21947
rect 21373 21913 21407 21947
rect 22477 21913 22511 21947
rect 23673 21913 23707 21947
rect 28825 21913 28859 21947
rect 13093 21845 13127 21879
rect 13553 21845 13587 21879
rect 16589 21845 16623 21879
rect 20913 21845 20947 21879
rect 22109 21845 22143 21879
rect 22569 21845 22603 21879
rect 25605 21845 25639 21879
rect 28457 21845 28491 21879
rect 28917 21845 28951 21879
rect 37657 21845 37691 21879
rect 10241 21641 10275 21675
rect 14289 21641 14323 21675
rect 25145 21641 25179 21675
rect 25513 21641 25547 21675
rect 29009 21641 29043 21675
rect 31585 21641 31619 21675
rect 29101 21573 29135 21607
rect 38761 21573 38795 21607
rect 9597 21505 9631 21539
rect 14473 21505 14507 21539
rect 19257 21505 19291 21539
rect 28181 21505 28215 21539
rect 32505 21505 32539 21539
rect 35265 21505 35299 21539
rect 36001 21505 36035 21539
rect 38485 21505 38519 21539
rect 47961 21505 47995 21539
rect 9781 21437 9815 21471
rect 19533 21437 19567 21471
rect 22477 21437 22511 21471
rect 22753 21437 22787 21471
rect 25605 21437 25639 21471
rect 25697 21437 25731 21471
rect 29285 21437 29319 21471
rect 29837 21437 29871 21471
rect 30113 21437 30147 21471
rect 32781 21437 32815 21471
rect 40233 21437 40267 21471
rect 49157 21437 49191 21471
rect 21005 21301 21039 21335
rect 24225 21301 24259 21335
rect 27997 21301 28031 21335
rect 28641 21301 28675 21335
rect 34253 21301 34287 21335
rect 35081 21301 35115 21335
rect 35817 21301 35851 21335
rect 9689 21097 9723 21131
rect 19441 21097 19475 21131
rect 36645 21029 36679 21063
rect 9137 20961 9171 20995
rect 20085 20961 20119 20995
rect 30941 20961 30975 20995
rect 38393 20961 38427 20995
rect 4169 20893 4203 20927
rect 9321 20893 9355 20927
rect 19809 20893 19843 20927
rect 30665 20893 30699 20927
rect 31677 20893 31711 20927
rect 32321 20893 32355 20927
rect 36829 20893 36863 20927
rect 38209 20893 38243 20927
rect 43821 20893 43855 20927
rect 47961 20893 47995 20927
rect 44005 20825 44039 20859
rect 49157 20825 49191 20859
rect 4261 20757 4295 20791
rect 19901 20757 19935 20791
rect 30297 20757 30331 20791
rect 30757 20757 30791 20791
rect 32137 20757 32171 20791
rect 37841 20757 37875 20791
rect 38301 20757 38335 20791
rect 21189 20553 21223 20587
rect 24869 20553 24903 20587
rect 26249 20553 26283 20587
rect 30021 20553 30055 20587
rect 30481 20553 30515 20587
rect 32873 20553 32907 20587
rect 23397 20485 23431 20519
rect 30389 20485 30423 20519
rect 32781 20485 32815 20519
rect 1777 20417 1811 20451
rect 21097 20417 21131 20451
rect 23121 20417 23155 20451
rect 26157 20417 26191 20451
rect 36921 20417 36955 20451
rect 47961 20417 47995 20451
rect 2053 20349 2087 20383
rect 21373 20349 21407 20383
rect 26433 20349 26467 20383
rect 30665 20349 30699 20383
rect 33057 20349 33091 20383
rect 49157 20349 49191 20383
rect 20729 20213 20763 20247
rect 25789 20213 25823 20247
rect 32413 20213 32447 20247
rect 36737 20213 36771 20247
rect 14289 20009 14323 20043
rect 18153 20009 18187 20043
rect 22096 20009 22130 20043
rect 25237 20009 25271 20043
rect 26801 20009 26835 20043
rect 35633 20009 35667 20043
rect 18613 19873 18647 19907
rect 18797 19873 18831 19907
rect 19625 19873 19659 19907
rect 21833 19873 21867 19907
rect 25789 19873 25823 19907
rect 27445 19873 27479 19907
rect 14473 19805 14507 19839
rect 18521 19805 18555 19839
rect 27169 19805 27203 19839
rect 32321 19805 32355 19839
rect 33149 19805 33183 19839
rect 33885 19805 33919 19839
rect 34989 19805 35023 19839
rect 35817 19805 35851 19839
rect 44189 19805 44223 19839
rect 19901 19737 19935 19771
rect 25605 19737 25639 19771
rect 34069 19737 34103 19771
rect 44373 19737 44407 19771
rect 21373 19669 21407 19703
rect 23581 19669 23615 19703
rect 25697 19669 25731 19703
rect 27261 19669 27295 19703
rect 32413 19669 32447 19703
rect 33241 19669 33275 19703
rect 35081 19669 35115 19703
rect 19533 19465 19567 19499
rect 19901 19465 19935 19499
rect 20729 19465 20763 19499
rect 21097 19465 21131 19499
rect 39221 19465 39255 19499
rect 21189 19397 21223 19431
rect 22017 19397 22051 19431
rect 22753 19397 22787 19431
rect 23857 19397 23891 19431
rect 28273 19397 28307 19431
rect 29653 19397 29687 19431
rect 19993 19329 20027 19363
rect 23765 19329 23799 19363
rect 24582 19329 24616 19363
rect 26617 19329 26651 19363
rect 33701 19329 33735 19363
rect 37473 19329 37507 19363
rect 47961 19329 47995 19363
rect 49157 19329 49191 19363
rect 20177 19261 20211 19295
rect 21281 19261 21315 19295
rect 24041 19261 24075 19295
rect 24869 19261 24903 19295
rect 29009 19261 29043 19295
rect 30389 19261 30423 19295
rect 33977 19261 34011 19295
rect 35449 19261 35483 19295
rect 37749 19261 37783 19295
rect 23397 19193 23431 19227
rect 18153 18921 18187 18955
rect 20545 18921 20579 18955
rect 23305 18921 23339 18955
rect 24593 18921 24627 18955
rect 27169 18921 27203 18955
rect 18337 18853 18371 18887
rect 31033 18853 31067 18887
rect 21189 18785 21223 18819
rect 23857 18785 23891 18819
rect 25145 18785 25179 18819
rect 26433 18785 26467 18819
rect 26617 18785 26651 18819
rect 27813 18785 27847 18819
rect 28825 18785 28859 18819
rect 28917 18785 28951 18819
rect 31493 18785 31527 18819
rect 31677 18785 31711 18819
rect 36921 18785 36955 18819
rect 4629 18717 4663 18751
rect 17877 18717 17911 18751
rect 21741 18717 21775 18751
rect 23673 18717 23707 18751
rect 27537 18717 27571 18751
rect 36277 18717 36311 18751
rect 44189 18717 44223 18751
rect 47961 18717 47995 18751
rect 20913 18649 20947 18683
rect 22569 18649 22603 18683
rect 23765 18649 23799 18683
rect 25053 18649 25087 18683
rect 28733 18649 28767 18683
rect 31401 18649 31435 18683
rect 36461 18649 36495 18683
rect 37197 18649 37231 18683
rect 44373 18649 44407 18683
rect 49157 18649 49191 18683
rect 4721 18581 4755 18615
rect 21005 18581 21039 18615
rect 24961 18581 24995 18615
rect 25973 18581 26007 18615
rect 26341 18581 26375 18615
rect 27629 18581 27663 18615
rect 28365 18581 28399 18615
rect 38669 18581 38703 18615
rect 19809 18377 19843 18411
rect 20729 18377 20763 18411
rect 21189 18377 21223 18411
rect 27353 18377 27387 18411
rect 27813 18377 27847 18411
rect 29837 18377 29871 18411
rect 34069 18377 34103 18411
rect 37841 18377 37875 18411
rect 37933 18377 37967 18411
rect 19901 18309 19935 18343
rect 23305 18309 23339 18343
rect 25053 18309 25087 18343
rect 30205 18309 30239 18343
rect 30297 18309 30331 18343
rect 32597 18309 32631 18343
rect 1777 18241 1811 18275
rect 21097 18241 21131 18275
rect 27721 18241 27755 18275
rect 47961 18241 47995 18275
rect 2053 18173 2087 18207
rect 20085 18173 20119 18207
rect 21281 18173 21315 18207
rect 23029 18173 23063 18207
rect 27905 18173 27939 18207
rect 30389 18173 30423 18207
rect 32321 18173 32355 18207
rect 34529 18173 34563 18207
rect 34805 18173 34839 18207
rect 38117 18173 38151 18207
rect 49157 18173 49191 18207
rect 19441 18037 19475 18071
rect 36277 18037 36311 18071
rect 37473 18037 37507 18071
rect 19901 17833 19935 17867
rect 27353 17833 27387 17867
rect 32413 17833 32447 17867
rect 37289 17833 37323 17867
rect 20545 17697 20579 17731
rect 21373 17697 21407 17731
rect 23121 17697 23155 17731
rect 27905 17697 27939 17731
rect 30665 17697 30699 17731
rect 33793 17697 33827 17731
rect 33977 17697 34011 17731
rect 35541 17697 35575 17731
rect 37749 17697 37783 17731
rect 38025 17697 38059 17731
rect 44649 17697 44683 17731
rect 21097 17629 21131 17663
rect 23765 17629 23799 17663
rect 27721 17629 27755 17663
rect 27813 17629 27847 17663
rect 42993 17629 43027 17663
rect 43729 17629 43763 17663
rect 43913 17629 43947 17663
rect 47961 17629 47995 17663
rect 30021 17561 30055 17595
rect 30941 17561 30975 17595
rect 35817 17561 35851 17595
rect 44465 17561 44499 17595
rect 49157 17561 49191 17595
rect 20269 17493 20303 17527
rect 20361 17493 20395 17527
rect 30113 17493 30147 17527
rect 33333 17493 33367 17527
rect 33701 17493 33735 17527
rect 39497 17493 39531 17527
rect 43085 17493 43119 17527
rect 21465 17289 21499 17323
rect 22845 17289 22879 17323
rect 23213 17289 23247 17323
rect 24409 17289 24443 17323
rect 27261 17289 27295 17323
rect 28825 17289 28859 17323
rect 33977 17289 34011 17323
rect 34069 17289 34103 17323
rect 19993 17221 20027 17255
rect 43729 17221 43763 17255
rect 23305 17153 23339 17187
rect 24501 17153 24535 17187
rect 27629 17153 27663 17187
rect 32505 17153 32539 17187
rect 35173 17153 35207 17187
rect 36185 17153 36219 17187
rect 19717 17085 19751 17119
rect 23397 17085 23431 17119
rect 24593 17085 24627 17119
rect 27721 17085 27755 17119
rect 27813 17085 27847 17119
rect 28917 17085 28951 17119
rect 29009 17085 29043 17119
rect 30021 17085 30055 17119
rect 30297 17085 30331 17119
rect 31769 17085 31803 17119
rect 34253 17085 34287 17119
rect 35265 17085 35299 17119
rect 35357 17085 35391 17119
rect 24041 17017 24075 17051
rect 33609 17017 33643 17051
rect 43913 17017 43947 17051
rect 28457 16949 28491 16983
rect 32321 16949 32355 16983
rect 34805 16949 34839 16983
rect 38117 16949 38151 16983
rect 23397 16745 23431 16779
rect 26525 16745 26559 16779
rect 19441 16609 19475 16643
rect 21649 16609 21683 16643
rect 21925 16609 21959 16643
rect 24777 16609 24811 16643
rect 25053 16609 25087 16643
rect 27721 16609 27755 16643
rect 34069 16609 34103 16643
rect 34253 16609 34287 16643
rect 34897 16609 34931 16643
rect 35173 16609 35207 16643
rect 38025 16609 38059 16643
rect 27537 16541 27571 16575
rect 33977 16541 34011 16575
rect 37841 16541 37875 16575
rect 47961 16541 47995 16575
rect 5549 16473 5583 16507
rect 19717 16473 19751 16507
rect 27629 16473 27663 16507
rect 37933 16473 37967 16507
rect 49157 16473 49191 16507
rect 5641 16405 5675 16439
rect 21189 16405 21223 16439
rect 27169 16405 27203 16439
rect 33609 16405 33643 16439
rect 36645 16405 36679 16439
rect 37473 16405 37507 16439
rect 25697 16201 25731 16235
rect 27169 16201 27203 16235
rect 27629 16201 27663 16235
rect 33425 16201 33459 16235
rect 23029 16133 23063 16167
rect 24777 16133 24811 16167
rect 27537 16133 27571 16167
rect 1777 16065 1811 16099
rect 33333 16065 33367 16099
rect 34345 16065 34379 16099
rect 36277 16065 36311 16099
rect 38945 16065 38979 16099
rect 47961 16065 47995 16099
rect 2053 15997 2087 16031
rect 22753 15997 22787 16031
rect 25789 15997 25823 16031
rect 25973 15997 26007 16031
rect 27721 15997 27755 16031
rect 28825 15997 28859 16031
rect 29101 15997 29135 16031
rect 33609 15997 33643 16031
rect 49157 15997 49191 16031
rect 32965 15929 32999 15963
rect 25329 15861 25363 15895
rect 30573 15861 30607 15895
rect 34989 15861 35023 15895
rect 36093 15861 36127 15895
rect 37657 15861 37691 15895
rect 38761 15861 38795 15895
rect 26525 15657 26559 15691
rect 31493 15657 31527 15691
rect 33057 15657 33091 15691
rect 27721 15589 27755 15623
rect 26065 15521 26099 15555
rect 27169 15521 27203 15555
rect 28273 15521 28307 15555
rect 29745 15521 29779 15555
rect 30021 15521 30055 15555
rect 33609 15521 33643 15555
rect 35817 15521 35851 15555
rect 36093 15521 36127 15555
rect 28089 15453 28123 15487
rect 28181 15453 28215 15487
rect 32597 15453 32631 15487
rect 33425 15453 33459 15487
rect 47961 15453 47995 15487
rect 24685 15385 24719 15419
rect 25881 15385 25915 15419
rect 26893 15385 26927 15419
rect 26985 15385 27019 15419
rect 29009 15385 29043 15419
rect 33517 15385 33551 15419
rect 49157 15385 49191 15419
rect 24777 15317 24811 15351
rect 29101 15317 29135 15351
rect 32413 15317 32447 15351
rect 37565 15317 37599 15351
rect 21005 15113 21039 15147
rect 24225 15113 24259 15147
rect 26341 15113 26375 15147
rect 29469 15113 29503 15147
rect 32781 15113 32815 15147
rect 37841 15113 37875 15147
rect 30021 15045 30055 15079
rect 31585 15045 31619 15079
rect 37933 15045 37967 15079
rect 20913 14977 20947 15011
rect 22477 14977 22511 15011
rect 26249 14977 26283 15011
rect 32689 14977 32723 15011
rect 41981 14977 42015 15011
rect 47961 14977 47995 15011
rect 21189 14909 21223 14943
rect 22753 14909 22787 14943
rect 26525 14909 26559 14943
rect 27721 14909 27755 14943
rect 27997 14909 28031 14943
rect 30205 14909 30239 14943
rect 32873 14909 32907 14943
rect 38025 14909 38059 14943
rect 49157 14909 49191 14943
rect 25881 14841 25915 14875
rect 31769 14841 31803 14875
rect 20545 14773 20579 14807
rect 30849 14773 30883 14807
rect 32321 14773 32355 14807
rect 37473 14773 37507 14807
rect 41797 14773 41831 14807
rect 32229 14569 32263 14603
rect 27629 14501 27663 14535
rect 29837 14501 29871 14535
rect 32689 14501 32723 14535
rect 37197 14501 37231 14535
rect 25881 14433 25915 14467
rect 30389 14433 30423 14467
rect 33149 14433 33183 14467
rect 33333 14433 33367 14467
rect 37657 14433 37691 14467
rect 37749 14433 37783 14467
rect 30205 14365 30239 14399
rect 33057 14365 33091 14399
rect 34989 14365 35023 14399
rect 37565 14365 37599 14399
rect 38577 14365 38611 14399
rect 40233 14365 40267 14399
rect 26157 14297 26191 14331
rect 35173 14297 35207 14331
rect 30297 14229 30331 14263
rect 40049 14229 40083 14263
rect 36737 14025 36771 14059
rect 38945 14025 38979 14059
rect 29009 13957 29043 13991
rect 37565 13957 37599 13991
rect 37749 13957 37783 13991
rect 1777 13889 1811 13923
rect 30573 13889 30607 13923
rect 33885 13889 33919 13923
rect 36921 13889 36955 13923
rect 38301 13889 38335 13923
rect 39129 13889 39163 13923
rect 41981 13889 42015 13923
rect 47961 13889 47995 13923
rect 2789 13821 2823 13855
rect 29193 13821 29227 13855
rect 35633 13821 35667 13855
rect 38485 13821 38519 13855
rect 49157 13821 49191 13855
rect 30389 13753 30423 13787
rect 41797 13753 41831 13787
rect 34148 13685 34182 13719
rect 28273 13481 28307 13515
rect 36645 13481 36679 13515
rect 28825 13345 28859 13379
rect 34897 13345 34931 13379
rect 35173 13345 35207 13379
rect 25697 13277 25731 13311
rect 28733 13277 28767 13311
rect 34161 13277 34195 13311
rect 37197 13277 37231 13311
rect 38117 13277 38151 13311
rect 40693 13277 40727 13311
rect 47961 13277 47995 13311
rect 28641 13209 28675 13243
rect 49157 13209 49191 13243
rect 25789 13141 25823 13175
rect 34253 13141 34287 13175
rect 37289 13141 37323 13175
rect 37933 13141 37967 13175
rect 40785 13141 40819 13175
rect 28825 12937 28859 12971
rect 29285 12937 29319 12971
rect 30481 12937 30515 12971
rect 35449 12937 35483 12971
rect 27261 12869 27295 12903
rect 27997 12869 28031 12903
rect 29193 12869 29227 12903
rect 33977 12869 34011 12903
rect 43821 12869 43855 12903
rect 30389 12801 30423 12835
rect 33701 12801 33735 12835
rect 36277 12801 36311 12835
rect 47961 12801 47995 12835
rect 29469 12733 29503 12767
rect 30573 12733 30607 12767
rect 36369 12733 36403 12767
rect 36461 12733 36495 12767
rect 49157 12733 49191 12767
rect 28181 12665 28215 12699
rect 30021 12665 30055 12699
rect 44005 12665 44039 12699
rect 27353 12597 27387 12631
rect 35909 12597 35943 12631
rect 36553 12393 36587 12427
rect 28825 12189 28859 12223
rect 39037 12189 39071 12223
rect 41429 12189 41463 12223
rect 44465 12189 44499 12223
rect 47961 12189 47995 12223
rect 29009 12121 29043 12155
rect 39221 12121 39255 12155
rect 49157 12121 49191 12155
rect 41245 12053 41279 12087
rect 44281 12053 44315 12087
rect 46213 11781 46247 11815
rect 41705 11713 41739 11747
rect 44741 11713 44775 11747
rect 45477 11713 45511 11747
rect 44925 11645 44959 11679
rect 45661 11577 45695 11611
rect 41521 11509 41555 11543
rect 46305 11509 46339 11543
rect 13001 11305 13035 11339
rect 13645 11169 13679 11203
rect 13369 11101 13403 11135
rect 14473 11101 14507 11135
rect 47961 11101 47995 11135
rect 49157 11101 49191 11135
rect 12449 11033 12483 11067
rect 13461 11033 13495 11067
rect 46305 11033 46339 11067
rect 46489 11033 46523 11067
rect 24409 10693 24443 10727
rect 40877 10625 40911 10659
rect 47961 10625 47995 10659
rect 49157 10557 49191 10591
rect 24593 10489 24627 10523
rect 40693 10421 40727 10455
rect 28733 10013 28767 10047
rect 31861 10013 31895 10047
rect 47961 10013 47995 10047
rect 28917 9945 28951 9979
rect 49157 9945 49191 9979
rect 31953 9877 31987 9911
rect 32413 9605 32447 9639
rect 36001 9605 36035 9639
rect 46213 9537 46247 9571
rect 47961 9537 47995 9571
rect 49157 9469 49191 9503
rect 32597 9401 32631 9435
rect 36185 9401 36219 9435
rect 46029 9333 46063 9367
rect 46029 8925 46063 8959
rect 46213 8857 46247 8891
rect 36553 8517 36587 8551
rect 37933 8517 37967 8551
rect 45753 8517 45787 8551
rect 9137 8449 9171 8483
rect 47961 8449 47995 8483
rect 9413 8381 9447 8415
rect 11161 8381 11195 8415
rect 36737 8381 36771 8415
rect 49157 8381 49191 8415
rect 38117 8313 38151 8347
rect 45937 8313 45971 8347
rect 47961 7837 47995 7871
rect 49157 7769 49191 7803
rect 35817 7429 35851 7463
rect 37565 7361 37599 7395
rect 47961 7361 47995 7395
rect 49157 7293 49191 7327
rect 37749 7225 37783 7259
rect 35909 7157 35943 7191
rect 37749 6749 37783 6783
rect 47409 6749 47443 6783
rect 47961 6749 47995 6783
rect 37565 6681 37599 6715
rect 38301 6681 38335 6715
rect 38485 6681 38519 6715
rect 49157 6681 49191 6715
rect 47225 6613 47259 6647
rect 48697 6273 48731 6307
rect 48789 6069 48823 6103
rect 47961 5661 47995 5695
rect 49157 5661 49191 5695
rect 29469 5185 29503 5219
rect 30113 5185 30147 5219
rect 30205 4981 30239 5015
rect 49341 4981 49375 5015
rect 47961 4573 47995 4607
rect 49157 4505 49191 4539
rect 33977 4097 34011 4131
rect 39129 4097 39163 4131
rect 43545 4097 43579 4131
rect 46029 4097 46063 4131
rect 48789 4097 48823 4131
rect 34437 4029 34471 4063
rect 39589 4029 39623 4063
rect 44005 4029 44039 4063
rect 48513 4029 48547 4063
rect 45845 3893 45879 3927
rect 1593 3689 1627 3723
rect 25053 3553 25087 3587
rect 30205 3553 30239 3587
rect 32045 3553 32079 3587
rect 35357 3553 35391 3587
rect 37197 3553 37231 3587
rect 40509 3553 40543 3587
rect 42349 3553 42383 3587
rect 45661 3553 45695 3587
rect 1777 3485 1811 3519
rect 24593 3485 24627 3519
rect 29745 3485 29779 3519
rect 31585 3485 31619 3519
rect 34897 3485 34931 3519
rect 36737 3485 36771 3519
rect 40049 3485 40083 3519
rect 41889 3485 41923 3519
rect 45201 3485 45235 3519
rect 48145 3485 48179 3519
rect 49157 3417 49191 3451
rect 6929 3145 6963 3179
rect 12817 3145 12851 3179
rect 14289 3145 14323 3179
rect 17969 3145 18003 3179
rect 4077 3077 4111 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 3893 3009 3927 3043
rect 5273 3009 5307 3043
rect 6837 3009 6871 3043
rect 10425 3009 10459 3043
rect 12725 3009 12759 3043
rect 14105 3009 14139 3043
rect 17785 3009 17819 3043
rect 19533 3009 19567 3043
rect 20913 3009 20947 3043
rect 22293 3009 22327 3043
rect 23397 3009 23431 3043
rect 25145 3009 25179 3043
rect 27353 3009 27387 3043
rect 29193 3009 29227 3043
rect 32505 3009 32539 3043
rect 34345 3009 34379 3043
rect 37657 3009 37691 3043
rect 39313 3009 39347 3043
rect 42625 3009 42659 3043
rect 44465 3009 44499 3043
rect 46673 3009 46707 3043
rect 47961 3009 47995 3043
rect 19257 2941 19291 2975
rect 20637 2941 20671 2975
rect 22017 2941 22051 2975
rect 23765 2941 23799 2975
rect 25605 2941 25639 2975
rect 27813 2941 27847 2975
rect 29653 2941 29687 2975
rect 32781 2941 32815 2975
rect 34621 2941 34655 2975
rect 37933 2941 37967 2975
rect 39773 2941 39807 2975
rect 43085 2941 43119 2975
rect 44925 2941 44959 2975
rect 46397 2941 46431 2975
rect 48421 2941 48455 2975
rect 1777 2873 1811 2907
rect 2329 2873 2363 2907
rect 5457 2873 5491 2907
rect 10609 2873 10643 2907
rect 7573 2601 7607 2635
rect 14565 2601 14599 2635
rect 46765 2601 46799 2635
rect 9505 2533 9539 2567
rect 20085 2533 20119 2567
rect 4905 2465 4939 2499
rect 18061 2465 18095 2499
rect 20637 2465 20671 2499
rect 23121 2465 23155 2499
rect 25789 2465 25823 2499
rect 27629 2465 27663 2499
rect 30205 2465 30239 2499
rect 32781 2465 32815 2499
rect 37933 2465 37967 2499
rect 40509 2465 40543 2499
rect 43085 2465 43119 2499
rect 48329 2465 48363 2499
rect 2145 2397 2179 2431
rect 7297 2397 7331 2431
rect 8585 2397 8619 2431
rect 10241 2397 10275 2431
rect 12357 2397 12391 2431
rect 14381 2397 14415 2431
rect 17509 2397 17543 2431
rect 18337 2397 18371 2431
rect 19809 2397 19843 2431
rect 20913 2397 20947 2431
rect 22661 2397 22695 2431
rect 25237 2397 25271 2431
rect 27169 2397 27203 2431
rect 29929 2397 29963 2431
rect 32321 2397 32355 2431
rect 34897 2397 34931 2431
rect 37473 2397 37507 2431
rect 40049 2397 40083 2431
rect 42625 2397 42659 2431
rect 47777 2397 47811 2431
rect 3065 2329 3099 2363
rect 4629 2329 4663 2363
rect 5641 2329 5675 2363
rect 6009 2329 6043 2363
rect 8217 2329 8251 2363
rect 9229 2329 9263 2363
rect 10793 2329 10827 2363
rect 11161 2329 11195 2363
rect 11989 2329 12023 2363
rect 13369 2329 13403 2363
rect 15209 2329 15243 2363
rect 15945 2329 15979 2363
rect 16313 2329 16347 2363
rect 17141 2329 17175 2363
rect 35817 2329 35851 2363
rect 45477 2329 45511 2363
rect 2421 2261 2455 2295
rect 3341 2261 3375 2295
rect 10057 2261 10091 2295
rect 13645 2261 13679 2295
rect 15301 2261 15335 2295
<< metal1 >>
rect 382 55700 388 55752
rect 440 55740 446 55752
rect 2866 55740 2872 55752
rect 440 55712 2872 55740
rect 440 55700 446 55712
rect 2866 55700 2872 55712
rect 2924 55700 2930 55752
rect 1104 54426 49864 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 27950 54426
rect 28002 54374 28014 54426
rect 28066 54374 28078 54426
rect 28130 54374 28142 54426
rect 28194 54374 28206 54426
rect 28258 54374 37950 54426
rect 38002 54374 38014 54426
rect 38066 54374 38078 54426
rect 38130 54374 38142 54426
rect 38194 54374 38206 54426
rect 38258 54374 47950 54426
rect 48002 54374 48014 54426
rect 48066 54374 48078 54426
rect 48130 54374 48142 54426
rect 48194 54374 48206 54426
rect 48258 54374 49864 54426
rect 1104 54352 49864 54374
rect 10042 54312 10048 54324
rect 4816 54284 10048 54312
rect 3237 54247 3295 54253
rect 3237 54213 3249 54247
rect 3283 54244 3295 54247
rect 3326 54244 3332 54256
rect 3283 54216 3332 54244
rect 3283 54213 3295 54216
rect 3237 54207 3295 54213
rect 3326 54204 3332 54216
rect 3384 54204 3390 54256
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54145 2283 54179
rect 2225 54139 2283 54145
rect 2240 54108 2268 54139
rect 2774 54136 2780 54188
rect 2832 54176 2838 54188
rect 4816 54185 4844 54284
rect 10042 54272 10048 54284
rect 10100 54272 10106 54324
rect 28902 54272 28908 54324
rect 28960 54312 28966 54324
rect 31573 54315 31631 54321
rect 31573 54312 31585 54315
rect 28960 54284 31585 54312
rect 28960 54272 28966 54284
rect 31573 54281 31585 54284
rect 31619 54281 31631 54315
rect 31573 54275 31631 54281
rect 37734 54272 37740 54324
rect 37792 54312 37798 54324
rect 41509 54315 41567 54321
rect 41509 54312 41521 54315
rect 37792 54284 41521 54312
rect 37792 54272 37798 54284
rect 41509 54281 41521 54284
rect 41555 54281 41567 54315
rect 41509 54275 41567 54281
rect 5813 54247 5871 54253
rect 5813 54213 5825 54247
rect 5859 54244 5871 54247
rect 6270 54244 6276 54256
rect 5859 54216 6276 54244
rect 5859 54213 5871 54216
rect 5813 54207 5871 54213
rect 6270 54204 6276 54216
rect 6328 54204 6334 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 8478 54244 8484 54256
rect 8435 54216 8484 54244
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 8478 54204 8484 54216
rect 8536 54204 8542 54256
rect 10965 54247 11023 54253
rect 9416 54216 9904 54244
rect 4157 54179 4215 54185
rect 4157 54176 4169 54179
rect 2832 54148 4169 54176
rect 2832 54136 2838 54148
rect 4157 54145 4169 54148
rect 4203 54145 4215 54179
rect 4157 54139 4215 54145
rect 4801 54179 4859 54185
rect 4801 54145 4813 54179
rect 4847 54145 4859 54179
rect 4801 54139 4859 54145
rect 7377 54179 7435 54185
rect 7377 54145 7389 54179
rect 7423 54176 7435 54179
rect 9416 54176 9444 54216
rect 7423 54148 9444 54176
rect 9769 54179 9827 54185
rect 7423 54145 7435 54148
rect 7377 54139 7435 54145
rect 9769 54145 9781 54179
rect 9815 54145 9827 54179
rect 9876 54176 9904 54216
rect 10965 54213 10977 54247
rect 11011 54244 11023 54247
rect 11422 54244 11428 54256
rect 11011 54216 11428 54244
rect 11011 54213 11023 54216
rect 10965 54207 11023 54213
rect 11422 54204 11428 54216
rect 11480 54204 11486 54256
rect 13541 54247 13599 54253
rect 13541 54213 13553 54247
rect 13587 54244 13599 54247
rect 13630 54244 13636 54256
rect 13587 54216 13636 54244
rect 13587 54213 13599 54216
rect 13541 54207 13599 54213
rect 13630 54204 13636 54216
rect 13688 54204 13694 54256
rect 16117 54247 16175 54253
rect 16117 54213 16129 54247
rect 16163 54244 16175 54247
rect 16574 54244 16580 54256
rect 16163 54216 16580 54244
rect 16163 54213 16175 54216
rect 16117 54207 16175 54213
rect 16574 54204 16580 54216
rect 16632 54204 16638 54256
rect 18693 54247 18751 54253
rect 18693 54213 18705 54247
rect 18739 54244 18751 54247
rect 18782 54244 18788 54256
rect 18739 54216 18788 54244
rect 18739 54213 18751 54216
rect 18693 54207 18751 54213
rect 18782 54204 18788 54216
rect 18840 54204 18846 54256
rect 20990 54204 20996 54256
rect 21048 54204 21054 54256
rect 24670 54204 24676 54256
rect 24728 54244 24734 54256
rect 24857 54247 24915 54253
rect 24857 54244 24869 54247
rect 24728 54216 24869 54244
rect 24728 54204 24734 54216
rect 24857 54213 24869 54216
rect 24903 54213 24915 54247
rect 24857 54207 24915 54213
rect 28350 54204 28356 54256
rect 28408 54244 28414 54256
rect 28721 54247 28779 54253
rect 28721 54244 28733 54247
rect 28408 54216 28733 54244
rect 28408 54204 28414 54216
rect 28721 54213 28733 54216
rect 28767 54213 28779 54247
rect 28721 54207 28779 54213
rect 32766 54204 32772 54256
rect 32824 54244 32830 54256
rect 32953 54247 33011 54253
rect 32953 54244 32965 54247
rect 32824 54216 32965 54244
rect 32824 54204 32830 54216
rect 32953 54213 32965 54216
rect 32999 54213 33011 54247
rect 32953 54207 33011 54213
rect 33502 54204 33508 54256
rect 33560 54244 33566 54256
rect 33689 54247 33747 54253
rect 33689 54244 33701 54247
rect 33560 54216 33701 54244
rect 33560 54204 33566 54216
rect 33689 54213 33701 54216
rect 33735 54213 33747 54247
rect 33689 54207 33747 54213
rect 37182 54204 37188 54256
rect 37240 54244 37246 54256
rect 37553 54247 37611 54253
rect 37553 54244 37565 54247
rect 37240 54216 37565 54244
rect 37240 54204 37246 54216
rect 37553 54213 37565 54216
rect 37599 54213 37611 54247
rect 37553 54207 37611 54213
rect 42334 54204 42340 54256
rect 42392 54244 42398 54256
rect 42705 54247 42763 54253
rect 42705 54244 42717 54247
rect 42392 54216 42717 54244
rect 42392 54204 42398 54216
rect 42705 54213 42717 54216
rect 42751 54213 42763 54247
rect 42705 54207 42763 54213
rect 11698 54176 11704 54188
rect 9876 54148 11704 54176
rect 9769 54139 9827 54145
rect 2240 54080 6914 54108
rect 3970 53932 3976 53984
rect 4028 53932 4034 53984
rect 6886 53972 6914 54080
rect 9784 54040 9812 54139
rect 11698 54136 11704 54148
rect 11756 54136 11762 54188
rect 12529 54179 12587 54185
rect 12529 54145 12541 54179
rect 12575 54176 12587 54179
rect 14550 54176 14556 54188
rect 12575 54148 14556 54176
rect 12575 54145 12587 54148
rect 12529 54139 12587 54145
rect 14550 54136 14556 54148
rect 14608 54136 14614 54188
rect 15105 54179 15163 54185
rect 15105 54145 15117 54179
rect 15151 54145 15163 54179
rect 15105 54139 15163 54145
rect 15120 54108 15148 54139
rect 17678 54136 17684 54188
rect 17736 54136 17742 54188
rect 20257 54179 20315 54185
rect 20257 54145 20269 54179
rect 20303 54176 20315 54179
rect 20346 54176 20352 54188
rect 20303 54148 20352 54176
rect 20303 54145 20315 54148
rect 20257 54139 20315 54145
rect 20346 54136 20352 54148
rect 20404 54136 20410 54188
rect 22738 54136 22744 54188
rect 22796 54136 22802 54188
rect 25406 54136 25412 54188
rect 25464 54176 25470 54188
rect 25501 54179 25559 54185
rect 25501 54176 25513 54179
rect 25464 54148 25513 54176
rect 25464 54136 25470 54148
rect 25501 54145 25513 54148
rect 25547 54145 25559 54179
rect 25501 54139 25559 54145
rect 26234 54136 26240 54188
rect 26292 54176 26298 54188
rect 26421 54179 26479 54185
rect 26421 54176 26433 54179
rect 26292 54148 26433 54176
rect 26292 54136 26298 54148
rect 26421 54145 26433 54148
rect 26467 54145 26479 54179
rect 26421 54139 26479 54145
rect 26878 54136 26884 54188
rect 26936 54176 26942 54188
rect 27157 54179 27215 54185
rect 27157 54176 27169 54179
rect 26936 54148 27169 54176
rect 26936 54136 26942 54148
rect 27157 54145 27169 54148
rect 27203 54145 27215 54179
rect 27157 54139 27215 54145
rect 27614 54136 27620 54188
rect 27672 54176 27678 54188
rect 27893 54179 27951 54185
rect 27893 54176 27905 54179
rect 27672 54148 27905 54176
rect 27672 54136 27678 54148
rect 27893 54145 27905 54148
rect 27939 54145 27951 54179
rect 27893 54139 27951 54145
rect 29822 54136 29828 54188
rect 29880 54176 29886 54188
rect 29917 54179 29975 54185
rect 29917 54176 29929 54179
rect 29880 54148 29929 54176
rect 29880 54136 29886 54148
rect 29917 54145 29929 54148
rect 29963 54145 29975 54179
rect 29917 54139 29975 54145
rect 30558 54136 30564 54188
rect 30616 54176 30622 54188
rect 30653 54179 30711 54185
rect 30653 54176 30665 54179
rect 30616 54148 30665 54176
rect 30616 54136 30622 54148
rect 30653 54145 30665 54148
rect 30699 54145 30711 54179
rect 30653 54139 30711 54145
rect 31294 54136 31300 54188
rect 31352 54176 31358 54188
rect 31389 54179 31447 54185
rect 31389 54176 31401 54179
rect 31352 54148 31401 54176
rect 31352 54136 31358 54148
rect 31389 54145 31401 54148
rect 31435 54145 31447 54179
rect 31389 54139 31447 54145
rect 34238 54136 34244 54188
rect 34296 54176 34302 54188
rect 34885 54179 34943 54185
rect 34885 54176 34897 54179
rect 34296 54148 34897 54176
rect 34296 54136 34302 54148
rect 34885 54145 34897 54148
rect 34931 54145 34943 54179
rect 34885 54139 34943 54145
rect 35710 54136 35716 54188
rect 35768 54176 35774 54188
rect 35805 54179 35863 54185
rect 35805 54176 35817 54179
rect 35768 54148 35817 54176
rect 35768 54136 35774 54148
rect 35805 54145 35817 54148
rect 35851 54145 35863 54179
rect 35805 54139 35863 54145
rect 36446 54136 36452 54188
rect 36504 54176 36510 54188
rect 36541 54179 36599 54185
rect 36541 54176 36553 54179
rect 36504 54148 36553 54176
rect 36504 54136 36510 54148
rect 36541 54145 36553 54148
rect 36587 54145 36599 54179
rect 36541 54139 36599 54145
rect 38654 54136 38660 54188
rect 38712 54176 38718 54188
rect 38749 54179 38807 54185
rect 38749 54176 38761 54179
rect 38712 54148 38761 54176
rect 38712 54136 38718 54148
rect 38749 54145 38761 54148
rect 38795 54145 38807 54179
rect 38749 54139 38807 54145
rect 39390 54136 39396 54188
rect 39448 54176 39454 54188
rect 40037 54179 40095 54185
rect 40037 54176 40049 54179
rect 39448 54148 40049 54176
rect 39448 54136 39454 54148
rect 40037 54145 40049 54148
rect 40083 54145 40095 54179
rect 40037 54139 40095 54145
rect 40126 54136 40132 54188
rect 40184 54176 40190 54188
rect 40773 54179 40831 54185
rect 40773 54176 40785 54179
rect 40184 54148 40785 54176
rect 40184 54136 40190 54148
rect 40773 54145 40785 54148
rect 40819 54145 40831 54179
rect 40773 54139 40831 54145
rect 40862 54136 40868 54188
rect 40920 54176 40926 54188
rect 41693 54179 41751 54185
rect 41693 54176 41705 54179
rect 40920 54148 41705 54176
rect 40920 54136 40926 54148
rect 41693 54145 41705 54148
rect 41739 54145 41751 54179
rect 41693 54139 41751 54145
rect 43070 54136 43076 54188
rect 43128 54176 43134 54188
rect 43717 54179 43775 54185
rect 43717 54176 43729 54179
rect 43128 54148 43729 54176
rect 43128 54136 43134 54148
rect 43717 54145 43729 54148
rect 43763 54145 43775 54179
rect 43717 54139 43775 54145
rect 44082 54136 44088 54188
rect 44140 54176 44146 54188
rect 44361 54179 44419 54185
rect 44361 54176 44373 54179
rect 44140 54148 44373 54176
rect 44140 54136 44146 54148
rect 44361 54145 44373 54148
rect 44407 54145 44419 54179
rect 44361 54139 44419 54145
rect 44542 54136 44548 54188
rect 44600 54176 44606 54188
rect 45373 54179 45431 54185
rect 45373 54176 45385 54179
rect 44600 54148 45385 54176
rect 44600 54136 44606 54148
rect 45373 54145 45385 54148
rect 45419 54145 45431 54179
rect 45373 54139 45431 54145
rect 47854 54136 47860 54188
rect 47912 54176 47918 54188
rect 47949 54179 48007 54185
rect 47949 54176 47961 54179
rect 47912 54148 47961 54176
rect 47912 54136 47918 54148
rect 47949 54145 47961 54148
rect 47995 54145 48007 54179
rect 47949 54139 48007 54145
rect 20162 54108 20168 54120
rect 15120 54080 20168 54108
rect 20162 54068 20168 54080
rect 20220 54068 20226 54120
rect 22462 54068 22468 54120
rect 22520 54108 22526 54120
rect 23017 54111 23075 54117
rect 23017 54108 23029 54111
rect 22520 54080 23029 54108
rect 22520 54068 22526 54080
rect 23017 54077 23029 54080
rect 23063 54077 23075 54111
rect 23017 54071 23075 54077
rect 42981 54111 43039 54117
rect 42981 54077 42993 54111
rect 43027 54108 43039 54111
rect 43990 54108 43996 54120
rect 43027 54080 43996 54108
rect 43027 54077 43039 54080
rect 42981 54071 43039 54077
rect 43990 54068 43996 54080
rect 44048 54068 44054 54120
rect 48222 54068 48228 54120
rect 48280 54108 48286 54120
rect 48409 54111 48467 54117
rect 48409 54108 48421 54111
rect 48280 54080 48421 54108
rect 48280 54068 48286 54080
rect 48409 54077 48421 54080
rect 48455 54077 48467 54111
rect 48409 54071 48467 54077
rect 14642 54040 14648 54052
rect 9784 54012 14648 54040
rect 14642 54000 14648 54012
rect 14700 54000 14706 54052
rect 25041 54043 25099 54049
rect 25041 54009 25053 54043
rect 25087 54040 25099 54043
rect 25222 54040 25228 54052
rect 25087 54012 25228 54040
rect 25087 54009 25099 54012
rect 25041 54003 25099 54009
rect 25222 54000 25228 54012
rect 25280 54000 25286 54052
rect 28905 54043 28963 54049
rect 28905 54009 28917 54043
rect 28951 54040 28963 54043
rect 29638 54040 29644 54052
rect 28951 54012 29644 54040
rect 28951 54009 28963 54012
rect 28905 54003 28963 54009
rect 29638 54000 29644 54012
rect 29696 54000 29702 54052
rect 33137 54043 33195 54049
rect 33137 54009 33149 54043
rect 33183 54040 33195 54043
rect 33410 54040 33416 54052
rect 33183 54012 33416 54040
rect 33183 54009 33195 54012
rect 33137 54003 33195 54009
rect 33410 54000 33416 54012
rect 33468 54000 33474 54052
rect 33873 54043 33931 54049
rect 33873 54009 33885 54043
rect 33919 54040 33931 54043
rect 33962 54040 33968 54052
rect 33919 54012 33968 54040
rect 33919 54009 33931 54012
rect 33873 54003 33931 54009
rect 33962 54000 33968 54012
rect 34020 54000 34026 54052
rect 40310 54000 40316 54052
rect 40368 54040 40374 54052
rect 40368 54012 41644 54040
rect 40368 54000 40374 54012
rect 12342 53972 12348 53984
rect 6886 53944 12348 53972
rect 12342 53932 12348 53944
rect 12400 53932 12406 53984
rect 25685 53975 25743 53981
rect 25685 53941 25697 53975
rect 25731 53972 25743 53975
rect 26050 53972 26056 53984
rect 25731 53944 26056 53972
rect 25731 53941 25743 53944
rect 25685 53935 25743 53941
rect 26050 53932 26056 53944
rect 26108 53932 26114 53984
rect 26234 53932 26240 53984
rect 26292 53932 26298 53984
rect 27341 53975 27399 53981
rect 27341 53941 27353 53975
rect 27387 53972 27399 53975
rect 27430 53972 27436 53984
rect 27387 53944 27436 53972
rect 27387 53941 27399 53944
rect 27341 53935 27399 53941
rect 27430 53932 27436 53944
rect 27488 53932 27494 53984
rect 28077 53975 28135 53981
rect 28077 53941 28089 53975
rect 28123 53972 28135 53975
rect 28534 53972 28540 53984
rect 28123 53944 28540 53972
rect 28123 53941 28135 53944
rect 28077 53935 28135 53941
rect 28534 53932 28540 53944
rect 28592 53932 28598 53984
rect 30098 53932 30104 53984
rect 30156 53932 30162 53984
rect 30466 53932 30472 53984
rect 30524 53972 30530 53984
rect 30837 53975 30895 53981
rect 30837 53972 30849 53975
rect 30524 53944 30849 53972
rect 30524 53932 30530 53944
rect 30837 53941 30849 53944
rect 30883 53941 30895 53975
rect 30837 53935 30895 53941
rect 35069 53975 35127 53981
rect 35069 53941 35081 53975
rect 35115 53972 35127 53975
rect 35250 53972 35256 53984
rect 35115 53944 35256 53972
rect 35115 53941 35127 53944
rect 35069 53935 35127 53941
rect 35250 53932 35256 53944
rect 35308 53932 35314 53984
rect 35989 53975 36047 53981
rect 35989 53941 36001 53975
rect 36035 53972 36047 53975
rect 36538 53972 36544 53984
rect 36035 53944 36544 53972
rect 36035 53941 36047 53944
rect 35989 53935 36047 53941
rect 36538 53932 36544 53944
rect 36596 53932 36602 53984
rect 36725 53975 36783 53981
rect 36725 53941 36737 53975
rect 36771 53972 36783 53975
rect 37182 53972 37188 53984
rect 36771 53944 37188 53972
rect 36771 53941 36783 53944
rect 36725 53935 36783 53941
rect 37182 53932 37188 53944
rect 37240 53932 37246 53984
rect 37642 53932 37648 53984
rect 37700 53932 37706 53984
rect 38930 53932 38936 53984
rect 38988 53932 38994 53984
rect 40221 53975 40279 53981
rect 40221 53941 40233 53975
rect 40267 53972 40279 53975
rect 40402 53972 40408 53984
rect 40267 53944 40408 53972
rect 40267 53941 40279 53944
rect 40221 53935 40279 53941
rect 40402 53932 40408 53944
rect 40460 53932 40466 53984
rect 40957 53975 41015 53981
rect 40957 53941 40969 53975
rect 41003 53972 41015 53975
rect 41046 53972 41052 53984
rect 41003 53944 41052 53972
rect 41003 53941 41015 53944
rect 40957 53935 41015 53941
rect 41046 53932 41052 53944
rect 41104 53932 41110 53984
rect 41616 53972 41644 54012
rect 43438 54000 43444 54052
rect 43496 54040 43502 54052
rect 44177 54043 44235 54049
rect 44177 54040 44189 54043
rect 43496 54012 44189 54040
rect 43496 54000 43502 54012
rect 44177 54009 44189 54012
rect 44223 54009 44235 54043
rect 44177 54003 44235 54009
rect 43533 53975 43591 53981
rect 43533 53972 43545 53975
rect 41616 53944 43545 53972
rect 43533 53941 43545 53944
rect 43579 53941 43591 53975
rect 43533 53935 43591 53941
rect 45186 53932 45192 53984
rect 45244 53932 45250 53984
rect 1104 53882 49864 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 32950 53882
rect 33002 53830 33014 53882
rect 33066 53830 33078 53882
rect 33130 53830 33142 53882
rect 33194 53830 33206 53882
rect 33258 53830 42950 53882
rect 43002 53830 43014 53882
rect 43066 53830 43078 53882
rect 43130 53830 43142 53882
rect 43194 53830 43206 53882
rect 43258 53830 49864 53882
rect 1104 53808 49864 53830
rect 15838 53660 15844 53712
rect 15896 53660 15902 53712
rect 23661 53703 23719 53709
rect 23661 53669 23673 53703
rect 23707 53700 23719 53703
rect 27062 53700 27068 53712
rect 23707 53672 27068 53700
rect 23707 53669 23719 53672
rect 23661 53663 23719 53669
rect 27062 53660 27068 53672
rect 27120 53660 27126 53712
rect 1854 53592 1860 53644
rect 1912 53632 1918 53644
rect 2409 53635 2467 53641
rect 2409 53632 2421 53635
rect 1912 53604 2421 53632
rect 1912 53592 1918 53604
rect 2409 53601 2421 53604
rect 2455 53601 2467 53635
rect 2409 53595 2467 53601
rect 5534 53592 5540 53644
rect 5592 53632 5598 53644
rect 5721 53635 5779 53641
rect 5721 53632 5733 53635
rect 5592 53604 5733 53632
rect 5592 53592 5598 53604
rect 5721 53601 5733 53604
rect 5767 53601 5779 53635
rect 5721 53595 5779 53601
rect 7006 53592 7012 53644
rect 7064 53632 7070 53644
rect 7561 53635 7619 53641
rect 7561 53632 7573 53635
rect 7064 53604 7573 53632
rect 7064 53592 7070 53604
rect 7561 53601 7573 53604
rect 7607 53601 7619 53635
rect 7561 53595 7619 53601
rect 10686 53592 10692 53644
rect 10744 53632 10750 53644
rect 10873 53635 10931 53641
rect 10873 53632 10885 53635
rect 10744 53604 10885 53632
rect 10744 53592 10750 53604
rect 10873 53601 10885 53604
rect 10919 53601 10931 53635
rect 10873 53595 10931 53601
rect 12158 53592 12164 53644
rect 12216 53632 12222 53644
rect 12713 53635 12771 53641
rect 12713 53632 12725 53635
rect 12216 53604 12725 53632
rect 12216 53592 12222 53604
rect 12713 53601 12725 53604
rect 12759 53601 12771 53635
rect 15856 53632 15884 53660
rect 16117 53635 16175 53641
rect 16117 53632 16129 53635
rect 15856 53604 16129 53632
rect 12713 53595 12771 53601
rect 16117 53601 16129 53604
rect 16163 53601 16175 53635
rect 16117 53595 16175 53601
rect 18322 53592 18328 53644
rect 18380 53592 18386 53644
rect 20254 53592 20260 53644
rect 20312 53632 20318 53644
rect 20441 53635 20499 53641
rect 20441 53632 20453 53635
rect 20312 53604 20453 53632
rect 20312 53592 20318 53604
rect 20441 53601 20453 53604
rect 20487 53601 20499 53635
rect 20441 53595 20499 53601
rect 21726 53592 21732 53644
rect 21784 53632 21790 53644
rect 22281 53635 22339 53641
rect 22281 53632 22293 53635
rect 21784 53604 22293 53632
rect 21784 53592 21790 53604
rect 22281 53601 22293 53604
rect 22327 53601 22339 53635
rect 22281 53595 22339 53601
rect 46750 53592 46756 53644
rect 46808 53632 46814 53644
rect 47305 53635 47363 53641
rect 47305 53632 47317 53635
rect 46808 53604 47317 53632
rect 46808 53592 46814 53604
rect 47305 53601 47317 53604
rect 47351 53601 47363 53635
rect 47305 53595 47363 53601
rect 2133 53567 2191 53573
rect 2133 53533 2145 53567
rect 2179 53533 2191 53567
rect 2133 53527 2191 53533
rect 5445 53567 5503 53573
rect 5445 53533 5457 53567
rect 5491 53564 5503 53567
rect 7285 53567 7343 53573
rect 5491 53536 6914 53564
rect 5491 53533 5503 53536
rect 5445 53527 5503 53533
rect 2148 53496 2176 53527
rect 6270 53496 6276 53508
rect 2148 53468 6276 53496
rect 6270 53456 6276 53468
rect 6328 53456 6334 53508
rect 6886 53496 6914 53536
rect 7285 53533 7297 53567
rect 7331 53564 7343 53567
rect 8938 53564 8944 53576
rect 7331 53536 8944 53564
rect 7331 53533 7343 53536
rect 7285 53527 7343 53533
rect 8938 53524 8944 53536
rect 8996 53524 9002 53576
rect 10410 53524 10416 53576
rect 10468 53524 10474 53576
rect 12345 53567 12403 53573
rect 12345 53533 12357 53567
rect 12391 53564 12403 53567
rect 14734 53564 14740 53576
rect 12391 53536 14740 53564
rect 12391 53533 12403 53536
rect 12345 53527 12403 53533
rect 14734 53524 14740 53536
rect 14792 53524 14798 53576
rect 15841 53567 15899 53573
rect 15841 53533 15853 53567
rect 15887 53533 15899 53567
rect 15841 53527 15899 53533
rect 17681 53567 17739 53573
rect 17681 53533 17693 53567
rect 17727 53564 17739 53567
rect 18414 53564 18420 53576
rect 17727 53536 18420 53564
rect 17727 53533 17739 53536
rect 17681 53527 17739 53533
rect 10778 53496 10784 53508
rect 6886 53468 10784 53496
rect 10778 53456 10784 53468
rect 10836 53456 10842 53508
rect 15856 53428 15884 53527
rect 18414 53524 18420 53536
rect 18472 53524 18478 53576
rect 20165 53567 20223 53573
rect 20165 53533 20177 53567
rect 20211 53533 20223 53567
rect 20165 53527 20223 53533
rect 22005 53567 22063 53573
rect 22005 53533 22017 53567
rect 22051 53564 22063 53567
rect 22830 53564 22836 53576
rect 22051 53536 22836 53564
rect 22051 53533 22063 53536
rect 22005 53527 22063 53533
rect 20180 53496 20208 53527
rect 22830 53524 22836 53536
rect 22888 53524 22894 53576
rect 23290 53524 23296 53576
rect 23348 53564 23354 53576
rect 23845 53567 23903 53573
rect 23845 53564 23857 53567
rect 23348 53536 23857 53564
rect 23348 53524 23354 53536
rect 23845 53533 23857 53536
rect 23891 53533 23903 53567
rect 23845 53527 23903 53533
rect 23934 53524 23940 53576
rect 23992 53564 23998 53576
rect 24673 53567 24731 53573
rect 24673 53564 24685 53567
rect 23992 53536 24685 53564
rect 23992 53524 23998 53536
rect 24673 53533 24685 53536
rect 24719 53533 24731 53567
rect 24673 53527 24731 53533
rect 29086 53524 29092 53576
rect 29144 53564 29150 53576
rect 29917 53567 29975 53573
rect 29917 53564 29929 53567
rect 29144 53536 29929 53564
rect 29144 53524 29150 53536
rect 29917 53533 29929 53536
rect 29963 53533 29975 53567
rect 29917 53527 29975 53533
rect 32030 53524 32036 53576
rect 32088 53564 32094 53576
rect 32309 53567 32367 53573
rect 32309 53564 32321 53567
rect 32088 53536 32321 53564
rect 32088 53524 32094 53536
rect 32309 53533 32321 53536
rect 32355 53533 32367 53567
rect 32309 53527 32367 53533
rect 34974 53524 34980 53576
rect 35032 53564 35038 53576
rect 35253 53567 35311 53573
rect 35253 53564 35265 53567
rect 35032 53536 35265 53564
rect 35032 53524 35038 53536
rect 35253 53533 35265 53536
rect 35299 53533 35311 53567
rect 35253 53527 35311 53533
rect 37826 53524 37832 53576
rect 37884 53564 37890 53576
rect 38197 53567 38255 53573
rect 38197 53564 38209 53567
rect 37884 53536 38209 53564
rect 37884 53524 37890 53536
rect 38197 53533 38209 53536
rect 38243 53533 38255 53567
rect 38197 53527 38255 53533
rect 41598 53524 41604 53576
rect 41656 53564 41662 53576
rect 41877 53567 41935 53573
rect 41877 53564 41889 53567
rect 41656 53536 41889 53564
rect 41656 53524 41662 53536
rect 41877 53533 41889 53536
rect 41923 53533 41935 53567
rect 41877 53527 41935 53533
rect 46198 53524 46204 53576
rect 46256 53564 46262 53576
rect 46845 53567 46903 53573
rect 46845 53564 46857 53567
rect 46256 53536 46857 53564
rect 46256 53524 46262 53536
rect 46845 53533 46857 53536
rect 46891 53533 46903 53567
rect 46845 53527 46903 53533
rect 22186 53496 22192 53508
rect 20180 53468 22192 53496
rect 22186 53456 22192 53468
rect 22244 53456 22250 53508
rect 24857 53499 24915 53505
rect 24857 53465 24869 53499
rect 24903 53496 24915 53499
rect 25774 53496 25780 53508
rect 24903 53468 25780 53496
rect 24903 53465 24915 53468
rect 24857 53459 24915 53465
rect 25774 53456 25780 53468
rect 25832 53456 25838 53508
rect 20438 53428 20444 53440
rect 15856 53400 20444 53428
rect 20438 53388 20444 53400
rect 20496 53388 20502 53440
rect 29730 53388 29736 53440
rect 29788 53388 29794 53440
rect 32122 53388 32128 53440
rect 32180 53388 32186 53440
rect 35069 53431 35127 53437
rect 35069 53397 35081 53431
rect 35115 53428 35127 53431
rect 35342 53428 35348 53440
rect 35115 53400 35348 53428
rect 35115 53397 35127 53400
rect 35069 53391 35127 53397
rect 35342 53388 35348 53400
rect 35400 53388 35406 53440
rect 37826 53388 37832 53440
rect 37884 53428 37890 53440
rect 38013 53431 38071 53437
rect 38013 53428 38025 53431
rect 37884 53400 38025 53428
rect 37884 53388 37890 53400
rect 38013 53397 38025 53400
rect 38059 53397 38071 53431
rect 38013 53391 38071 53397
rect 40678 53388 40684 53440
rect 40736 53428 40742 53440
rect 41693 53431 41751 53437
rect 41693 53428 41705 53431
rect 40736 53400 41705 53428
rect 40736 53388 40742 53400
rect 41693 53397 41705 53400
rect 41739 53397 41751 53431
rect 41693 53391 41751 53397
rect 1104 53338 49864 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 27950 53338
rect 28002 53286 28014 53338
rect 28066 53286 28078 53338
rect 28130 53286 28142 53338
rect 28194 53286 28206 53338
rect 28258 53286 37950 53338
rect 38002 53286 38014 53338
rect 38066 53286 38078 53338
rect 38130 53286 38142 53338
rect 38194 53286 38206 53338
rect 38258 53286 47950 53338
rect 48002 53286 48014 53338
rect 48066 53286 48078 53338
rect 48130 53286 48142 53338
rect 48194 53286 48206 53338
rect 48258 53286 49864 53338
rect 1104 53264 49864 53286
rect 46198 53184 46204 53236
rect 46256 53184 46262 53236
rect 6362 53156 6368 53168
rect 2884 53128 6368 53156
rect 934 53048 940 53100
rect 992 53088 998 53100
rect 2884 53097 2912 53128
rect 6362 53116 6368 53128
rect 6420 53116 6426 53168
rect 9858 53156 9864 53168
rect 6886 53128 9864 53156
rect 1673 53091 1731 53097
rect 1673 53088 1685 53091
rect 992 53060 1685 53088
rect 992 53048 998 53060
rect 1673 53057 1685 53060
rect 1719 53057 1731 53091
rect 1673 53051 1731 53057
rect 2869 53091 2927 53097
rect 2869 53057 2881 53091
rect 2915 53057 2927 53091
rect 2869 53051 2927 53057
rect 4801 53091 4859 53097
rect 4801 53057 4813 53091
rect 4847 53088 4859 53091
rect 6886 53088 6914 53128
rect 9858 53116 9864 53128
rect 9916 53116 9922 53168
rect 16942 53156 16948 53168
rect 13188 53128 16948 53156
rect 4847 53060 6914 53088
rect 8021 53091 8079 53097
rect 4847 53057 4859 53060
rect 4801 53051 4859 53057
rect 8021 53057 8033 53091
rect 8067 53088 8079 53091
rect 9030 53088 9036 53100
rect 8067 53060 9036 53088
rect 8067 53057 8079 53060
rect 8021 53051 8079 53057
rect 9030 53048 9036 53060
rect 9088 53048 9094 53100
rect 9766 53048 9772 53100
rect 9824 53048 9830 53100
rect 13188 53097 13216 53128
rect 16942 53116 16948 53128
rect 17000 53116 17006 53168
rect 21266 53156 21272 53168
rect 17604 53128 21272 53156
rect 13173 53091 13231 53097
rect 13173 53057 13185 53091
rect 13219 53057 13231 53091
rect 13173 53051 13231 53057
rect 15013 53091 15071 53097
rect 15013 53057 15025 53091
rect 15059 53088 15071 53091
rect 15194 53088 15200 53100
rect 15059 53060 15200 53088
rect 15059 53057 15071 53060
rect 15013 53051 15071 53057
rect 15194 53048 15200 53060
rect 15252 53048 15258 53100
rect 17604 53097 17632 53128
rect 21266 53116 21272 53128
rect 21324 53116 21330 53168
rect 49145 53159 49203 53165
rect 49145 53125 49157 53159
rect 49191 53156 49203 53159
rect 49694 53156 49700 53168
rect 49191 53128 49700 53156
rect 49191 53125 49203 53128
rect 49145 53119 49203 53125
rect 49694 53116 49700 53128
rect 49752 53116 49758 53168
rect 17589 53091 17647 53097
rect 17589 53057 17601 53091
rect 17635 53057 17647 53091
rect 17589 53051 17647 53057
rect 19610 53048 19616 53100
rect 19668 53048 19674 53100
rect 46382 53048 46388 53100
rect 46440 53048 46446 53100
rect 47670 53048 47676 53100
rect 47728 53088 47734 53100
rect 47949 53091 48007 53097
rect 47949 53088 47961 53091
rect 47728 53060 47961 53088
rect 47728 53048 47734 53060
rect 47949 53057 47961 53060
rect 47995 53057 48007 53091
rect 47949 53051 48007 53057
rect 2590 52980 2596 53032
rect 2648 53020 2654 53032
rect 3145 53023 3203 53029
rect 3145 53020 3157 53023
rect 2648 52992 3157 53020
rect 2648 52980 2654 52992
rect 3145 52989 3157 52992
rect 3191 52989 3203 53023
rect 3145 52983 3203 52989
rect 4890 52980 4896 53032
rect 4948 53020 4954 53032
rect 5077 53023 5135 53029
rect 5077 53020 5089 53023
rect 4948 52992 5089 53020
rect 4948 52980 4954 52992
rect 5077 52989 5089 52992
rect 5123 52989 5135 53023
rect 5077 52983 5135 52989
rect 7742 52980 7748 53032
rect 7800 53020 7806 53032
rect 8297 53023 8355 53029
rect 8297 53020 8309 53023
rect 7800 52992 8309 53020
rect 7800 52980 7806 52992
rect 8297 52989 8309 52992
rect 8343 52989 8355 53023
rect 8297 52983 8355 52989
rect 9950 52980 9956 53032
rect 10008 53020 10014 53032
rect 10229 53023 10287 53029
rect 10229 53020 10241 53023
rect 10008 52992 10241 53020
rect 10008 52980 10014 52992
rect 10229 52989 10241 52992
rect 10275 52989 10287 53023
rect 10229 52983 10287 52989
rect 12802 52980 12808 53032
rect 12860 53020 12866 53032
rect 13449 53023 13507 53029
rect 13449 53020 13461 53023
rect 12860 52992 13461 53020
rect 12860 52980 12866 52992
rect 13449 52989 13461 52992
rect 13495 52989 13507 53023
rect 13449 52983 13507 52989
rect 15102 52980 15108 53032
rect 15160 53020 15166 53032
rect 15381 53023 15439 53029
rect 15381 53020 15393 53023
rect 15160 52992 15393 53020
rect 15160 52980 15166 52992
rect 15381 52989 15393 52992
rect 15427 52989 15439 53023
rect 15381 52983 15439 52989
rect 17310 52980 17316 53032
rect 17368 53020 17374 53032
rect 17865 53023 17923 53029
rect 17865 53020 17877 53023
rect 17368 52992 17877 53020
rect 17368 52980 17374 52992
rect 17865 52989 17877 52992
rect 17911 52989 17923 53023
rect 17865 52983 17923 52989
rect 19518 52980 19524 53032
rect 19576 53020 19582 53032
rect 20073 53023 20131 53029
rect 20073 53020 20085 53023
rect 19576 52992 20085 53020
rect 19576 52980 19582 52992
rect 20073 52989 20085 52992
rect 20119 52989 20131 53023
rect 20073 52983 20131 52989
rect 1857 52955 1915 52961
rect 1857 52921 1869 52955
rect 1903 52952 1915 52955
rect 1946 52952 1952 52964
rect 1903 52924 1952 52952
rect 1903 52921 1915 52924
rect 1857 52915 1915 52921
rect 1946 52912 1952 52924
rect 2004 52912 2010 52964
rect 1104 52794 49864 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 32950 52794
rect 33002 52742 33014 52794
rect 33066 52742 33078 52794
rect 33130 52742 33142 52794
rect 33194 52742 33206 52794
rect 33258 52742 42950 52794
rect 43002 52742 43014 52794
rect 43066 52742 43078 52794
rect 43130 52742 43142 52794
rect 43194 52742 43206 52794
rect 43258 52742 49864 52794
rect 1104 52720 49864 52742
rect 5810 52612 5816 52624
rect 3712 52584 5816 52612
rect 1118 52504 1124 52556
rect 1176 52544 1182 52556
rect 2041 52547 2099 52553
rect 2041 52544 2053 52547
rect 1176 52516 2053 52544
rect 1176 52504 1182 52516
rect 2041 52513 2053 52516
rect 2087 52513 2099 52547
rect 2041 52507 2099 52513
rect 1765 52479 1823 52485
rect 1765 52445 1777 52479
rect 1811 52476 1823 52479
rect 3712 52476 3740 52584
rect 5810 52572 5816 52584
rect 5868 52572 5874 52624
rect 4062 52504 4068 52556
rect 4120 52544 4126 52556
rect 4617 52547 4675 52553
rect 4617 52544 4629 52547
rect 4120 52516 4629 52544
rect 4120 52504 4126 52516
rect 4617 52513 4629 52516
rect 4663 52513 4675 52547
rect 4617 52507 4675 52513
rect 9214 52504 9220 52556
rect 9272 52544 9278 52556
rect 9769 52547 9827 52553
rect 9769 52544 9781 52547
rect 9272 52516 9781 52544
rect 9272 52504 9278 52516
rect 9769 52513 9781 52516
rect 9815 52513 9827 52547
rect 9769 52507 9827 52513
rect 14366 52504 14372 52556
rect 14424 52544 14430 52556
rect 14921 52547 14979 52553
rect 14921 52544 14933 52547
rect 14424 52516 14933 52544
rect 14424 52504 14430 52516
rect 14921 52513 14933 52516
rect 14967 52513 14979 52547
rect 14921 52507 14979 52513
rect 1811 52448 3740 52476
rect 4341 52479 4399 52485
rect 1811 52445 1823 52448
rect 1765 52439 1823 52445
rect 4341 52445 4353 52479
rect 4387 52476 4399 52479
rect 9122 52476 9128 52488
rect 4387 52448 9128 52476
rect 4387 52445 4399 52448
rect 4341 52439 4399 52445
rect 9122 52436 9128 52448
rect 9180 52436 9186 52488
rect 9493 52479 9551 52485
rect 9493 52445 9505 52479
rect 9539 52476 9551 52479
rect 14458 52476 14464 52488
rect 9539 52448 14464 52476
rect 9539 52445 9551 52448
rect 9493 52439 9551 52445
rect 14458 52436 14464 52448
rect 14516 52436 14522 52488
rect 14645 52479 14703 52485
rect 14645 52445 14657 52479
rect 14691 52476 14703 52479
rect 19150 52476 19156 52488
rect 14691 52448 19156 52476
rect 14691 52445 14703 52448
rect 14645 52439 14703 52445
rect 19150 52436 19156 52448
rect 19208 52436 19214 52488
rect 1104 52250 49864 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 27950 52250
rect 28002 52198 28014 52250
rect 28066 52198 28078 52250
rect 28130 52198 28142 52250
rect 28194 52198 28206 52250
rect 28258 52198 37950 52250
rect 38002 52198 38014 52250
rect 38066 52198 38078 52250
rect 38130 52198 38142 52250
rect 38194 52198 38206 52250
rect 38258 52198 47950 52250
rect 48002 52198 48014 52250
rect 48066 52198 48078 52250
rect 48130 52198 48142 52250
rect 48194 52198 48206 52250
rect 48258 52198 49864 52250
rect 1104 52176 49864 52198
rect 22738 52096 22744 52148
rect 22796 52136 22802 52148
rect 23569 52139 23627 52145
rect 23569 52136 23581 52139
rect 22796 52108 23581 52136
rect 22796 52096 22802 52108
rect 23569 52105 23581 52108
rect 23615 52105 23627 52139
rect 23569 52099 23627 52105
rect 2777 52071 2835 52077
rect 2777 52037 2789 52071
rect 2823 52068 2835 52071
rect 2866 52068 2872 52080
rect 2823 52040 2872 52068
rect 2823 52037 2835 52040
rect 2777 52031 2835 52037
rect 2866 52028 2872 52040
rect 2924 52028 2930 52080
rect 1578 51960 1584 52012
rect 1636 51960 1642 52012
rect 23750 51960 23756 52012
rect 23808 51960 23814 52012
rect 49050 51960 49056 52012
rect 49108 51960 49114 52012
rect 49234 51756 49240 51808
rect 49292 51756 49298 51808
rect 1104 51706 49864 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 32950 51706
rect 33002 51654 33014 51706
rect 33066 51654 33078 51706
rect 33130 51654 33142 51706
rect 33194 51654 33206 51706
rect 33258 51654 42950 51706
rect 43002 51654 43014 51706
rect 43066 51654 43078 51706
rect 43130 51654 43142 51706
rect 43194 51654 43206 51706
rect 43258 51654 49864 51706
rect 1104 51632 49864 51654
rect 10042 51552 10048 51604
rect 10100 51592 10106 51604
rect 13081 51595 13139 51601
rect 13081 51592 13093 51595
rect 10100 51564 13093 51592
rect 10100 51552 10106 51564
rect 13081 51561 13093 51564
rect 13127 51561 13139 51595
rect 13081 51555 13139 51561
rect 14458 51552 14464 51604
rect 14516 51552 14522 51604
rect 22830 51552 22836 51604
rect 22888 51592 22894 51604
rect 24673 51595 24731 51601
rect 24673 51592 24685 51595
rect 22888 51564 24685 51592
rect 22888 51552 22894 51564
rect 24673 51561 24685 51564
rect 24719 51561 24731 51595
rect 24673 51555 24731 51561
rect 24857 51391 24915 51397
rect 24857 51357 24869 51391
rect 24903 51388 24915 51391
rect 26694 51388 26700 51400
rect 24903 51360 26700 51388
rect 24903 51357 24915 51360
rect 24857 51351 24915 51357
rect 26694 51348 26700 51360
rect 26752 51348 26758 51400
rect 49050 51348 49056 51400
rect 49108 51348 49114 51400
rect 12989 51323 13047 51329
rect 12989 51289 13001 51323
rect 13035 51320 13047 51323
rect 14274 51320 14280 51332
rect 13035 51292 14280 51320
rect 13035 51289 13047 51292
rect 12989 51283 13047 51289
rect 14274 51280 14280 51292
rect 14332 51280 14338 51332
rect 14369 51323 14427 51329
rect 14369 51289 14381 51323
rect 14415 51320 14427 51323
rect 15930 51320 15936 51332
rect 14415 51292 15936 51320
rect 14415 51289 14427 51292
rect 14369 51283 14427 51289
rect 15930 51280 15936 51292
rect 15988 51280 15994 51332
rect 49142 51212 49148 51264
rect 49200 51252 49206 51264
rect 49237 51255 49295 51261
rect 49237 51252 49249 51255
rect 49200 51224 49249 51252
rect 49200 51212 49206 51224
rect 49237 51221 49249 51224
rect 49283 51221 49295 51255
rect 49237 51215 49295 51221
rect 1104 51162 49864 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 27950 51162
rect 28002 51110 28014 51162
rect 28066 51110 28078 51162
rect 28130 51110 28142 51162
rect 28194 51110 28206 51162
rect 28258 51110 37950 51162
rect 38002 51110 38014 51162
rect 38066 51110 38078 51162
rect 38130 51110 38142 51162
rect 38194 51110 38206 51162
rect 38258 51110 47950 51162
rect 48002 51110 48014 51162
rect 48066 51110 48078 51162
rect 48130 51110 48142 51162
rect 48194 51110 48206 51162
rect 48258 51110 49864 51162
rect 1104 51088 49864 51110
rect 22186 51008 22192 51060
rect 22244 51008 22250 51060
rect 20346 50940 20352 50992
rect 20404 50980 20410 50992
rect 23293 50983 23351 50989
rect 23293 50980 23305 50983
rect 20404 50952 23305 50980
rect 20404 50940 20410 50952
rect 23293 50949 23305 50952
rect 23339 50949 23351 50983
rect 23293 50943 23351 50949
rect 934 50872 940 50924
rect 992 50912 998 50924
rect 1673 50915 1731 50921
rect 1673 50912 1685 50915
rect 992 50884 1685 50912
rect 992 50872 998 50884
rect 1673 50881 1685 50884
rect 1719 50881 1731 50915
rect 1673 50875 1731 50881
rect 22097 50915 22155 50921
rect 22097 50881 22109 50915
rect 22143 50912 22155 50915
rect 22738 50912 22744 50924
rect 22143 50884 22744 50912
rect 22143 50881 22155 50884
rect 22097 50875 22155 50881
rect 22738 50872 22744 50884
rect 22796 50872 22802 50924
rect 23109 50915 23167 50921
rect 23109 50881 23121 50915
rect 23155 50912 23167 50915
rect 24118 50912 24124 50924
rect 23155 50884 24124 50912
rect 23155 50881 23167 50884
rect 23109 50875 23167 50881
rect 24118 50872 24124 50884
rect 24176 50872 24182 50924
rect 48958 50872 48964 50924
rect 49016 50872 49022 50924
rect 1670 50668 1676 50720
rect 1728 50708 1734 50720
rect 1765 50711 1823 50717
rect 1765 50708 1777 50711
rect 1728 50680 1777 50708
rect 1728 50668 1734 50680
rect 1765 50677 1777 50680
rect 1811 50677 1823 50711
rect 1765 50671 1823 50677
rect 49237 50711 49295 50717
rect 49237 50677 49249 50711
rect 49283 50708 49295 50711
rect 49418 50708 49424 50720
rect 49283 50680 49424 50708
rect 49283 50677 49295 50680
rect 49237 50671 49295 50677
rect 49418 50668 49424 50680
rect 49476 50668 49482 50720
rect 1104 50618 49864 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 32950 50618
rect 33002 50566 33014 50618
rect 33066 50566 33078 50618
rect 33130 50566 33142 50618
rect 33194 50566 33206 50618
rect 33258 50566 42950 50618
rect 43002 50566 43014 50618
rect 43066 50566 43078 50618
rect 43130 50566 43142 50618
rect 43194 50566 43206 50618
rect 43258 50566 49864 50618
rect 1104 50544 49864 50566
rect 17678 50464 17684 50516
rect 17736 50504 17742 50516
rect 20257 50507 20315 50513
rect 20257 50504 20269 50507
rect 17736 50476 20269 50504
rect 17736 50464 17742 50476
rect 20257 50473 20269 50476
rect 20303 50473 20315 50507
rect 20257 50467 20315 50473
rect 49050 50260 49056 50312
rect 49108 50260 49114 50312
rect 20165 50235 20223 50241
rect 20165 50201 20177 50235
rect 20211 50232 20223 50235
rect 21818 50232 21824 50244
rect 20211 50204 21824 50232
rect 20211 50201 20223 50204
rect 20165 50195 20223 50201
rect 21818 50192 21824 50204
rect 21876 50192 21882 50244
rect 48406 50124 48412 50176
rect 48464 50164 48470 50176
rect 49237 50167 49295 50173
rect 49237 50164 49249 50167
rect 48464 50136 49249 50164
rect 48464 50124 48470 50136
rect 49237 50133 49249 50136
rect 49283 50133 49295 50167
rect 49237 50127 49295 50133
rect 1104 50074 49864 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 27950 50074
rect 28002 50022 28014 50074
rect 28066 50022 28078 50074
rect 28130 50022 28142 50074
rect 28194 50022 28206 50074
rect 28258 50022 37950 50074
rect 38002 50022 38014 50074
rect 38066 50022 38078 50074
rect 38130 50022 38142 50074
rect 38194 50022 38206 50074
rect 38258 50022 47950 50074
rect 48002 50022 48014 50074
rect 48066 50022 48078 50074
rect 48130 50022 48142 50074
rect 48194 50022 48206 50074
rect 48258 50022 49864 50074
rect 1104 50000 49864 50022
rect 12342 49920 12348 49972
rect 12400 49920 12406 49972
rect 14734 49920 14740 49972
rect 14792 49920 14798 49972
rect 12253 49895 12311 49901
rect 12253 49861 12265 49895
rect 12299 49892 12311 49895
rect 20898 49892 20904 49904
rect 12299 49864 20904 49892
rect 12299 49861 12311 49864
rect 12253 49855 12311 49861
rect 20898 49852 20904 49864
rect 20956 49852 20962 49904
rect 14645 49827 14703 49833
rect 14645 49793 14657 49827
rect 14691 49824 14703 49827
rect 16850 49824 16856 49836
rect 14691 49796 16856 49824
rect 14691 49793 14703 49796
rect 14645 49787 14703 49793
rect 16850 49784 16856 49796
rect 16908 49784 16914 49836
rect 1104 49530 49864 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 32950 49530
rect 33002 49478 33014 49530
rect 33066 49478 33078 49530
rect 33130 49478 33142 49530
rect 33194 49478 33206 49530
rect 33258 49478 42950 49530
rect 43002 49478 43014 49530
rect 43066 49478 43078 49530
rect 43130 49478 43142 49530
rect 43194 49478 43206 49530
rect 43258 49478 49864 49530
rect 1104 49456 49864 49478
rect 15194 49376 15200 49428
rect 15252 49416 15258 49428
rect 18141 49419 18199 49425
rect 18141 49416 18153 49419
rect 15252 49388 18153 49416
rect 15252 49376 15258 49388
rect 18141 49385 18153 49388
rect 18187 49385 18199 49419
rect 18141 49379 18199 49385
rect 18414 49376 18420 49428
rect 18472 49416 18478 49428
rect 20349 49419 20407 49425
rect 20349 49416 20361 49419
rect 18472 49388 20361 49416
rect 18472 49376 18478 49388
rect 20349 49385 20361 49388
rect 20395 49385 20407 49419
rect 20349 49379 20407 49385
rect 18049 49215 18107 49221
rect 18049 49181 18061 49215
rect 18095 49212 18107 49215
rect 20714 49212 20720 49224
rect 18095 49184 20720 49212
rect 18095 49181 18107 49184
rect 18049 49175 18107 49181
rect 20714 49172 20720 49184
rect 20772 49172 20778 49224
rect 49050 49172 49056 49224
rect 49108 49172 49114 49224
rect 20257 49147 20315 49153
rect 20257 49113 20269 49147
rect 20303 49144 20315 49147
rect 22094 49144 22100 49156
rect 20303 49116 22100 49144
rect 20303 49113 20315 49116
rect 20257 49107 20315 49113
rect 22094 49104 22100 49116
rect 22152 49104 22158 49156
rect 48866 49036 48872 49088
rect 48924 49076 48930 49088
rect 49237 49079 49295 49085
rect 49237 49076 49249 49079
rect 48924 49048 49249 49076
rect 48924 49036 48930 49048
rect 49237 49045 49249 49048
rect 49283 49045 49295 49079
rect 49237 49039 49295 49045
rect 1104 48986 49864 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 27950 48986
rect 28002 48934 28014 48986
rect 28066 48934 28078 48986
rect 28130 48934 28142 48986
rect 28194 48934 28206 48986
rect 28258 48934 37950 48986
rect 38002 48934 38014 48986
rect 38066 48934 38078 48986
rect 38130 48934 38142 48986
rect 38194 48934 38206 48986
rect 38258 48934 47950 48986
rect 48002 48934 48014 48986
rect 48066 48934 48078 48986
rect 48130 48934 48142 48986
rect 48194 48934 48206 48986
rect 48258 48934 49864 48986
rect 1104 48912 49864 48934
rect 49050 48696 49056 48748
rect 49108 48696 49114 48748
rect 48958 48492 48964 48544
rect 49016 48532 49022 48544
rect 49237 48535 49295 48541
rect 49237 48532 49249 48535
rect 49016 48504 49249 48532
rect 49016 48492 49022 48504
rect 49237 48501 49249 48504
rect 49283 48501 49295 48535
rect 49237 48495 49295 48501
rect 1104 48442 49864 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 32950 48442
rect 33002 48390 33014 48442
rect 33066 48390 33078 48442
rect 33130 48390 33142 48442
rect 33194 48390 33206 48442
rect 33258 48390 42950 48442
rect 43002 48390 43014 48442
rect 43066 48390 43078 48442
rect 43130 48390 43142 48442
rect 43194 48390 43206 48442
rect 43258 48390 49864 48442
rect 1104 48368 49864 48390
rect 10137 48195 10195 48201
rect 10137 48161 10149 48195
rect 10183 48192 10195 48195
rect 21082 48192 21088 48204
rect 10183 48164 21088 48192
rect 10183 48161 10195 48164
rect 10137 48155 10195 48161
rect 21082 48152 21088 48164
rect 21140 48152 21146 48204
rect 49050 48084 49056 48136
rect 49108 48084 49114 48136
rect 934 48016 940 48068
rect 992 48056 998 48068
rect 1673 48059 1731 48065
rect 1673 48056 1685 48059
rect 992 48028 1685 48056
rect 992 48016 998 48028
rect 1673 48025 1685 48028
rect 1719 48025 1731 48059
rect 1673 48019 1731 48025
rect 1854 48016 1860 48068
rect 1912 48016 1918 48068
rect 3970 48016 3976 48068
rect 4028 48056 4034 48068
rect 10413 48059 10471 48065
rect 10413 48056 10425 48059
rect 4028 48028 10425 48056
rect 4028 48016 4034 48028
rect 10413 48025 10425 48028
rect 10459 48025 10471 48059
rect 12161 48059 12219 48065
rect 11638 48028 12112 48056
rect 10413 48019 10471 48025
rect 12084 47988 12112 48028
rect 12161 48025 12173 48059
rect 12207 48056 12219 48059
rect 21910 48056 21916 48068
rect 12207 48028 21916 48056
rect 12207 48025 12219 48028
rect 12161 48019 12219 48025
rect 21910 48016 21916 48028
rect 21968 48016 21974 48068
rect 20530 47988 20536 48000
rect 12084 47960 20536 47988
rect 20530 47948 20536 47960
rect 20588 47948 20594 48000
rect 40126 47948 40132 48000
rect 40184 47988 40190 48000
rect 49237 47991 49295 47997
rect 49237 47988 49249 47991
rect 40184 47960 49249 47988
rect 40184 47948 40190 47960
rect 49237 47957 49249 47960
rect 49283 47957 49295 47991
rect 49237 47951 49295 47957
rect 1104 47898 49864 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 27950 47898
rect 28002 47846 28014 47898
rect 28066 47846 28078 47898
rect 28130 47846 28142 47898
rect 28194 47846 28206 47898
rect 28258 47846 37950 47898
rect 38002 47846 38014 47898
rect 38066 47846 38078 47898
rect 38130 47846 38142 47898
rect 38194 47846 38206 47898
rect 38258 47846 47950 47898
rect 48002 47846 48014 47898
rect 48066 47846 48078 47898
rect 48130 47846 48142 47898
rect 48194 47846 48206 47898
rect 48258 47846 49864 47898
rect 1104 47824 49864 47846
rect 23750 47744 23756 47796
rect 23808 47784 23814 47796
rect 24581 47787 24639 47793
rect 24581 47784 24593 47787
rect 23808 47756 24593 47784
rect 23808 47744 23814 47756
rect 24581 47753 24593 47756
rect 24627 47753 24639 47787
rect 24581 47747 24639 47753
rect 24765 47651 24823 47657
rect 24765 47617 24777 47651
rect 24811 47648 24823 47651
rect 25866 47648 25872 47660
rect 24811 47620 25872 47648
rect 24811 47617 24823 47620
rect 24765 47611 24823 47617
rect 25866 47608 25872 47620
rect 25924 47608 25930 47660
rect 49050 47608 49056 47660
rect 49108 47608 49114 47660
rect 48682 47404 48688 47456
rect 48740 47444 48746 47456
rect 49237 47447 49295 47453
rect 49237 47444 49249 47447
rect 48740 47416 49249 47444
rect 48740 47404 48746 47416
rect 49237 47413 49249 47416
rect 49283 47413 49295 47447
rect 49237 47407 49295 47413
rect 1104 47354 49864 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 32950 47354
rect 33002 47302 33014 47354
rect 33066 47302 33078 47354
rect 33130 47302 33142 47354
rect 33194 47302 33206 47354
rect 33258 47302 42950 47354
rect 43002 47302 43014 47354
rect 43066 47302 43078 47354
rect 43130 47302 43142 47354
rect 43194 47302 43206 47354
rect 43258 47302 49864 47354
rect 1104 47280 49864 47302
rect 1104 46810 49864 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 27950 46810
rect 28002 46758 28014 46810
rect 28066 46758 28078 46810
rect 28130 46758 28142 46810
rect 28194 46758 28206 46810
rect 28258 46758 37950 46810
rect 38002 46758 38014 46810
rect 38066 46758 38078 46810
rect 38130 46758 38142 46810
rect 38194 46758 38206 46810
rect 38258 46758 47950 46810
rect 48002 46758 48014 46810
rect 48066 46758 48078 46810
rect 48130 46758 48142 46810
rect 48194 46758 48206 46810
rect 48258 46758 49864 46810
rect 1104 46736 49864 46758
rect 1104 46266 49864 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 32950 46266
rect 33002 46214 33014 46266
rect 33066 46214 33078 46266
rect 33130 46214 33142 46266
rect 33194 46214 33206 46266
rect 33258 46214 42950 46266
rect 43002 46214 43014 46266
rect 43066 46214 43078 46266
rect 43130 46214 43142 46266
rect 43194 46214 43206 46266
rect 43258 46214 49864 46266
rect 1104 46192 49864 46214
rect 15930 46112 15936 46164
rect 15988 46152 15994 46164
rect 18417 46155 18475 46161
rect 18417 46152 18429 46155
rect 15988 46124 18429 46152
rect 15988 46112 15994 46124
rect 18417 46121 18429 46124
rect 18463 46121 18475 46155
rect 18417 46115 18475 46121
rect 26694 46112 26700 46164
rect 26752 46112 26758 46164
rect 18601 45951 18659 45957
rect 18601 45917 18613 45951
rect 18647 45948 18659 45951
rect 19705 45951 19763 45957
rect 18647 45920 19656 45948
rect 18647 45917 18659 45920
rect 18601 45911 18659 45917
rect 934 45840 940 45892
rect 992 45880 998 45892
rect 1673 45883 1731 45889
rect 1673 45880 1685 45883
rect 992 45852 1685 45880
rect 992 45840 998 45852
rect 1673 45849 1685 45852
rect 1719 45849 1731 45883
rect 1673 45843 1731 45849
rect 14274 45840 14280 45892
rect 14332 45880 14338 45892
rect 19628 45880 19656 45920
rect 19705 45917 19717 45951
rect 19751 45948 19763 45951
rect 22002 45948 22008 45960
rect 19751 45920 22008 45948
rect 19751 45917 19763 45920
rect 19705 45911 19763 45917
rect 22002 45908 22008 45920
rect 22060 45908 22066 45960
rect 26881 45951 26939 45957
rect 26881 45917 26893 45951
rect 26927 45948 26939 45951
rect 27798 45948 27804 45960
rect 26927 45920 27804 45948
rect 26927 45917 26939 45920
rect 26881 45911 26939 45917
rect 27798 45908 27804 45920
rect 27856 45908 27862 45960
rect 48133 45951 48191 45957
rect 48133 45917 48145 45951
rect 48179 45948 48191 45951
rect 48590 45948 48596 45960
rect 48179 45920 48596 45948
rect 48179 45917 48191 45920
rect 48133 45911 48191 45917
rect 48590 45908 48596 45920
rect 48648 45908 48654 45960
rect 20622 45880 20628 45892
rect 14332 45852 19564 45880
rect 19628 45852 20628 45880
rect 14332 45840 14338 45852
rect 1762 45772 1768 45824
rect 1820 45772 1826 45824
rect 19536 45821 19564 45852
rect 20622 45840 20628 45852
rect 20680 45840 20686 45892
rect 49142 45840 49148 45892
rect 49200 45840 49206 45892
rect 19521 45815 19579 45821
rect 19521 45781 19533 45815
rect 19567 45781 19579 45815
rect 19521 45775 19579 45781
rect 1104 45722 49864 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 27950 45722
rect 28002 45670 28014 45722
rect 28066 45670 28078 45722
rect 28130 45670 28142 45722
rect 28194 45670 28206 45722
rect 28258 45670 37950 45722
rect 38002 45670 38014 45722
rect 38066 45670 38078 45722
rect 38130 45670 38142 45722
rect 38194 45670 38206 45722
rect 38258 45670 47950 45722
rect 48002 45670 48014 45722
rect 48066 45670 48078 45722
rect 48130 45670 48142 45722
rect 48194 45670 48206 45722
rect 48258 45670 49864 45722
rect 1104 45648 49864 45670
rect 1762 45568 1768 45620
rect 1820 45608 1826 45620
rect 22462 45608 22468 45620
rect 1820 45580 22468 45608
rect 1820 45568 1826 45580
rect 22462 45568 22468 45580
rect 22520 45568 22526 45620
rect 48590 45568 48596 45620
rect 48648 45568 48654 45620
rect 10410 45500 10416 45552
rect 10468 45540 10474 45552
rect 15105 45543 15163 45549
rect 15105 45540 15117 45543
rect 10468 45512 15117 45540
rect 10468 45500 10474 45512
rect 15105 45509 15117 45512
rect 15151 45509 15163 45543
rect 15105 45503 15163 45509
rect 32122 45500 32128 45552
rect 32180 45540 32186 45552
rect 33873 45543 33931 45549
rect 33873 45540 33885 45543
rect 32180 45512 33885 45540
rect 32180 45500 32186 45512
rect 33873 45509 33885 45512
rect 33919 45509 33931 45543
rect 33873 45503 33931 45509
rect 46382 45500 46388 45552
rect 46440 45540 46446 45552
rect 46440 45512 48820 45540
rect 46440 45500 46446 45512
rect 14921 45475 14979 45481
rect 14921 45441 14933 45475
rect 14967 45472 14979 45475
rect 21542 45472 21548 45484
rect 14967 45444 21548 45472
rect 14967 45441 14979 45444
rect 14921 45435 14979 45441
rect 21542 45432 21548 45444
rect 21600 45432 21606 45484
rect 29730 45432 29736 45484
rect 29788 45472 29794 45484
rect 32677 45475 32735 45481
rect 32677 45472 32689 45475
rect 29788 45444 32689 45472
rect 29788 45432 29794 45444
rect 32677 45441 32689 45444
rect 32723 45441 32735 45475
rect 32677 45435 32735 45441
rect 32769 45475 32827 45481
rect 32769 45441 32781 45475
rect 32815 45472 32827 45475
rect 33410 45472 33416 45484
rect 32815 45444 33416 45472
rect 32815 45441 32827 45444
rect 32769 45435 32827 45441
rect 33410 45432 33416 45444
rect 33468 45432 33474 45484
rect 48133 45475 48191 45481
rect 48133 45441 48145 45475
rect 48179 45472 48191 45475
rect 48314 45472 48320 45484
rect 48179 45444 48320 45472
rect 48179 45441 48191 45444
rect 48133 45435 48191 45441
rect 48314 45432 48320 45444
rect 48372 45432 48378 45484
rect 48792 45481 48820 45512
rect 48777 45475 48835 45481
rect 48777 45441 48789 45475
rect 48823 45441 48835 45475
rect 48777 45435 48835 45441
rect 32858 45364 32864 45416
rect 32916 45364 32922 45416
rect 33962 45364 33968 45416
rect 34020 45364 34026 45416
rect 34146 45364 34152 45416
rect 34204 45364 34210 45416
rect 32309 45271 32367 45277
rect 32309 45237 32321 45271
rect 32355 45268 32367 45271
rect 32674 45268 32680 45280
rect 32355 45240 32680 45268
rect 32355 45237 32367 45240
rect 32309 45231 32367 45237
rect 32674 45228 32680 45240
rect 32732 45228 32738 45280
rect 33502 45228 33508 45280
rect 33560 45228 33566 45280
rect 46934 45228 46940 45280
rect 46992 45268 46998 45280
rect 47949 45271 48007 45277
rect 47949 45268 47961 45271
rect 46992 45240 47961 45268
rect 46992 45228 46998 45240
rect 47949 45237 47961 45240
rect 47995 45237 48007 45271
rect 47949 45231 48007 45237
rect 1104 45178 49864 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 32950 45178
rect 33002 45126 33014 45178
rect 33066 45126 33078 45178
rect 33130 45126 33142 45178
rect 33194 45126 33206 45178
rect 33258 45126 42950 45178
rect 43002 45126 43014 45178
rect 43066 45126 43078 45178
rect 43130 45126 43142 45178
rect 43194 45126 43206 45178
rect 43258 45126 49864 45178
rect 1104 45104 49864 45126
rect 22738 45024 22744 45076
rect 22796 45064 22802 45076
rect 22925 45067 22983 45073
rect 22925 45064 22937 45067
rect 22796 45036 22937 45064
rect 22796 45024 22802 45036
rect 22925 45033 22937 45036
rect 22971 45033 22983 45067
rect 22925 45027 22983 45033
rect 24118 45024 24124 45076
rect 24176 45064 24182 45076
rect 25041 45067 25099 45073
rect 25041 45064 25053 45067
rect 24176 45036 25053 45064
rect 24176 45024 24182 45036
rect 25041 45033 25053 45036
rect 25087 45033 25099 45067
rect 25041 45027 25099 45033
rect 34885 44999 34943 45005
rect 34885 44965 34897 44999
rect 34931 44996 34943 44999
rect 35986 44996 35992 45008
rect 34931 44968 35992 44996
rect 34931 44965 34943 44968
rect 34885 44959 34943 44965
rect 35986 44956 35992 44968
rect 36044 44956 36050 45008
rect 35342 44888 35348 44940
rect 35400 44888 35406 44940
rect 35526 44888 35532 44940
rect 35584 44888 35590 44940
rect 48777 44931 48835 44937
rect 48777 44928 48789 44931
rect 45526 44900 48789 44928
rect 23109 44863 23167 44869
rect 23109 44829 23121 44863
rect 23155 44860 23167 44863
rect 24486 44860 24492 44872
rect 23155 44832 24492 44860
rect 23155 44829 23167 44832
rect 23109 44823 23167 44829
rect 24486 44820 24492 44832
rect 24544 44820 24550 44872
rect 25225 44863 25283 44869
rect 25225 44829 25237 44863
rect 25271 44860 25283 44863
rect 27154 44860 27160 44872
rect 25271 44832 27160 44860
rect 25271 44829 25283 44832
rect 25225 44823 25283 44829
rect 27154 44820 27160 44832
rect 27212 44820 27218 44872
rect 38378 44820 38384 44872
rect 38436 44860 38442 44872
rect 45526 44860 45554 44900
rect 48777 44897 48789 44900
rect 48823 44897 48835 44931
rect 48777 44891 48835 44897
rect 38436 44832 45554 44860
rect 38436 44820 38442 44832
rect 48498 44820 48504 44872
rect 48556 44820 48562 44872
rect 35250 44684 35256 44736
rect 35308 44684 35314 44736
rect 1104 44634 49864 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 27950 44634
rect 28002 44582 28014 44634
rect 28066 44582 28078 44634
rect 28130 44582 28142 44634
rect 28194 44582 28206 44634
rect 28258 44582 37950 44634
rect 38002 44582 38014 44634
rect 38066 44582 38078 44634
rect 38130 44582 38142 44634
rect 38194 44582 38206 44634
rect 38258 44582 47950 44634
rect 48002 44582 48014 44634
rect 48066 44582 48078 44634
rect 48130 44582 48142 44634
rect 48194 44582 48206 44634
rect 48258 44582 49864 44634
rect 1104 44560 49864 44582
rect 9766 44480 9772 44532
rect 9824 44520 9830 44532
rect 14369 44523 14427 44529
rect 14369 44520 14381 44523
rect 9824 44492 14381 44520
rect 9824 44480 9830 44492
rect 14369 44489 14381 44492
rect 14415 44489 14427 44523
rect 14369 44483 14427 44489
rect 36633 44523 36691 44529
rect 36633 44489 36645 44523
rect 36679 44520 36691 44523
rect 37826 44520 37832 44532
rect 36679 44492 37832 44520
rect 36679 44489 36691 44492
rect 36633 44483 36691 44489
rect 37826 44480 37832 44492
rect 37884 44480 37890 44532
rect 39209 44523 39267 44529
rect 39209 44489 39221 44523
rect 39255 44520 39267 44523
rect 40678 44520 40684 44532
rect 39255 44492 40684 44520
rect 39255 44489 39267 44492
rect 39209 44483 39267 44489
rect 40678 44480 40684 44492
rect 40736 44480 40742 44532
rect 14277 44387 14335 44393
rect 14277 44353 14289 44387
rect 14323 44384 14335 44387
rect 14458 44384 14464 44396
rect 14323 44356 14464 44384
rect 14323 44353 14335 44356
rect 14277 44347 14335 44353
rect 14458 44344 14464 44356
rect 14516 44344 14522 44396
rect 36538 44344 36544 44396
rect 36596 44344 36602 44396
rect 37642 44344 37648 44396
rect 37700 44384 37706 44396
rect 39117 44387 39175 44393
rect 39117 44384 39129 44387
rect 37700 44356 39129 44384
rect 37700 44344 37706 44356
rect 39117 44353 39129 44356
rect 39163 44353 39175 44387
rect 39117 44347 39175 44353
rect 36817 44319 36875 44325
rect 36817 44285 36829 44319
rect 36863 44316 36875 44319
rect 36906 44316 36912 44328
rect 36863 44288 36912 44316
rect 36863 44285 36875 44288
rect 36817 44279 36875 44285
rect 36906 44276 36912 44288
rect 36964 44276 36970 44328
rect 38654 44276 38660 44328
rect 38712 44316 38718 44328
rect 39301 44319 39359 44325
rect 39301 44316 39313 44319
rect 38712 44288 39313 44316
rect 38712 44276 38718 44288
rect 39301 44285 39313 44288
rect 39347 44285 39359 44319
rect 39301 44279 39359 44285
rect 36170 44140 36176 44192
rect 36228 44140 36234 44192
rect 38746 44140 38752 44192
rect 38804 44140 38810 44192
rect 1104 44090 49864 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 32950 44090
rect 33002 44038 33014 44090
rect 33066 44038 33078 44090
rect 33130 44038 33142 44090
rect 33194 44038 33206 44090
rect 33258 44038 42950 44090
rect 43002 44038 43014 44090
rect 43066 44038 43078 44090
rect 43130 44038 43142 44090
rect 43194 44038 43206 44090
rect 43258 44038 49864 44090
rect 1104 44016 49864 44038
rect 11698 43936 11704 43988
rect 11756 43976 11762 43988
rect 13541 43979 13599 43985
rect 13541 43976 13553 43979
rect 11756 43948 13553 43976
rect 11756 43936 11762 43948
rect 13541 43945 13553 43948
rect 13587 43945 13599 43979
rect 13541 43939 13599 43945
rect 14642 43936 14648 43988
rect 14700 43976 14706 43988
rect 16209 43979 16267 43985
rect 16209 43976 16221 43979
rect 14700 43948 16221 43976
rect 14700 43936 14706 43948
rect 16209 43945 16221 43948
rect 16255 43945 16267 43979
rect 16209 43939 16267 43945
rect 16942 43936 16948 43988
rect 17000 43936 17006 43988
rect 20438 43936 20444 43988
rect 20496 43936 20502 43988
rect 21266 43936 21272 43988
rect 21324 43936 21330 43988
rect 21818 43936 21824 43988
rect 21876 43936 21882 43988
rect 28445 43979 28503 43985
rect 28445 43945 28457 43979
rect 28491 43976 28503 43979
rect 32582 43976 32588 43988
rect 28491 43948 32588 43976
rect 28491 43945 28503 43948
rect 28445 43939 28503 43945
rect 32582 43936 32588 43948
rect 32640 43936 32646 43988
rect 9030 43868 9036 43920
rect 9088 43908 9094 43920
rect 12345 43911 12403 43917
rect 12345 43908 12357 43911
rect 9088 43880 12357 43908
rect 9088 43868 9094 43880
rect 12345 43877 12357 43880
rect 12391 43877 12403 43911
rect 12345 43871 12403 43877
rect 19610 43868 19616 43920
rect 19668 43908 19674 43920
rect 22925 43911 22983 43917
rect 22925 43908 22937 43911
rect 19668 43880 22937 43908
rect 19668 43868 19674 43880
rect 22925 43877 22937 43880
rect 22971 43877 22983 43911
rect 22925 43871 22983 43877
rect 20364 43812 22876 43840
rect 20364 43781 20392 43812
rect 19797 43775 19855 43781
rect 19797 43741 19809 43775
rect 19843 43772 19855 43775
rect 20349 43775 20407 43781
rect 20349 43772 20361 43775
rect 19843 43744 20361 43772
rect 19843 43741 19855 43744
rect 19797 43735 19855 43741
rect 20349 43741 20361 43744
rect 20395 43741 20407 43775
rect 20349 43735 20407 43741
rect 22005 43775 22063 43781
rect 22005 43741 22017 43775
rect 22051 43772 22063 43775
rect 22278 43772 22284 43784
rect 22051 43744 22284 43772
rect 22051 43741 22063 43744
rect 22005 43735 22063 43741
rect 22278 43732 22284 43744
rect 22336 43732 22342 43784
rect 12158 43664 12164 43716
rect 12216 43664 12222 43716
rect 13446 43664 13452 43716
rect 13504 43664 13510 43716
rect 15565 43707 15623 43713
rect 15565 43673 15577 43707
rect 15611 43704 15623 43707
rect 16114 43704 16120 43716
rect 15611 43676 16120 43704
rect 15611 43673 15623 43676
rect 15565 43667 15623 43673
rect 16114 43664 16120 43676
rect 16172 43664 16178 43716
rect 16853 43707 16911 43713
rect 16853 43673 16865 43707
rect 16899 43704 16911 43707
rect 17034 43704 17040 43716
rect 16899 43676 17040 43704
rect 16899 43673 16911 43676
rect 16853 43667 16911 43673
rect 17034 43664 17040 43676
rect 17092 43664 17098 43716
rect 21174 43664 21180 43716
rect 21232 43664 21238 43716
rect 22738 43664 22744 43716
rect 22796 43664 22802 43716
rect 22848 43704 22876 43812
rect 28442 43800 28448 43852
rect 28500 43840 28506 43852
rect 28997 43843 29055 43849
rect 28997 43840 29009 43843
rect 28500 43812 29009 43840
rect 28500 43800 28506 43812
rect 28997 43809 29009 43812
rect 29043 43809 29055 43843
rect 28997 43803 29055 43809
rect 30285 43843 30343 43849
rect 30285 43809 30297 43843
rect 30331 43840 30343 43843
rect 32858 43840 32864 43852
rect 30331 43812 32864 43840
rect 30331 43809 30343 43812
rect 30285 43803 30343 43809
rect 32858 43800 32864 43812
rect 32916 43840 32922 43852
rect 33965 43843 34023 43849
rect 33965 43840 33977 43843
rect 32916 43812 33977 43840
rect 32916 43800 32922 43812
rect 33965 43809 33977 43812
rect 34011 43809 34023 43843
rect 33965 43803 34023 43809
rect 37734 43800 37740 43852
rect 37792 43800 37798 43852
rect 37921 43843 37979 43849
rect 37921 43809 37933 43843
rect 37967 43840 37979 43843
rect 38286 43840 38292 43852
rect 37967 43812 38292 43840
rect 37967 43809 37979 43812
rect 37921 43803 37979 43809
rect 38286 43800 38292 43812
rect 38344 43800 38350 43852
rect 48777 43843 48835 43849
rect 48777 43840 48789 43843
rect 45526 43812 48789 43840
rect 26234 43732 26240 43784
rect 26292 43772 26298 43784
rect 26292 43744 27568 43772
rect 26292 43732 26298 43744
rect 27540 43704 27568 43744
rect 28718 43732 28724 43784
rect 28776 43772 28782 43784
rect 30009 43775 30067 43781
rect 30009 43772 30021 43775
rect 28776 43744 30021 43772
rect 28776 43732 28782 43744
rect 30009 43741 30021 43744
rect 30055 43741 30067 43775
rect 30009 43735 30067 43741
rect 32214 43732 32220 43784
rect 32272 43732 32278 43784
rect 40770 43732 40776 43784
rect 40828 43772 40834 43784
rect 45526 43772 45554 43812
rect 48777 43809 48789 43812
rect 48823 43809 48835 43843
rect 48777 43803 48835 43809
rect 40828 43744 45554 43772
rect 40828 43732 40834 43744
rect 48498 43732 48504 43784
rect 48556 43732 48562 43784
rect 28813 43707 28871 43713
rect 28813 43704 28825 43707
rect 22848 43676 26234 43704
rect 27540 43676 28825 43704
rect 26206 43636 26234 43676
rect 28813 43673 28825 43676
rect 28859 43673 28871 43707
rect 28813 43667 28871 43673
rect 31294 43664 31300 43716
rect 31352 43664 31358 43716
rect 32493 43707 32551 43713
rect 32493 43673 32505 43707
rect 32539 43673 32551 43707
rect 32493 43667 32551 43673
rect 27614 43636 27620 43648
rect 26206 43608 27620 43636
rect 27614 43596 27620 43608
rect 27672 43596 27678 43648
rect 28902 43596 28908 43648
rect 28960 43596 28966 43648
rect 31754 43596 31760 43648
rect 31812 43596 31818 43648
rect 32508 43636 32536 43667
rect 33226 43664 33232 43716
rect 33284 43664 33290 43716
rect 37182 43664 37188 43716
rect 37240 43704 37246 43716
rect 37645 43707 37703 43713
rect 37645 43704 37657 43707
rect 37240 43676 37657 43704
rect 37240 43664 37246 43676
rect 37645 43673 37657 43676
rect 37691 43673 37703 43707
rect 37645 43667 37703 43673
rect 33318 43636 33324 43648
rect 32508 43608 33324 43636
rect 33318 43596 33324 43608
rect 33376 43596 33382 43648
rect 37274 43596 37280 43648
rect 37332 43596 37338 43648
rect 1104 43546 49864 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 27950 43546
rect 28002 43494 28014 43546
rect 28066 43494 28078 43546
rect 28130 43494 28142 43546
rect 28194 43494 28206 43546
rect 28258 43494 37950 43546
rect 38002 43494 38014 43546
rect 38066 43494 38078 43546
rect 38130 43494 38142 43546
rect 38194 43494 38206 43546
rect 38258 43494 47950 43546
rect 48002 43494 48014 43546
rect 48066 43494 48078 43546
rect 48130 43494 48142 43546
rect 48194 43494 48206 43546
rect 48258 43494 49864 43546
rect 1104 43472 49864 43494
rect 16850 43392 16856 43444
rect 16908 43392 16914 43444
rect 19150 43392 19156 43444
rect 19208 43392 19214 43444
rect 20346 43392 20352 43444
rect 20404 43392 20410 43444
rect 20898 43392 20904 43444
rect 20956 43392 20962 43444
rect 25866 43392 25872 43444
rect 25924 43392 25930 43444
rect 32324 43404 34560 43432
rect 12158 43324 12164 43376
rect 12216 43364 12222 43376
rect 21910 43364 21916 43376
rect 12216 43336 21916 43364
rect 12216 43324 12222 43336
rect 21910 43324 21916 43336
rect 21968 43324 21974 43376
rect 29178 43364 29184 43376
rect 28276 43336 29184 43364
rect 12066 43256 12072 43308
rect 12124 43256 12130 43308
rect 17037 43299 17095 43305
rect 17037 43265 17049 43299
rect 17083 43265 17095 43299
rect 17037 43259 17095 43265
rect 8938 43188 8944 43240
rect 8996 43228 9002 43240
rect 12253 43231 12311 43237
rect 12253 43228 12265 43231
rect 8996 43200 12265 43228
rect 8996 43188 9002 43200
rect 12253 43197 12265 43200
rect 12299 43197 12311 43231
rect 17052 43228 17080 43259
rect 19058 43256 19064 43308
rect 19116 43256 19122 43308
rect 20254 43256 20260 43308
rect 20312 43256 20318 43308
rect 21085 43299 21143 43305
rect 21085 43265 21097 43299
rect 21131 43265 21143 43299
rect 21085 43259 21143 43265
rect 19426 43228 19432 43240
rect 17052 43200 19432 43228
rect 12253 43191 12311 43197
rect 19426 43188 19432 43200
rect 19484 43188 19490 43240
rect 21100 43160 21128 43259
rect 25958 43256 25964 43308
rect 26016 43296 26022 43308
rect 26237 43299 26295 43305
rect 26237 43296 26249 43299
rect 26016 43268 26249 43296
rect 26016 43256 26022 43268
rect 26237 43265 26249 43268
rect 26283 43265 26295 43299
rect 26237 43259 26295 43265
rect 26326 43188 26332 43240
rect 26384 43188 26390 43240
rect 26513 43231 26571 43237
rect 26513 43197 26525 43231
rect 26559 43228 26571 43231
rect 27338 43228 27344 43240
rect 26559 43200 27344 43228
rect 26559 43197 26571 43200
rect 26513 43191 26571 43197
rect 27338 43188 27344 43200
rect 27396 43188 27402 43240
rect 28276 43160 28304 43336
rect 29178 43324 29184 43336
rect 29236 43324 29242 43376
rect 30374 43364 30380 43376
rect 30314 43336 30380 43364
rect 30374 43324 30380 43336
rect 30432 43364 30438 43376
rect 31294 43364 31300 43376
rect 30432 43336 31300 43364
rect 30432 43324 30438 43336
rect 31294 43324 31300 43336
rect 31352 43324 31358 43376
rect 32214 43256 32220 43308
rect 32272 43296 32278 43308
rect 32324 43305 32352 43404
rect 33226 43324 33232 43376
rect 33284 43324 33290 43376
rect 34532 43308 34560 43404
rect 40310 43392 40316 43444
rect 40368 43392 40374 43444
rect 34790 43324 34796 43376
rect 34848 43324 34854 43376
rect 32309 43299 32367 43305
rect 32309 43296 32321 43299
rect 32272 43268 32321 43296
rect 32272 43256 32278 43268
rect 32309 43265 32321 43268
rect 32355 43265 32367 43299
rect 32309 43259 32367 43265
rect 34514 43256 34520 43308
rect 34572 43256 34578 43308
rect 28718 43188 28724 43240
rect 28776 43228 28782 43240
rect 28813 43231 28871 43237
rect 28813 43228 28825 43231
rect 28776 43200 28825 43228
rect 28776 43188 28782 43200
rect 28813 43197 28825 43200
rect 28859 43197 28871 43231
rect 28813 43191 28871 43197
rect 29089 43231 29147 43237
rect 29089 43197 29101 43231
rect 29135 43228 29147 43231
rect 31938 43228 31944 43240
rect 29135 43200 31944 43228
rect 29135 43197 29147 43200
rect 29089 43191 29147 43197
rect 31938 43188 31944 43200
rect 31996 43188 32002 43240
rect 33226 43188 33232 43240
rect 33284 43228 33290 43240
rect 35912 43228 35940 43282
rect 38930 43256 38936 43308
rect 38988 43296 38994 43308
rect 39758 43296 39764 43308
rect 38988 43268 39764 43296
rect 38988 43256 38994 43268
rect 39758 43256 39764 43268
rect 39816 43296 39822 43308
rect 40221 43299 40279 43305
rect 40221 43296 40233 43299
rect 39816 43268 40233 43296
rect 39816 43256 39822 43268
rect 40221 43265 40233 43268
rect 40267 43265 40279 43299
rect 48777 43299 48835 43305
rect 48777 43296 48789 43299
rect 40221 43259 40279 43265
rect 45526 43268 48789 43296
rect 33284 43200 35940 43228
rect 33284 43188 33290 43200
rect 34146 43160 34152 43172
rect 21100 43132 28304 43160
rect 33980 43132 34152 43160
rect 28442 43052 28448 43104
rect 28500 43092 28506 43104
rect 30561 43095 30619 43101
rect 30561 43092 30573 43095
rect 28500 43064 30573 43092
rect 28500 43052 28506 43064
rect 30561 43061 30573 43064
rect 30607 43061 30619 43095
rect 30561 43055 30619 43061
rect 32572 43095 32630 43101
rect 32572 43061 32584 43095
rect 32618 43092 32630 43095
rect 33980 43092 34008 43132
rect 34146 43120 34152 43132
rect 34204 43120 34210 43172
rect 35820 43160 35848 43200
rect 40494 43188 40500 43240
rect 40552 43188 40558 43240
rect 41598 43188 41604 43240
rect 41656 43228 41662 43240
rect 45526 43228 45554 43268
rect 48777 43265 48789 43268
rect 48823 43265 48835 43299
rect 48777 43259 48835 43265
rect 41656 43200 45554 43228
rect 41656 43188 41662 43200
rect 48498 43188 48504 43240
rect 48556 43188 48562 43240
rect 35894 43160 35900 43172
rect 35820 43132 35900 43160
rect 35894 43120 35900 43132
rect 35952 43120 35958 43172
rect 32618 43064 34008 43092
rect 32618 43061 32630 43064
rect 32572 43055 32630 43061
rect 34054 43052 34060 43104
rect 34112 43052 34118 43104
rect 34164 43092 34192 43120
rect 36265 43095 36323 43101
rect 36265 43092 36277 43095
rect 34164 43064 36277 43092
rect 36265 43061 36277 43064
rect 36311 43061 36323 43095
rect 36265 43055 36323 43061
rect 39853 43095 39911 43101
rect 39853 43061 39865 43095
rect 39899 43092 39911 43095
rect 41230 43092 41236 43104
rect 39899 43064 41236 43092
rect 39899 43061 39911 43064
rect 39853 43055 39911 43061
rect 41230 43052 41236 43064
rect 41288 43052 41294 43104
rect 1104 43002 49864 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 32950 43002
rect 33002 42950 33014 43002
rect 33066 42950 33078 43002
rect 33130 42950 33142 43002
rect 33194 42950 33206 43002
rect 33258 42950 42950 43002
rect 43002 42950 43014 43002
rect 43066 42950 43078 43002
rect 43130 42950 43142 43002
rect 43194 42950 43206 43002
rect 43258 42950 49864 43002
rect 1104 42928 49864 42950
rect 27338 42848 27344 42900
rect 27396 42848 27402 42900
rect 9122 42712 9128 42764
rect 9180 42752 9186 42764
rect 9401 42755 9459 42761
rect 9401 42752 9413 42755
rect 9180 42724 9413 42752
rect 9180 42712 9186 42724
rect 9401 42721 9413 42724
rect 9447 42721 9459 42755
rect 9401 42715 9459 42721
rect 14550 42712 14556 42764
rect 14608 42752 14614 42764
rect 17405 42755 17463 42761
rect 17405 42752 17417 42755
rect 14608 42724 17417 42752
rect 14608 42712 14614 42724
rect 17405 42721 17417 42724
rect 17451 42721 17463 42755
rect 17405 42715 17463 42721
rect 35897 42755 35955 42761
rect 35897 42721 35909 42755
rect 35943 42752 35955 42755
rect 36906 42752 36912 42764
rect 35943 42724 36912 42752
rect 35943 42721 35955 42724
rect 35897 42715 35955 42721
rect 36906 42712 36912 42724
rect 36964 42712 36970 42764
rect 40678 42712 40684 42764
rect 40736 42712 40742 42764
rect 24670 42644 24676 42696
rect 24728 42684 24734 42696
rect 25593 42687 25651 42693
rect 25593 42684 25605 42687
rect 24728 42656 25605 42684
rect 24728 42644 24734 42656
rect 25593 42653 25605 42656
rect 25639 42653 25651 42687
rect 25593 42647 25651 42653
rect 34514 42644 34520 42696
rect 34572 42684 34578 42696
rect 35621 42687 35679 42693
rect 35621 42684 35633 42687
rect 34572 42656 35633 42684
rect 34572 42644 34578 42656
rect 35621 42653 35633 42656
rect 35667 42653 35679 42687
rect 35621 42647 35679 42653
rect 36998 42644 37004 42696
rect 37056 42644 37062 42696
rect 40497 42687 40555 42693
rect 40497 42653 40509 42687
rect 40543 42684 40555 42687
rect 43438 42684 43444 42696
rect 40543 42656 43444 42684
rect 40543 42653 40555 42656
rect 40497 42647 40555 42653
rect 43438 42644 43444 42656
rect 43496 42644 43502 42696
rect 48498 42644 48504 42696
rect 48556 42644 48562 42696
rect 48777 42687 48835 42693
rect 48777 42653 48789 42687
rect 48823 42653 48835 42687
rect 48777 42647 48835 42653
rect 9214 42576 9220 42628
rect 9272 42576 9278 42628
rect 17221 42619 17279 42625
rect 17221 42585 17233 42619
rect 17267 42616 17279 42619
rect 17402 42616 17408 42628
rect 17267 42588 17408 42616
rect 17267 42585 17279 42588
rect 17221 42579 17279 42585
rect 17402 42576 17408 42588
rect 17460 42576 17466 42628
rect 25866 42576 25872 42628
rect 25924 42576 25930 42628
rect 26206 42588 26358 42616
rect 24854 42508 24860 42560
rect 24912 42548 24918 42560
rect 26206 42548 26234 42588
rect 24912 42520 26234 42548
rect 24912 42508 24918 42520
rect 37182 42508 37188 42560
rect 37240 42548 37246 42560
rect 37369 42551 37427 42557
rect 37369 42548 37381 42551
rect 37240 42520 37381 42548
rect 37240 42508 37246 42520
rect 37369 42517 37381 42520
rect 37415 42517 37427 42551
rect 37369 42511 37427 42517
rect 40034 42508 40040 42560
rect 40092 42508 40098 42560
rect 40402 42508 40408 42560
rect 40460 42508 40466 42560
rect 40586 42508 40592 42560
rect 40644 42548 40650 42560
rect 48792 42548 48820 42647
rect 40644 42520 48820 42548
rect 40644 42508 40650 42520
rect 1104 42458 49864 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 27950 42458
rect 28002 42406 28014 42458
rect 28066 42406 28078 42458
rect 28130 42406 28142 42458
rect 28194 42406 28206 42458
rect 28258 42406 37950 42458
rect 38002 42406 38014 42458
rect 38066 42406 38078 42458
rect 38130 42406 38142 42458
rect 38194 42406 38206 42458
rect 38258 42406 47950 42458
rect 48002 42406 48014 42458
rect 48066 42406 48078 42458
rect 48130 42406 48142 42458
rect 48194 42406 48206 42458
rect 48258 42406 49864 42458
rect 1104 42384 49864 42406
rect 6270 42304 6276 42356
rect 6328 42344 6334 42356
rect 7193 42347 7251 42353
rect 7193 42344 7205 42347
rect 6328 42316 7205 42344
rect 6328 42304 6334 42316
rect 7193 42313 7205 42316
rect 7239 42313 7251 42347
rect 7193 42307 7251 42313
rect 20714 42304 20720 42356
rect 20772 42304 20778 42356
rect 22094 42304 22100 42356
rect 22152 42304 22158 42356
rect 30190 42344 30196 42356
rect 29288 42316 30196 42344
rect 6362 42236 6368 42288
rect 6420 42276 6426 42288
rect 8021 42279 8079 42285
rect 8021 42276 8033 42279
rect 6420 42248 8033 42276
rect 6420 42236 6426 42248
rect 8021 42245 8033 42248
rect 8067 42245 8079 42279
rect 24670 42276 24676 42288
rect 8021 42239 8079 42245
rect 24136 42248 24676 42276
rect 7098 42168 7104 42220
rect 7156 42168 7162 42220
rect 7834 42168 7840 42220
rect 7892 42168 7898 42220
rect 20901 42211 20959 42217
rect 20901 42177 20913 42211
rect 20947 42208 20959 42211
rect 20990 42208 20996 42220
rect 20947 42180 20996 42208
rect 20947 42177 20959 42180
rect 20901 42171 20959 42177
rect 20990 42168 20996 42180
rect 21048 42168 21054 42220
rect 22281 42211 22339 42217
rect 22281 42177 22293 42211
rect 22327 42208 22339 42211
rect 22554 42208 22560 42220
rect 22327 42180 22560 42208
rect 22327 42177 22339 42180
rect 22281 42171 22339 42177
rect 22554 42168 22560 42180
rect 22612 42168 22618 42220
rect 24136 42217 24164 42248
rect 24670 42236 24676 42248
rect 24728 42236 24734 42288
rect 24854 42236 24860 42288
rect 24912 42236 24918 42288
rect 27338 42236 27344 42288
rect 27396 42276 27402 42288
rect 27985 42279 28043 42285
rect 27985 42276 27997 42279
rect 27396 42248 27997 42276
rect 27396 42236 27402 42248
rect 27985 42245 27997 42248
rect 28031 42245 28043 42279
rect 29288 42276 29316 42316
rect 30190 42304 30196 42316
rect 30248 42304 30254 42356
rect 31754 42344 31760 42356
rect 30300 42316 31760 42344
rect 29210 42248 29316 42276
rect 27985 42239 28043 42245
rect 29362 42236 29368 42288
rect 29420 42276 29426 42288
rect 30300 42285 30328 42316
rect 31754 42304 31760 42316
rect 31812 42344 31818 42356
rect 32766 42344 32772 42356
rect 31812 42316 32772 42344
rect 31812 42304 31818 42316
rect 32766 42304 32772 42316
rect 32824 42304 32830 42356
rect 34514 42304 34520 42356
rect 34572 42304 34578 42356
rect 38286 42304 38292 42356
rect 38344 42344 38350 42356
rect 40037 42347 40095 42353
rect 40037 42344 40049 42347
rect 38344 42316 40049 42344
rect 38344 42304 38350 42316
rect 40037 42313 40049 42316
rect 40083 42313 40095 42347
rect 40037 42307 40095 42313
rect 41693 42347 41751 42353
rect 41693 42313 41705 42347
rect 41739 42344 41751 42347
rect 45186 42344 45192 42356
rect 41739 42316 45192 42344
rect 41739 42313 41751 42316
rect 41693 42307 41751 42313
rect 45186 42304 45192 42316
rect 45244 42304 45250 42356
rect 30285 42279 30343 42285
rect 30285 42276 30297 42279
rect 29420 42248 30297 42276
rect 29420 42236 29426 42248
rect 30285 42245 30297 42248
rect 30331 42245 30343 42279
rect 30285 42239 30343 42245
rect 31294 42236 31300 42288
rect 31352 42236 31358 42288
rect 34532 42276 34560 42304
rect 35894 42276 35900 42288
rect 33888 42248 34560 42276
rect 35374 42248 35900 42276
rect 33888 42217 33916 42248
rect 35894 42236 35900 42248
rect 35952 42276 35958 42288
rect 36998 42276 37004 42288
rect 35952 42248 37004 42276
rect 35952 42236 35958 42248
rect 36998 42236 37004 42248
rect 37056 42236 37062 42288
rect 39574 42236 39580 42288
rect 39632 42236 39638 42288
rect 24121 42211 24179 42217
rect 24121 42177 24133 42211
rect 24167 42177 24179 42211
rect 24121 42171 24179 42177
rect 33873 42211 33931 42217
rect 33873 42177 33885 42211
rect 33919 42177 33931 42211
rect 33873 42171 33931 42177
rect 41046 42168 41052 42220
rect 41104 42208 41110 42220
rect 41322 42208 41328 42220
rect 41104 42180 41328 42208
rect 41104 42168 41110 42180
rect 41322 42168 41328 42180
rect 41380 42208 41386 42220
rect 41601 42211 41659 42217
rect 41601 42208 41613 42211
rect 41380 42180 41613 42208
rect 41380 42168 41386 42180
rect 41601 42177 41613 42180
rect 41647 42177 41659 42211
rect 41601 42171 41659 42177
rect 24394 42100 24400 42152
rect 24452 42100 24458 42152
rect 27246 42100 27252 42152
rect 27304 42140 27310 42152
rect 27709 42143 27767 42149
rect 27709 42140 27721 42143
rect 27304 42112 27721 42140
rect 27304 42100 27310 42112
rect 27709 42109 27721 42112
rect 27755 42140 27767 42143
rect 28718 42140 28724 42152
rect 27755 42112 28724 42140
rect 27755 42109 27767 42112
rect 27709 42103 27767 42109
rect 28718 42100 28724 42112
rect 28776 42140 28782 42152
rect 30009 42143 30067 42149
rect 28776 42112 29776 42140
rect 28776 42100 28782 42112
rect 29748 42084 29776 42112
rect 30009 42109 30021 42143
rect 30055 42109 30067 42143
rect 30009 42103 30067 42109
rect 34149 42143 34207 42149
rect 34149 42109 34161 42143
rect 34195 42140 34207 42143
rect 35526 42140 35532 42152
rect 34195 42112 35532 42140
rect 34195 42109 34207 42112
rect 34149 42103 34207 42109
rect 29730 42032 29736 42084
rect 29788 42072 29794 42084
rect 30024 42072 30052 42103
rect 35526 42100 35532 42112
rect 35584 42100 35590 42152
rect 37826 42100 37832 42152
rect 37884 42140 37890 42152
rect 38289 42143 38347 42149
rect 38289 42140 38301 42143
rect 37884 42112 38301 42140
rect 37884 42100 37890 42112
rect 38289 42109 38301 42112
rect 38335 42109 38347 42143
rect 38289 42103 38347 42109
rect 38565 42143 38623 42149
rect 38565 42109 38577 42143
rect 38611 42140 38623 42143
rect 39298 42140 39304 42152
rect 38611 42112 39304 42140
rect 38611 42109 38623 42112
rect 38565 42103 38623 42109
rect 39298 42100 39304 42112
rect 39356 42100 39362 42152
rect 41874 42100 41880 42152
rect 41932 42100 41938 42152
rect 48498 42100 48504 42152
rect 48556 42100 48562 42152
rect 48777 42143 48835 42149
rect 48777 42109 48789 42143
rect 48823 42109 48835 42143
rect 48777 42103 48835 42109
rect 29788 42044 30052 42072
rect 29788 42032 29794 42044
rect 39850 42032 39856 42084
rect 39908 42072 39914 42084
rect 48792 42072 48820 42103
rect 39908 42044 48820 42072
rect 39908 42032 39914 42044
rect 20530 41964 20536 42016
rect 20588 42004 20594 42016
rect 22370 42004 22376 42016
rect 20588 41976 22376 42004
rect 20588 41964 20594 41976
rect 22370 41964 22376 41976
rect 22428 42004 22434 42016
rect 24854 42004 24860 42016
rect 22428 41976 24860 42004
rect 22428 41964 22434 41976
rect 24854 41964 24860 41976
rect 24912 41964 24918 42016
rect 25866 41964 25872 42016
rect 25924 41964 25930 42016
rect 29454 41964 29460 42016
rect 29512 41964 29518 42016
rect 31757 42007 31815 42013
rect 31757 41973 31769 42007
rect 31803 42004 31815 42007
rect 31938 42004 31944 42016
rect 31803 41976 31944 42004
rect 31803 41973 31815 41976
rect 31757 41967 31815 41973
rect 31938 41964 31944 41976
rect 31996 41964 32002 42016
rect 34882 41964 34888 42016
rect 34940 42004 34946 42016
rect 35621 42007 35679 42013
rect 35621 42004 35633 42007
rect 34940 41976 35633 42004
rect 34940 41964 34946 41976
rect 35621 41973 35633 41976
rect 35667 41973 35679 42007
rect 35621 41967 35679 41973
rect 41233 42007 41291 42013
rect 41233 41973 41245 42007
rect 41279 42004 41291 42007
rect 42334 42004 42340 42016
rect 41279 41976 42340 42004
rect 41279 41973 41291 41976
rect 41233 41967 41291 41973
rect 42334 41964 42340 41976
rect 42392 41964 42398 42016
rect 1104 41914 49864 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 32950 41914
rect 33002 41862 33014 41914
rect 33066 41862 33078 41914
rect 33130 41862 33142 41914
rect 33194 41862 33206 41914
rect 33258 41862 42950 41914
rect 43002 41862 43014 41914
rect 43066 41862 43078 41914
rect 43130 41862 43142 41914
rect 43194 41862 43206 41914
rect 43258 41862 49864 41914
rect 1104 41840 49864 41862
rect 1578 41760 1584 41812
rect 1636 41800 1642 41812
rect 23658 41800 23664 41812
rect 1636 41772 23664 41800
rect 1636 41760 1642 41772
rect 23658 41760 23664 41772
rect 23716 41760 23722 41812
rect 26326 41760 26332 41812
rect 26384 41800 26390 41812
rect 26973 41803 27031 41809
rect 26973 41800 26985 41803
rect 26384 41772 26985 41800
rect 26384 41760 26390 41772
rect 26973 41769 26985 41772
rect 27019 41769 27031 41803
rect 32858 41800 32864 41812
rect 26973 41763 27031 41769
rect 29656 41772 32864 41800
rect 22922 41692 22928 41744
rect 22980 41732 22986 41744
rect 22980 41704 23796 41732
rect 22980 41692 22986 41704
rect 21637 41667 21695 41673
rect 21637 41633 21649 41667
rect 21683 41664 21695 41667
rect 22646 41664 22652 41676
rect 21683 41636 22652 41664
rect 21683 41633 21695 41636
rect 21637 41627 21695 41633
rect 22646 41624 22652 41636
rect 22704 41624 22710 41676
rect 23658 41624 23664 41676
rect 23716 41624 23722 41676
rect 23768 41664 23796 41704
rect 25866 41692 25872 41744
rect 25924 41732 25930 41744
rect 25924 41704 27568 41732
rect 25924 41692 25930 41704
rect 27540 41673 27568 41704
rect 27433 41667 27491 41673
rect 27433 41664 27445 41667
rect 23768 41636 27445 41664
rect 27433 41633 27445 41636
rect 27479 41633 27491 41667
rect 27433 41627 27491 41633
rect 27525 41667 27583 41673
rect 27525 41633 27537 41667
rect 27571 41633 27583 41667
rect 27525 41627 27583 41633
rect 23676 41596 23704 41624
rect 26418 41596 26424 41608
rect 23676 41568 26424 41596
rect 26418 41556 26424 41568
rect 26476 41556 26482 41608
rect 1670 41488 1676 41540
rect 1728 41488 1734 41540
rect 21177 41531 21235 41537
rect 21177 41497 21189 41531
rect 21223 41528 21235 41531
rect 21913 41531 21971 41537
rect 21913 41528 21925 41531
rect 21223 41500 21925 41528
rect 21223 41497 21235 41500
rect 21177 41491 21235 41497
rect 21913 41497 21925 41500
rect 21959 41497 21971 41531
rect 21913 41491 21971 41497
rect 1765 41463 1823 41469
rect 1765 41429 1777 41463
rect 1811 41460 1823 41463
rect 10594 41460 10600 41472
rect 1811 41432 10600 41460
rect 1811 41429 1823 41432
rect 1765 41423 1823 41429
rect 10594 41420 10600 41432
rect 10652 41420 10658 41472
rect 21928 41460 21956 41491
rect 22370 41488 22376 41540
rect 22428 41488 22434 41540
rect 29656 41528 29684 41772
rect 32858 41760 32864 41772
rect 32916 41760 32922 41812
rect 35526 41760 35532 41812
rect 35584 41800 35590 41812
rect 36633 41803 36691 41809
rect 36633 41800 36645 41803
rect 35584 41772 36645 41800
rect 35584 41760 35590 41772
rect 36633 41769 36645 41772
rect 36679 41769 36691 41803
rect 36633 41763 36691 41769
rect 36906 41760 36912 41812
rect 36964 41800 36970 41812
rect 38841 41803 38899 41809
rect 38841 41800 38853 41803
rect 36964 41772 38853 41800
rect 36964 41760 36970 41772
rect 38841 41769 38853 41772
rect 38887 41769 38899 41803
rect 38841 41763 38899 41769
rect 31662 41624 31668 41676
rect 31720 41664 31726 41676
rect 34146 41664 34152 41676
rect 31720 41636 34152 41664
rect 31720 41624 31726 41636
rect 34146 41624 34152 41636
rect 34204 41624 34210 41676
rect 34514 41624 34520 41676
rect 34572 41664 34578 41676
rect 34698 41664 34704 41676
rect 34572 41636 34704 41664
rect 34572 41624 34578 41636
rect 34698 41624 34704 41636
rect 34756 41664 34762 41676
rect 34885 41667 34943 41673
rect 34885 41664 34897 41667
rect 34756 41636 34897 41664
rect 34756 41624 34762 41636
rect 34885 41633 34897 41636
rect 34931 41664 34943 41667
rect 37093 41667 37151 41673
rect 37093 41664 37105 41667
rect 34931 41636 37105 41664
rect 34931 41633 34943 41636
rect 34885 41627 34943 41633
rect 37093 41633 37105 41636
rect 37139 41664 37151 41667
rect 37826 41664 37832 41676
rect 37139 41636 37832 41664
rect 37139 41633 37151 41636
rect 37093 41627 37151 41633
rect 37826 41624 37832 41636
rect 37884 41624 37890 41676
rect 29730 41556 29736 41608
rect 29788 41596 29794 41608
rect 31389 41599 31447 41605
rect 31389 41596 31401 41599
rect 29788 41568 31401 41596
rect 29788 41556 29794 41568
rect 31389 41565 31401 41568
rect 31435 41565 31447 41599
rect 31389 41559 31447 41565
rect 23768 41500 29684 41528
rect 23768 41460 23796 41500
rect 31202 41488 31208 41540
rect 31260 41528 31266 41540
rect 31662 41528 31668 41540
rect 31260 41500 31668 41528
rect 31260 41488 31266 41500
rect 31662 41488 31668 41500
rect 31720 41488 31726 41540
rect 32950 41528 32956 41540
rect 32890 41500 32956 41528
rect 32950 41488 32956 41500
rect 33008 41488 33014 41540
rect 34422 41528 34428 41540
rect 33060 41500 34428 41528
rect 21928 41432 23796 41460
rect 24670 41420 24676 41472
rect 24728 41460 24734 41472
rect 27246 41460 27252 41472
rect 24728 41432 27252 41460
rect 24728 41420 24734 41432
rect 27246 41420 27252 41432
rect 27304 41420 27310 41472
rect 27341 41463 27399 41469
rect 27341 41429 27353 41463
rect 27387 41460 27399 41463
rect 33060 41460 33088 41500
rect 34422 41488 34428 41500
rect 34480 41488 34486 41540
rect 35161 41531 35219 41537
rect 35161 41497 35173 41531
rect 35207 41497 35219 41531
rect 36386 41500 36584 41528
rect 35161 41491 35219 41497
rect 27387 41432 33088 41460
rect 33137 41463 33195 41469
rect 27387 41429 27399 41432
rect 27341 41423 27399 41429
rect 33137 41429 33149 41463
rect 33183 41460 33195 41463
rect 33318 41460 33324 41472
rect 33183 41432 33324 41460
rect 33183 41429 33195 41432
rect 33137 41423 33195 41429
rect 33318 41420 33324 41432
rect 33376 41460 33382 41472
rect 34238 41460 34244 41472
rect 33376 41432 34244 41460
rect 33376 41420 33382 41432
rect 34238 41420 34244 41432
rect 34296 41420 34302 41472
rect 35176 41460 35204 41491
rect 35802 41460 35808 41472
rect 35176 41432 35808 41460
rect 35802 41420 35808 41432
rect 35860 41420 35866 41472
rect 36556 41460 36584 41500
rect 36630 41488 36636 41540
rect 36688 41528 36694 41540
rect 37369 41531 37427 41537
rect 37369 41528 37381 41531
rect 36688 41500 37381 41528
rect 36688 41488 36694 41500
rect 37369 41497 37381 41500
rect 37415 41497 37427 41531
rect 39574 41528 39580 41540
rect 38594 41500 39580 41528
rect 37369 41491 37427 41497
rect 36998 41460 37004 41472
rect 36556 41432 37004 41460
rect 36998 41420 37004 41432
rect 37056 41460 37062 41472
rect 38672 41460 38700 41500
rect 39574 41488 39580 41500
rect 39632 41488 39638 41540
rect 37056 41432 38700 41460
rect 37056 41420 37062 41432
rect 1104 41370 49864 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 27950 41370
rect 28002 41318 28014 41370
rect 28066 41318 28078 41370
rect 28130 41318 28142 41370
rect 28194 41318 28206 41370
rect 28258 41318 37950 41370
rect 38002 41318 38014 41370
rect 38066 41318 38078 41370
rect 38130 41318 38142 41370
rect 38194 41318 38206 41370
rect 38258 41318 47950 41370
rect 48002 41318 48014 41370
rect 48066 41318 48078 41370
rect 48130 41318 48142 41370
rect 48194 41318 48206 41370
rect 48258 41318 49864 41370
rect 1104 41296 49864 41318
rect 5810 41216 5816 41268
rect 5868 41216 5874 41268
rect 9858 41216 9864 41268
rect 9916 41216 9922 41268
rect 10778 41216 10784 41268
rect 10836 41216 10842 41268
rect 22005 41259 22063 41265
rect 22005 41225 22017 41259
rect 22051 41256 22063 41259
rect 22922 41256 22928 41268
rect 22051 41228 22928 41256
rect 22051 41225 22063 41228
rect 22005 41219 22063 41225
rect 22922 41216 22928 41228
rect 22980 41216 22986 41268
rect 24854 41216 24860 41268
rect 24912 41216 24918 41268
rect 25424 41228 27752 41256
rect 1946 41148 1952 41200
rect 2004 41188 2010 41200
rect 21177 41191 21235 41197
rect 21177 41188 21189 41191
rect 2004 41160 21189 41188
rect 2004 41148 2010 41160
rect 21177 41157 21189 41160
rect 21223 41188 21235 41191
rect 22373 41191 22431 41197
rect 22373 41188 22385 41191
rect 21223 41160 22385 41188
rect 21223 41157 21235 41160
rect 21177 41151 21235 41157
rect 22373 41157 22385 41160
rect 22419 41188 22431 41191
rect 22462 41188 22468 41200
rect 22419 41160 22468 41188
rect 22419 41157 22431 41160
rect 22373 41151 22431 41157
rect 22462 41148 22468 41160
rect 22520 41148 22526 41200
rect 24872 41188 24900 41216
rect 25314 41188 25320 41200
rect 24872 41160 25320 41188
rect 25314 41148 25320 41160
rect 25372 41188 25378 41200
rect 25424 41188 25452 41228
rect 27724 41188 27752 41228
rect 27798 41216 27804 41268
rect 27856 41256 27862 41268
rect 29457 41259 29515 41265
rect 29457 41256 29469 41259
rect 27856 41228 29469 41256
rect 27856 41216 27862 41228
rect 29457 41225 29469 41228
rect 29503 41225 29515 41259
rect 34882 41256 34888 41268
rect 29457 41219 29515 41225
rect 33428 41228 34888 41256
rect 29825 41191 29883 41197
rect 25372 41160 25530 41188
rect 27724 41160 28014 41188
rect 25372 41148 25378 41160
rect 29825 41157 29837 41191
rect 29871 41188 29883 41191
rect 30742 41188 30748 41200
rect 29871 41160 30748 41188
rect 29871 41157 29883 41160
rect 29825 41151 29883 41157
rect 30742 41148 30748 41160
rect 30800 41148 30806 41200
rect 32858 41148 32864 41200
rect 32916 41188 32922 41200
rect 33428 41197 33456 41228
rect 34882 41216 34888 41228
rect 34940 41216 34946 41268
rect 33413 41191 33471 41197
rect 33413 41188 33425 41191
rect 32916 41160 33425 41188
rect 32916 41148 32922 41160
rect 33413 41157 33425 41160
rect 33459 41157 33471 41191
rect 33413 41151 33471 41157
rect 5721 41123 5779 41129
rect 5721 41089 5733 41123
rect 5767 41120 5779 41123
rect 5767 41092 6914 41120
rect 5767 41089 5779 41092
rect 5721 41083 5779 41089
rect 6886 41052 6914 41092
rect 9766 41080 9772 41132
rect 9824 41080 9830 41132
rect 10686 41080 10692 41132
rect 10744 41080 10750 41132
rect 22066 41092 22692 41120
rect 17678 41052 17684 41064
rect 6886 41024 17684 41052
rect 17678 41012 17684 41024
rect 17736 41012 17742 41064
rect 21818 41012 21824 41064
rect 21876 41052 21882 41064
rect 22066 41052 22094 41092
rect 21876 41024 22094 41052
rect 21876 41012 21882 41024
rect 22370 41012 22376 41064
rect 22428 41052 22434 41064
rect 22664 41061 22692 41092
rect 27246 41080 27252 41132
rect 27304 41080 27310 41132
rect 29917 41123 29975 41129
rect 29917 41089 29929 41123
rect 29963 41120 29975 41123
rect 30834 41120 30840 41132
rect 29963 41092 30840 41120
rect 29963 41089 29975 41092
rect 29917 41083 29975 41089
rect 30834 41080 30840 41092
rect 30892 41080 30898 41132
rect 36998 41120 37004 41132
rect 34546 41106 37004 41120
rect 34532 41092 37004 41106
rect 22465 41055 22523 41061
rect 22465 41052 22477 41055
rect 22428 41024 22477 41052
rect 22428 41012 22434 41024
rect 22465 41021 22477 41024
rect 22511 41021 22523 41055
rect 22465 41015 22523 41021
rect 22649 41055 22707 41061
rect 22649 41021 22661 41055
rect 22695 41052 22707 41055
rect 24302 41052 24308 41064
rect 22695 41024 24308 41052
rect 22695 41021 22707 41024
rect 22649 41015 22707 41021
rect 22480 40916 22508 41015
rect 24302 41012 24308 41024
rect 24360 41012 24366 41064
rect 24578 41012 24584 41064
rect 24636 41052 24642 41064
rect 24765 41055 24823 41061
rect 24765 41052 24777 41055
rect 24636 41024 24777 41052
rect 24636 41012 24642 41024
rect 24765 41021 24777 41024
rect 24811 41021 24823 41055
rect 24765 41015 24823 41021
rect 25038 41012 25044 41064
rect 25096 41012 25102 41064
rect 27525 41055 27583 41061
rect 27525 41052 27537 41055
rect 27264 41024 27537 41052
rect 27264 40996 27292 41024
rect 27525 41021 27537 41024
rect 27571 41021 27583 41055
rect 27525 41015 27583 41021
rect 30006 41012 30012 41064
rect 30064 41012 30070 41064
rect 32306 41012 32312 41064
rect 32364 41052 32370 41064
rect 33137 41055 33195 41061
rect 33137 41052 33149 41055
rect 32364 41024 33149 41052
rect 32364 41012 32370 41024
rect 33137 41021 33149 41024
rect 33183 41021 33195 41055
rect 33870 41052 33876 41064
rect 33137 41015 33195 41021
rect 33244 41024 33876 41052
rect 26513 40987 26571 40993
rect 26513 40953 26525 40987
rect 26559 40984 26571 40987
rect 27246 40984 27252 40996
rect 26559 40956 27252 40984
rect 26559 40953 26571 40956
rect 26513 40947 26571 40953
rect 27246 40944 27252 40956
rect 27304 40944 27310 40996
rect 31294 40944 31300 40996
rect 31352 40984 31358 40996
rect 33042 40984 33048 40996
rect 31352 40956 33048 40984
rect 31352 40944 31358 40956
rect 33042 40944 33048 40956
rect 33100 40984 33106 40996
rect 33244 40984 33272 41024
rect 33870 41012 33876 41024
rect 33928 41052 33934 41064
rect 34532 41052 34560 41092
rect 36998 41080 37004 41092
rect 37056 41080 37062 41132
rect 37826 41080 37832 41132
rect 37884 41120 37890 41132
rect 38197 41123 38255 41129
rect 38197 41120 38209 41123
rect 37884 41092 38209 41120
rect 37884 41080 37890 41092
rect 38197 41089 38209 41092
rect 38243 41089 38255 41123
rect 38197 41083 38255 41089
rect 39574 41080 39580 41132
rect 39632 41080 39638 41132
rect 33928 41024 34560 41052
rect 33928 41012 33934 41024
rect 38470 41012 38476 41064
rect 38528 41012 38534 41064
rect 48498 41012 48504 41064
rect 48556 41012 48562 41064
rect 48590 41012 48596 41064
rect 48648 41052 48654 41064
rect 48777 41055 48835 41061
rect 48777 41052 48789 41055
rect 48648 41024 48789 41052
rect 48648 41012 48654 41024
rect 48777 41021 48789 41024
rect 48823 41021 48835 41055
rect 48777 41015 48835 41021
rect 33100 40956 33272 40984
rect 33100 40944 33106 40956
rect 23293 40919 23351 40925
rect 23293 40916 23305 40919
rect 22480 40888 23305 40916
rect 23293 40885 23305 40888
rect 23339 40916 23351 40919
rect 23382 40916 23388 40928
rect 23339 40888 23388 40916
rect 23339 40885 23351 40888
rect 23293 40879 23351 40885
rect 23382 40876 23388 40888
rect 23440 40876 23446 40928
rect 26602 40876 26608 40928
rect 26660 40916 26666 40928
rect 28997 40919 29055 40925
rect 28997 40916 29009 40919
rect 26660 40888 29009 40916
rect 26660 40876 26666 40888
rect 28997 40885 29009 40888
rect 29043 40916 29055 40919
rect 30374 40916 30380 40928
rect 29043 40888 30380 40916
rect 29043 40885 29055 40888
rect 28997 40879 29055 40885
rect 30374 40876 30380 40888
rect 30432 40876 30438 40928
rect 32582 40876 32588 40928
rect 32640 40916 32646 40928
rect 32950 40916 32956 40928
rect 32640 40888 32956 40916
rect 32640 40876 32646 40888
rect 32950 40876 32956 40888
rect 33008 40876 33014 40928
rect 34790 40876 34796 40928
rect 34848 40916 34854 40928
rect 34885 40919 34943 40925
rect 34885 40916 34897 40919
rect 34848 40888 34897 40916
rect 34848 40876 34854 40888
rect 34885 40885 34897 40888
rect 34931 40916 34943 40919
rect 35710 40916 35716 40928
rect 34931 40888 35716 40916
rect 34931 40885 34943 40888
rect 34885 40879 34943 40885
rect 35710 40876 35716 40888
rect 35768 40876 35774 40928
rect 39942 40876 39948 40928
rect 40000 40876 40006 40928
rect 1104 40826 49864 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 32950 40826
rect 33002 40774 33014 40826
rect 33066 40774 33078 40826
rect 33130 40774 33142 40826
rect 33194 40774 33206 40826
rect 33258 40774 42950 40826
rect 43002 40774 43014 40826
rect 43066 40774 43078 40826
rect 43130 40774 43142 40826
rect 43194 40774 43206 40826
rect 43258 40774 49864 40826
rect 1104 40752 49864 40774
rect 22002 40672 22008 40724
rect 22060 40712 22066 40724
rect 25501 40715 25559 40721
rect 25501 40712 25513 40715
rect 22060 40684 25513 40712
rect 22060 40672 22066 40684
rect 25501 40681 25513 40684
rect 25547 40681 25559 40715
rect 25501 40675 25559 40681
rect 31018 40672 31024 40724
rect 31076 40712 31082 40724
rect 31076 40684 35848 40712
rect 31076 40672 31082 40684
rect 20622 40604 20628 40656
rect 20680 40644 20686 40656
rect 23201 40647 23259 40653
rect 23201 40644 23213 40647
rect 20680 40616 23213 40644
rect 20680 40604 20686 40616
rect 23201 40613 23213 40616
rect 23247 40613 23259 40647
rect 23201 40607 23259 40613
rect 34422 40604 34428 40656
rect 34480 40644 34486 40656
rect 35253 40647 35311 40653
rect 35253 40644 35265 40647
rect 34480 40616 35265 40644
rect 34480 40604 34486 40616
rect 35253 40613 35265 40616
rect 35299 40613 35311 40647
rect 35253 40607 35311 40613
rect 23845 40579 23903 40585
rect 23845 40545 23857 40579
rect 23891 40576 23903 40579
rect 25038 40576 25044 40588
rect 23891 40548 25044 40576
rect 23891 40545 23903 40548
rect 23845 40539 23903 40545
rect 25038 40536 25044 40548
rect 25096 40536 25102 40588
rect 26145 40579 26203 40585
rect 26145 40545 26157 40579
rect 26191 40576 26203 40579
rect 26602 40576 26608 40588
rect 26191 40548 26608 40576
rect 26191 40545 26203 40548
rect 26145 40539 26203 40545
rect 26602 40536 26608 40548
rect 26660 40536 26666 40588
rect 27341 40579 27399 40585
rect 27341 40545 27353 40579
rect 27387 40576 27399 40579
rect 27430 40576 27436 40588
rect 27387 40548 27436 40576
rect 27387 40545 27399 40548
rect 27341 40539 27399 40545
rect 27430 40536 27436 40548
rect 27488 40536 27494 40588
rect 27706 40536 27712 40588
rect 27764 40576 27770 40588
rect 28902 40576 28908 40588
rect 27764 40548 28908 40576
rect 27764 40536 27770 40548
rect 28902 40536 28908 40548
rect 28960 40536 28966 40588
rect 30006 40536 30012 40588
rect 30064 40576 30070 40588
rect 31481 40579 31539 40585
rect 31481 40576 31493 40579
rect 30064 40548 31493 40576
rect 30064 40536 30070 40548
rect 31481 40545 31493 40548
rect 31527 40545 31539 40579
rect 31481 40539 31539 40545
rect 32674 40536 32680 40588
rect 32732 40536 32738 40588
rect 32766 40536 32772 40588
rect 32824 40536 32830 40588
rect 33502 40536 33508 40588
rect 33560 40576 33566 40588
rect 34057 40579 34115 40585
rect 34057 40576 34069 40579
rect 33560 40548 34069 40576
rect 33560 40536 33566 40548
rect 34057 40545 34069 40548
rect 34103 40545 34115 40579
rect 34057 40539 34115 40545
rect 34146 40536 34152 40588
rect 34204 40536 34210 40588
rect 35820 40585 35848 40684
rect 35805 40579 35863 40585
rect 35805 40545 35817 40579
rect 35851 40545 35863 40579
rect 35805 40539 35863 40545
rect 38746 40536 38752 40588
rect 38804 40576 38810 40588
rect 39209 40579 39267 40585
rect 39209 40576 39221 40579
rect 38804 40548 39221 40576
rect 38804 40536 38810 40548
rect 39209 40545 39221 40548
rect 39255 40545 39267 40579
rect 39209 40539 39267 40545
rect 39393 40579 39451 40585
rect 39393 40545 39405 40579
rect 39439 40576 39451 40579
rect 39942 40576 39948 40588
rect 39439 40548 39948 40576
rect 39439 40545 39451 40548
rect 39393 40539 39451 40545
rect 23661 40511 23719 40517
rect 23661 40477 23673 40511
rect 23707 40508 23719 40511
rect 26970 40508 26976 40520
rect 23707 40480 26976 40508
rect 23707 40477 23719 40480
rect 23661 40471 23719 40477
rect 26970 40468 26976 40480
rect 27028 40468 27034 40520
rect 27062 40468 27068 40520
rect 27120 40468 27126 40520
rect 27157 40511 27215 40517
rect 27157 40477 27169 40511
rect 27203 40508 27215 40511
rect 27522 40508 27528 40520
rect 27203 40480 27528 40508
rect 27203 40477 27215 40480
rect 27157 40471 27215 40477
rect 27522 40468 27528 40480
rect 27580 40468 27586 40520
rect 29730 40468 29736 40520
rect 29788 40468 29794 40520
rect 32585 40511 32643 40517
rect 32585 40477 32597 40511
rect 32631 40508 32643 40511
rect 32631 40480 38792 40508
rect 32631 40477 32643 40480
rect 32585 40471 32643 40477
rect 23474 40400 23480 40452
rect 23532 40440 23538 40452
rect 25869 40443 25927 40449
rect 25869 40440 25881 40443
rect 23532 40412 25881 40440
rect 23532 40400 23538 40412
rect 25869 40409 25881 40412
rect 25915 40409 25927 40443
rect 25869 40403 25927 40409
rect 25961 40443 26019 40449
rect 25961 40409 25973 40443
rect 26007 40440 26019 40443
rect 28902 40440 28908 40452
rect 26007 40412 28908 40440
rect 26007 40409 26019 40412
rect 25961 40403 26019 40409
rect 28902 40400 28908 40412
rect 28960 40400 28966 40452
rect 30009 40443 30067 40449
rect 30009 40409 30021 40443
rect 30055 40409 30067 40443
rect 30009 40403 30067 40409
rect 22186 40332 22192 40384
rect 22244 40372 22250 40384
rect 23569 40375 23627 40381
rect 23569 40372 23581 40375
rect 22244 40344 23581 40372
rect 22244 40332 22250 40344
rect 23569 40341 23581 40344
rect 23615 40341 23627 40375
rect 23569 40335 23627 40341
rect 26697 40375 26755 40381
rect 26697 40341 26709 40375
rect 26743 40372 26755 40375
rect 26878 40372 26884 40384
rect 26743 40344 26884 40372
rect 26743 40341 26755 40344
rect 26697 40335 26755 40341
rect 26878 40332 26884 40344
rect 26936 40332 26942 40384
rect 30024 40372 30052 40403
rect 30466 40400 30472 40452
rect 30524 40400 30530 40452
rect 34146 40440 34152 40452
rect 32232 40412 34152 40440
rect 31478 40372 31484 40384
rect 30024 40344 31484 40372
rect 31478 40332 31484 40344
rect 31536 40332 31542 40384
rect 32232 40381 32260 40412
rect 34146 40400 34152 40412
rect 34204 40400 34210 40452
rect 35621 40443 35679 40449
rect 35621 40409 35633 40443
rect 35667 40440 35679 40443
rect 37642 40440 37648 40452
rect 35667 40412 37648 40440
rect 35667 40409 35679 40412
rect 35621 40403 35679 40409
rect 37642 40400 37648 40412
rect 37700 40400 37706 40452
rect 38764 40440 38792 40480
rect 38838 40468 38844 40520
rect 38896 40508 38902 40520
rect 39408 40508 39436 40539
rect 39942 40536 39948 40548
rect 40000 40536 40006 40588
rect 48406 40536 48412 40588
rect 48464 40576 48470 40588
rect 48777 40579 48835 40585
rect 48777 40576 48789 40579
rect 48464 40548 48789 40576
rect 48464 40536 48470 40548
rect 48777 40545 48789 40548
rect 48823 40545 48835 40579
rect 48777 40539 48835 40545
rect 38896 40480 39436 40508
rect 38896 40468 38902 40480
rect 48498 40468 48504 40520
rect 48556 40468 48562 40520
rect 39206 40440 39212 40452
rect 38764 40412 39212 40440
rect 39206 40400 39212 40412
rect 39264 40400 39270 40452
rect 32217 40375 32275 40381
rect 32217 40341 32229 40375
rect 32263 40341 32275 40375
rect 32217 40335 32275 40341
rect 33594 40332 33600 40384
rect 33652 40332 33658 40384
rect 33686 40332 33692 40384
rect 33744 40372 33750 40384
rect 33965 40375 34023 40381
rect 33965 40372 33977 40375
rect 33744 40344 33977 40372
rect 33744 40332 33750 40344
rect 33965 40341 33977 40344
rect 34011 40341 34023 40375
rect 33965 40335 34023 40341
rect 35713 40375 35771 40381
rect 35713 40341 35725 40375
rect 35759 40372 35771 40375
rect 37366 40372 37372 40384
rect 35759 40344 37372 40372
rect 35759 40341 35771 40344
rect 35713 40335 35771 40341
rect 37366 40332 37372 40344
rect 37424 40372 37430 40384
rect 38378 40372 38384 40384
rect 37424 40344 38384 40372
rect 37424 40332 37430 40344
rect 38378 40332 38384 40344
rect 38436 40332 38442 40384
rect 38746 40332 38752 40384
rect 38804 40332 38810 40384
rect 39114 40332 39120 40384
rect 39172 40332 39178 40384
rect 1104 40282 49864 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 27950 40282
rect 28002 40230 28014 40282
rect 28066 40230 28078 40282
rect 28130 40230 28142 40282
rect 28194 40230 28206 40282
rect 28258 40230 37950 40282
rect 38002 40230 38014 40282
rect 38066 40230 38078 40282
rect 38130 40230 38142 40282
rect 38194 40230 38206 40282
rect 38258 40230 47950 40282
rect 48002 40230 48014 40282
rect 48066 40230 48078 40282
rect 48130 40230 48142 40282
rect 48194 40230 48206 40282
rect 48258 40230 49864 40282
rect 1104 40208 49864 40230
rect 24949 40171 25007 40177
rect 24949 40137 24961 40171
rect 24995 40168 25007 40171
rect 25038 40168 25044 40180
rect 24995 40140 25044 40168
rect 24995 40137 25007 40140
rect 24949 40131 25007 40137
rect 25038 40128 25044 40140
rect 25096 40128 25102 40180
rect 30466 40168 30472 40180
rect 28828 40140 30472 40168
rect 25314 40100 25320 40112
rect 24702 40072 25320 40100
rect 25314 40060 25320 40072
rect 25372 40100 25378 40112
rect 28828 40100 28856 40140
rect 30466 40128 30472 40140
rect 30524 40168 30530 40180
rect 31294 40168 31300 40180
rect 30524 40140 31300 40168
rect 30524 40128 30530 40140
rect 31294 40128 31300 40140
rect 31352 40128 31358 40180
rect 34057 40171 34115 40177
rect 34057 40137 34069 40171
rect 34103 40168 34115 40171
rect 35066 40168 35072 40180
rect 34103 40140 35072 40168
rect 34103 40137 34115 40140
rect 34057 40131 34115 40137
rect 35066 40128 35072 40140
rect 35124 40128 35130 40180
rect 35894 40128 35900 40180
rect 35952 40168 35958 40180
rect 36449 40171 36507 40177
rect 36449 40168 36461 40171
rect 35952 40140 36461 40168
rect 35952 40128 35958 40140
rect 36449 40137 36461 40140
rect 36495 40168 36507 40171
rect 36814 40168 36820 40180
rect 36495 40140 36820 40168
rect 36495 40137 36507 40140
rect 36449 40131 36507 40137
rect 36814 40128 36820 40140
rect 36872 40128 36878 40180
rect 39482 40128 39488 40180
rect 39540 40168 39546 40180
rect 40313 40171 40371 40177
rect 40313 40168 40325 40171
rect 39540 40140 40325 40168
rect 39540 40128 39546 40140
rect 40313 40137 40325 40140
rect 40359 40137 40371 40171
rect 40313 40131 40371 40137
rect 40773 40171 40831 40177
rect 40773 40137 40785 40171
rect 40819 40168 40831 40171
rect 42702 40168 42708 40180
rect 40819 40140 42708 40168
rect 40819 40137 40831 40140
rect 40773 40131 40831 40137
rect 42702 40128 42708 40140
rect 42760 40128 42766 40180
rect 33870 40100 33876 40112
rect 25372 40072 28934 40100
rect 33810 40072 33876 40100
rect 25372 40060 25378 40072
rect 33870 40060 33876 40072
rect 33928 40100 33934 40112
rect 33928 40072 35466 40100
rect 33928 40060 33934 40072
rect 38838 40060 38844 40112
rect 38896 40060 38902 40112
rect 39574 40060 39580 40112
rect 39632 40060 39638 40112
rect 41138 40060 41144 40112
rect 41196 40060 41202 40112
rect 22646 39992 22652 40044
rect 22704 40032 22710 40044
rect 23201 40035 23259 40041
rect 23201 40032 23213 40035
rect 22704 40004 23213 40032
rect 22704 39992 22710 40004
rect 23201 40001 23213 40004
rect 23247 40001 23259 40035
rect 23201 39995 23259 40001
rect 34698 39992 34704 40044
rect 34756 39992 34762 40044
rect 37826 39992 37832 40044
rect 37884 40032 37890 40044
rect 38562 40032 38568 40044
rect 37884 40004 38568 40032
rect 37884 39992 37890 40004
rect 38562 39992 38568 40004
rect 38620 39992 38626 40044
rect 41230 39992 41236 40044
rect 41288 39992 41294 40044
rect 23477 39967 23535 39973
rect 23477 39933 23489 39967
rect 23523 39964 23535 39967
rect 23566 39964 23572 39976
rect 23523 39936 23572 39964
rect 23523 39933 23535 39936
rect 23477 39927 23535 39933
rect 23566 39924 23572 39936
rect 23624 39924 23630 39976
rect 28169 39967 28227 39973
rect 28169 39933 28181 39967
rect 28215 39933 28227 39967
rect 28169 39927 28227 39933
rect 23658 39788 23664 39840
rect 23716 39828 23722 39840
rect 27798 39828 27804 39840
rect 23716 39800 27804 39828
rect 23716 39788 23722 39800
rect 27798 39788 27804 39800
rect 27856 39788 27862 39840
rect 28184 39828 28212 39927
rect 28442 39924 28448 39976
rect 28500 39924 28506 39976
rect 32306 39924 32312 39976
rect 32364 39924 32370 39976
rect 32585 39967 32643 39973
rect 32585 39964 32597 39967
rect 32416 39936 32597 39964
rect 30374 39856 30380 39908
rect 30432 39896 30438 39908
rect 32416 39896 32444 39936
rect 32585 39933 32597 39936
rect 32631 39933 32643 39967
rect 32585 39927 32643 39933
rect 33778 39924 33784 39976
rect 33836 39964 33842 39976
rect 34977 39967 35035 39973
rect 34977 39964 34989 39967
rect 33836 39936 34989 39964
rect 33836 39924 33842 39936
rect 34977 39933 34989 39936
rect 35023 39933 35035 39967
rect 34977 39927 35035 39933
rect 35618 39924 35624 39976
rect 35676 39964 35682 39976
rect 40126 39964 40132 39976
rect 35676 39936 40132 39964
rect 35676 39924 35682 39936
rect 40126 39924 40132 39936
rect 40184 39924 40190 39976
rect 41417 39967 41475 39973
rect 41417 39933 41429 39967
rect 41463 39964 41475 39967
rect 41782 39964 41788 39976
rect 41463 39936 41788 39964
rect 41463 39933 41475 39936
rect 41417 39927 41475 39933
rect 41782 39924 41788 39936
rect 41840 39924 41846 39976
rect 48498 39924 48504 39976
rect 48556 39924 48562 39976
rect 48777 39967 48835 39973
rect 48777 39933 48789 39967
rect 48823 39933 48835 39967
rect 48777 39927 48835 39933
rect 41598 39896 41604 39908
rect 30432 39868 32444 39896
rect 39868 39868 41604 39896
rect 30432 39856 30438 39868
rect 29730 39828 29736 39840
rect 28184 39800 29736 39828
rect 29730 39788 29736 39800
rect 29788 39788 29794 39840
rect 29822 39788 29828 39840
rect 29880 39828 29886 39840
rect 29917 39831 29975 39837
rect 29917 39828 29929 39831
rect 29880 39800 29929 39828
rect 29880 39788 29886 39800
rect 29917 39797 29929 39800
rect 29963 39797 29975 39831
rect 29917 39791 29975 39797
rect 30098 39788 30104 39840
rect 30156 39828 30162 39840
rect 34054 39828 34060 39840
rect 30156 39800 34060 39828
rect 30156 39788 30162 39800
rect 34054 39788 34060 39800
rect 34112 39788 34118 39840
rect 34330 39788 34336 39840
rect 34388 39828 34394 39840
rect 39868 39828 39896 39868
rect 41598 39856 41604 39868
rect 41656 39856 41662 39908
rect 34388 39800 39896 39828
rect 34388 39788 34394 39800
rect 39942 39788 39948 39840
rect 40000 39828 40006 39840
rect 48792 39828 48820 39927
rect 40000 39800 48820 39828
rect 40000 39788 40006 39800
rect 1104 39738 49864 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 32950 39738
rect 33002 39686 33014 39738
rect 33066 39686 33078 39738
rect 33130 39686 33142 39738
rect 33194 39686 33206 39738
rect 33258 39686 42950 39738
rect 43002 39686 43014 39738
rect 43066 39686 43078 39738
rect 43130 39686 43142 39738
rect 43194 39686 43206 39738
rect 43258 39686 49864 39738
rect 1104 39664 49864 39686
rect 28718 39624 28724 39636
rect 24504 39596 28724 39624
rect 22005 39559 22063 39565
rect 22005 39525 22017 39559
rect 22051 39556 22063 39559
rect 24394 39556 24400 39568
rect 22051 39528 24400 39556
rect 22051 39525 22063 39528
rect 22005 39519 22063 39525
rect 24394 39516 24400 39528
rect 24452 39516 24458 39568
rect 22278 39448 22284 39500
rect 22336 39488 22342 39500
rect 22557 39491 22615 39497
rect 22557 39488 22569 39491
rect 22336 39460 22569 39488
rect 22336 39448 22342 39460
rect 22557 39457 22569 39460
rect 22603 39457 22615 39491
rect 22557 39451 22615 39457
rect 22373 39423 22431 39429
rect 22373 39389 22385 39423
rect 22419 39420 22431 39423
rect 22462 39420 22468 39432
rect 22419 39392 22468 39420
rect 22419 39389 22431 39392
rect 22373 39383 22431 39389
rect 22462 39380 22468 39392
rect 22520 39420 22526 39432
rect 24504 39420 24532 39596
rect 28718 39584 28724 39596
rect 28776 39584 28782 39636
rect 30834 39584 30840 39636
rect 30892 39624 30898 39636
rect 32677 39627 32735 39633
rect 32677 39624 32689 39627
rect 30892 39596 32689 39624
rect 30892 39584 30898 39596
rect 32677 39593 32689 39596
rect 32723 39593 32735 39627
rect 38654 39624 38660 39636
rect 32677 39587 32735 39593
rect 36004 39596 38660 39624
rect 31478 39516 31484 39568
rect 31536 39556 31542 39568
rect 31941 39559 31999 39565
rect 31941 39556 31953 39559
rect 31536 39528 31953 39556
rect 31536 39516 31542 39528
rect 31941 39525 31953 39528
rect 31987 39556 31999 39559
rect 31987 39528 32720 39556
rect 31987 39525 31999 39528
rect 31941 39519 31999 39525
rect 24578 39448 24584 39500
rect 24636 39448 24642 39500
rect 24857 39491 24915 39497
rect 24857 39457 24869 39491
rect 24903 39488 24915 39491
rect 24946 39488 24952 39500
rect 24903 39460 24952 39488
rect 24903 39457 24915 39460
rect 24857 39451 24915 39457
rect 24946 39448 24952 39460
rect 25004 39488 25010 39500
rect 28350 39488 28356 39500
rect 25004 39460 28356 39488
rect 25004 39448 25010 39460
rect 28350 39448 28356 39460
rect 28408 39448 28414 39500
rect 30193 39491 30251 39497
rect 30193 39457 30205 39491
rect 30239 39488 30251 39491
rect 32582 39488 32588 39500
rect 30239 39460 32588 39488
rect 30239 39457 30251 39460
rect 30193 39451 30251 39457
rect 32582 39448 32588 39460
rect 32640 39448 32646 39500
rect 32692 39488 32720 39528
rect 34054 39516 34060 39568
rect 34112 39556 34118 39568
rect 35894 39556 35900 39568
rect 34112 39528 35900 39556
rect 34112 39516 34118 39528
rect 35894 39516 35900 39528
rect 35952 39516 35958 39568
rect 33229 39491 33287 39497
rect 33229 39488 33241 39491
rect 32692 39460 33241 39488
rect 33229 39457 33241 39460
rect 33275 39457 33287 39491
rect 33229 39451 33287 39457
rect 33502 39448 33508 39500
rect 33560 39488 33566 39500
rect 34241 39491 34299 39497
rect 34241 39488 34253 39491
rect 33560 39460 34253 39488
rect 33560 39448 33566 39460
rect 34241 39457 34253 39460
rect 34287 39488 34299 39491
rect 36004 39488 36032 39596
rect 38654 39584 38660 39596
rect 38712 39584 38718 39636
rect 38749 39627 38807 39633
rect 38749 39593 38761 39627
rect 38795 39624 38807 39627
rect 43806 39624 43812 39636
rect 38795 39596 43812 39624
rect 38795 39593 38807 39596
rect 38749 39587 38807 39593
rect 43806 39584 43812 39596
rect 43864 39584 43870 39636
rect 43898 39584 43904 39636
rect 43956 39624 43962 39636
rect 48314 39624 48320 39636
rect 43956 39596 48320 39624
rect 43956 39584 43962 39596
rect 48314 39584 48320 39596
rect 48372 39584 48378 39636
rect 38378 39516 38384 39568
rect 38436 39556 38442 39568
rect 39942 39556 39948 39568
rect 38436 39528 39948 39556
rect 38436 39516 38442 39528
rect 39942 39516 39948 39528
rect 40000 39516 40006 39568
rect 34287 39460 36032 39488
rect 36265 39491 36323 39497
rect 34287 39457 34299 39460
rect 34241 39451 34299 39457
rect 36265 39457 36277 39491
rect 36311 39488 36323 39491
rect 37550 39488 37556 39500
rect 36311 39460 37556 39488
rect 36311 39457 36323 39460
rect 36265 39451 36323 39457
rect 37550 39448 37556 39460
rect 37608 39488 37614 39500
rect 38286 39488 38292 39500
rect 37608 39460 38292 39488
rect 37608 39448 37614 39460
rect 38286 39448 38292 39460
rect 38344 39448 38350 39500
rect 38746 39448 38752 39500
rect 38804 39488 38810 39500
rect 39209 39491 39267 39497
rect 39209 39488 39221 39491
rect 38804 39460 39221 39488
rect 38804 39448 38810 39460
rect 39209 39457 39221 39460
rect 39255 39457 39267 39491
rect 39209 39451 39267 39457
rect 39298 39448 39304 39500
rect 39356 39448 39362 39500
rect 41233 39491 41291 39497
rect 41233 39457 41245 39491
rect 41279 39488 41291 39491
rect 42794 39488 42800 39500
rect 41279 39460 42800 39488
rect 41279 39457 41291 39460
rect 41233 39451 41291 39457
rect 42794 39448 42800 39460
rect 42852 39448 42858 39500
rect 48774 39448 48780 39500
rect 48832 39448 48838 39500
rect 22520 39392 24532 39420
rect 22520 39380 22526 39392
rect 28442 39380 28448 39432
rect 28500 39420 28506 39432
rect 28810 39420 28816 39432
rect 28500 39392 28816 39420
rect 28500 39380 28506 39392
rect 28810 39380 28816 39392
rect 28868 39380 28874 39432
rect 33045 39423 33103 39429
rect 33045 39389 33057 39423
rect 33091 39420 33103 39423
rect 34514 39420 34520 39432
rect 33091 39392 34520 39420
rect 33091 39389 33103 39392
rect 33045 39383 33103 39389
rect 34514 39380 34520 39392
rect 34572 39380 34578 39432
rect 34698 39380 34704 39432
rect 34756 39420 34762 39432
rect 35989 39423 36047 39429
rect 35989 39420 36001 39423
rect 34756 39392 36001 39420
rect 34756 39380 34762 39392
rect 35989 39389 36001 39392
rect 36035 39389 36047 39423
rect 35989 39383 36047 39389
rect 40310 39380 40316 39432
rect 40368 39420 40374 39432
rect 40957 39423 41015 39429
rect 40957 39420 40969 39423
rect 40368 39392 40969 39420
rect 40368 39380 40374 39392
rect 40957 39389 40969 39392
rect 41003 39389 41015 39423
rect 40957 39383 41015 39389
rect 48498 39380 48504 39432
rect 48556 39380 48562 39432
rect 25130 39352 25136 39364
rect 21468 39324 25136 39352
rect 1854 39244 1860 39296
rect 1912 39284 1918 39296
rect 21468 39293 21496 39324
rect 22480 39293 22508 39324
rect 25130 39312 25136 39324
rect 25188 39312 25194 39364
rect 25314 39312 25320 39364
rect 25372 39312 25378 39364
rect 26142 39312 26148 39364
rect 26200 39352 26206 39364
rect 26200 39324 28764 39352
rect 26200 39312 26206 39324
rect 21453 39287 21511 39293
rect 21453 39284 21465 39287
rect 1912 39256 21465 39284
rect 1912 39244 1918 39256
rect 21453 39253 21465 39256
rect 21499 39253 21511 39287
rect 21453 39247 21511 39253
rect 22465 39287 22523 39293
rect 22465 39253 22477 39287
rect 22511 39253 22523 39287
rect 22465 39247 22523 39253
rect 23566 39244 23572 39296
rect 23624 39284 23630 39296
rect 26329 39287 26387 39293
rect 26329 39284 26341 39287
rect 23624 39256 26341 39284
rect 23624 39244 23630 39256
rect 26329 39253 26341 39256
rect 26375 39284 26387 39287
rect 28626 39284 28632 39296
rect 26375 39256 28632 39284
rect 26375 39253 26387 39256
rect 26329 39247 26387 39253
rect 28626 39244 28632 39256
rect 28684 39244 28690 39296
rect 28736 39284 28764 39324
rect 28994 39312 29000 39364
rect 29052 39352 29058 39364
rect 29454 39352 29460 39364
rect 29052 39324 29460 39352
rect 29052 39312 29058 39324
rect 29454 39312 29460 39324
rect 29512 39352 29518 39364
rect 30466 39352 30472 39364
rect 29512 39324 30472 39352
rect 29512 39312 29518 39324
rect 30466 39312 30472 39324
rect 30524 39312 30530 39364
rect 30558 39312 30564 39364
rect 30616 39352 30622 39364
rect 34057 39355 34115 39361
rect 34057 39352 34069 39355
rect 30616 39324 30958 39352
rect 32968 39324 34069 39352
rect 30616 39312 30622 39324
rect 31110 39284 31116 39296
rect 28736 39256 31116 39284
rect 31110 39244 31116 39256
rect 31168 39284 31174 39296
rect 32968 39284 32996 39324
rect 34057 39321 34069 39324
rect 34103 39352 34115 39355
rect 35345 39355 35403 39361
rect 35345 39352 35357 39355
rect 34103 39324 35357 39352
rect 34103 39321 34115 39324
rect 34057 39315 34115 39321
rect 35345 39321 35357 39324
rect 35391 39321 35403 39355
rect 35345 39315 35403 39321
rect 36998 39312 37004 39364
rect 37056 39312 37062 39364
rect 39390 39312 39396 39364
rect 39448 39352 39454 39364
rect 41230 39352 41236 39364
rect 39448 39324 41236 39352
rect 39448 39312 39454 39324
rect 41230 39312 41236 39324
rect 41288 39312 41294 39364
rect 43438 39352 43444 39364
rect 42458 39324 43444 39352
rect 43438 39312 43444 39324
rect 43496 39352 43502 39364
rect 46382 39352 46388 39364
rect 43496 39324 46388 39352
rect 43496 39312 43502 39324
rect 46382 39312 46388 39324
rect 46440 39312 46446 39364
rect 31168 39256 32996 39284
rect 33137 39287 33195 39293
rect 31168 39244 31174 39256
rect 33137 39253 33149 39287
rect 33183 39284 33195 39287
rect 33597 39287 33655 39293
rect 33597 39284 33609 39287
rect 33183 39256 33609 39284
rect 33183 39253 33195 39256
rect 33137 39247 33195 39253
rect 33597 39253 33609 39256
rect 33643 39253 33655 39287
rect 33597 39247 33655 39253
rect 33965 39287 34023 39293
rect 33965 39253 33977 39287
rect 34011 39284 34023 39287
rect 34974 39284 34980 39296
rect 34011 39256 34980 39284
rect 34011 39253 34023 39256
rect 33965 39247 34023 39253
rect 34974 39244 34980 39256
rect 35032 39244 35038 39296
rect 35250 39244 35256 39296
rect 35308 39284 35314 39296
rect 37734 39284 37740 39296
rect 35308 39256 37740 39284
rect 35308 39244 35314 39256
rect 37734 39244 37740 39256
rect 37792 39244 37798 39296
rect 38838 39244 38844 39296
rect 38896 39284 38902 39296
rect 39117 39287 39175 39293
rect 39117 39284 39129 39287
rect 38896 39256 39129 39284
rect 38896 39244 38902 39256
rect 39117 39253 39129 39256
rect 39163 39253 39175 39287
rect 39117 39247 39175 39253
rect 39942 39244 39948 39296
rect 40000 39284 40006 39296
rect 42705 39287 42763 39293
rect 42705 39284 42717 39287
rect 40000 39256 42717 39284
rect 40000 39244 40006 39256
rect 42705 39253 42717 39256
rect 42751 39253 42763 39287
rect 42705 39247 42763 39253
rect 1104 39194 49864 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 27950 39194
rect 28002 39142 28014 39194
rect 28066 39142 28078 39194
rect 28130 39142 28142 39194
rect 28194 39142 28206 39194
rect 28258 39142 37950 39194
rect 38002 39142 38014 39194
rect 38066 39142 38078 39194
rect 38130 39142 38142 39194
rect 38194 39142 38206 39194
rect 38258 39142 47950 39194
rect 48002 39142 48014 39194
rect 48066 39142 48078 39194
rect 48130 39142 48142 39194
rect 48194 39142 48206 39194
rect 48258 39142 49864 39194
rect 1104 39120 49864 39142
rect 22373 39083 22431 39089
rect 22373 39080 22385 39083
rect 22066 39052 22385 39080
rect 934 38904 940 38956
rect 992 38944 998 38956
rect 1765 38947 1823 38953
rect 1765 38944 1777 38947
rect 992 38916 1777 38944
rect 992 38904 998 38916
rect 1765 38913 1777 38916
rect 1811 38913 1823 38947
rect 1765 38907 1823 38913
rect 1854 38904 1860 38956
rect 1912 38944 1918 38956
rect 22066 38944 22094 39052
rect 22373 39049 22385 39052
rect 22419 39080 22431 39083
rect 23201 39083 23259 39089
rect 23201 39080 23213 39083
rect 22419 39052 23213 39080
rect 22419 39049 22431 39052
rect 22373 39043 22431 39049
rect 23201 39049 23213 39052
rect 23247 39080 23259 39083
rect 23658 39080 23664 39092
rect 23247 39052 23664 39080
rect 23247 39049 23259 39052
rect 23201 39043 23259 39049
rect 23658 39040 23664 39052
rect 23716 39040 23722 39092
rect 24486 39040 24492 39092
rect 24544 39040 24550 39092
rect 25869 39083 25927 39089
rect 25869 39049 25881 39083
rect 25915 39080 25927 39083
rect 25958 39080 25964 39092
rect 25915 39052 25964 39080
rect 25915 39049 25927 39052
rect 25869 39043 25927 39049
rect 25958 39040 25964 39052
rect 26016 39040 26022 39092
rect 26234 39080 26240 39092
rect 26206 39040 26240 39080
rect 26292 39040 26298 39092
rect 27154 39040 27160 39092
rect 27212 39080 27218 39092
rect 27341 39083 27399 39089
rect 27341 39080 27353 39083
rect 27212 39052 27353 39080
rect 27212 39040 27218 39052
rect 27341 39049 27353 39052
rect 27387 39049 27399 39083
rect 28905 39083 28963 39089
rect 27341 39043 27399 39049
rect 27724 39052 28580 39080
rect 23293 39015 23351 39021
rect 23293 38981 23305 39015
rect 23339 39012 23351 39015
rect 23382 39012 23388 39024
rect 23339 38984 23388 39012
rect 23339 38981 23351 38984
rect 23293 38975 23351 38981
rect 23382 38972 23388 38984
rect 23440 38972 23446 39024
rect 24949 39015 25007 39021
rect 24949 38981 24961 39015
rect 24995 39012 25007 39015
rect 26206 39012 26234 39040
rect 27724 39012 27752 39052
rect 24995 38984 26234 39012
rect 26344 38984 27752 39012
rect 27801 39015 27859 39021
rect 24995 38981 25007 38984
rect 24949 38975 25007 38981
rect 1912 38916 22094 38944
rect 1912 38904 1918 38916
rect 24854 38904 24860 38956
rect 24912 38904 24918 38956
rect 25130 38904 25136 38956
rect 25188 38944 25194 38956
rect 26142 38944 26148 38956
rect 25188 38916 26148 38944
rect 25188 38904 25194 38916
rect 26142 38904 26148 38916
rect 26200 38904 26206 38956
rect 26234 38904 26240 38956
rect 26292 38904 26298 38956
rect 26344 38953 26372 38984
rect 27801 38981 27813 39015
rect 27847 39012 27859 39015
rect 28442 39012 28448 39024
rect 27847 38984 28448 39012
rect 27847 38981 27859 38984
rect 27801 38975 27859 38981
rect 28442 38972 28448 38984
rect 28500 38972 28506 39024
rect 28552 39012 28580 39052
rect 28905 39049 28917 39083
rect 28951 39080 28963 39083
rect 30098 39080 30104 39092
rect 28951 39052 30104 39080
rect 28951 39049 28963 39052
rect 28905 39043 28963 39049
rect 30098 39040 30104 39052
rect 30156 39040 30162 39092
rect 30466 39040 30472 39092
rect 30524 39080 30530 39092
rect 33502 39080 33508 39092
rect 30524 39052 33508 39080
rect 30524 39040 30530 39052
rect 33502 39040 33508 39052
rect 33560 39040 33566 39092
rect 33594 39040 33600 39092
rect 33652 39080 33658 39092
rect 34149 39083 34207 39089
rect 34149 39080 34161 39083
rect 33652 39052 34161 39080
rect 33652 39040 33658 39052
rect 34149 39049 34161 39052
rect 34195 39049 34207 39083
rect 34149 39043 34207 39049
rect 34422 39040 34428 39092
rect 34480 39080 34486 39092
rect 35342 39080 35348 39092
rect 34480 39052 35348 39080
rect 34480 39040 34486 39052
rect 35342 39040 35348 39052
rect 35400 39040 35406 39092
rect 35529 39083 35587 39089
rect 35529 39080 35541 39083
rect 35452 39052 35541 39080
rect 35452 39024 35480 39052
rect 35529 39049 35541 39052
rect 35575 39049 35587 39083
rect 35529 39043 35587 39049
rect 35618 39040 35624 39092
rect 35676 39080 35682 39092
rect 35897 39083 35955 39089
rect 35897 39080 35909 39083
rect 35676 39052 35909 39080
rect 35676 39040 35682 39052
rect 35897 39049 35909 39052
rect 35943 39049 35955 39083
rect 35897 39043 35955 39049
rect 35986 39040 35992 39092
rect 36044 39040 36050 39092
rect 36357 39083 36415 39089
rect 36357 39049 36369 39083
rect 36403 39049 36415 39083
rect 36357 39043 36415 39049
rect 29914 39012 29920 39024
rect 28552 38984 29920 39012
rect 29914 38972 29920 38984
rect 29972 38972 29978 39024
rect 31573 39015 31631 39021
rect 31573 38981 31585 39015
rect 31619 39012 31631 39015
rect 32769 39015 32827 39021
rect 32769 39012 32781 39015
rect 31619 38984 32781 39012
rect 31619 38981 31631 38984
rect 31573 38975 31631 38981
rect 32769 38981 32781 38984
rect 32815 39012 32827 39015
rect 34330 39012 34336 39024
rect 32815 38984 34336 39012
rect 32815 38981 32827 38984
rect 32769 38975 32827 38981
rect 34330 38972 34336 38984
rect 34388 38972 34394 39024
rect 35434 38972 35440 39024
rect 35492 38972 35498 39024
rect 36078 39012 36084 39024
rect 35820 38984 36084 39012
rect 26329 38947 26387 38953
rect 26329 38913 26341 38947
rect 26375 38913 26387 38947
rect 26329 38907 26387 38913
rect 27709 38947 27767 38953
rect 27709 38913 27721 38947
rect 27755 38944 27767 38947
rect 27755 38916 28028 38944
rect 27755 38913 27767 38916
rect 27709 38907 27767 38913
rect 23385 38879 23443 38885
rect 23385 38845 23397 38879
rect 23431 38876 23443 38879
rect 24762 38876 24768 38888
rect 23431 38848 24768 38876
rect 23431 38845 23443 38848
rect 23385 38839 23443 38845
rect 24762 38836 24768 38848
rect 24820 38836 24826 38888
rect 24946 38836 24952 38888
rect 25004 38876 25010 38888
rect 25041 38879 25099 38885
rect 25041 38876 25053 38879
rect 25004 38848 25053 38876
rect 25004 38836 25010 38848
rect 25041 38845 25053 38848
rect 25087 38845 25099 38879
rect 25041 38839 25099 38845
rect 25866 38836 25872 38888
rect 25924 38876 25930 38888
rect 26421 38879 26479 38885
rect 26421 38876 26433 38879
rect 25924 38848 26433 38876
rect 25924 38836 25930 38848
rect 26421 38845 26433 38848
rect 26467 38845 26479 38879
rect 26421 38839 26479 38845
rect 27890 38836 27896 38888
rect 27948 38836 27954 38888
rect 25958 38768 25964 38820
rect 26016 38808 26022 38820
rect 26016 38780 27660 38808
rect 26016 38768 26022 38780
rect 1581 38743 1639 38749
rect 1581 38709 1593 38743
rect 1627 38740 1639 38743
rect 7374 38740 7380 38752
rect 1627 38712 7380 38740
rect 1627 38709 1639 38712
rect 1581 38703 1639 38709
rect 7374 38700 7380 38712
rect 7432 38700 7438 38752
rect 22833 38743 22891 38749
rect 22833 38709 22845 38743
rect 22879 38740 22891 38743
rect 27522 38740 27528 38752
rect 22879 38712 27528 38740
rect 22879 38709 22891 38712
rect 22833 38703 22891 38709
rect 27522 38700 27528 38712
rect 27580 38700 27586 38752
rect 27632 38740 27660 38780
rect 28000 38740 28028 38916
rect 28350 38904 28356 38956
rect 28408 38944 28414 38956
rect 28408 38916 29132 38944
rect 28408 38904 28414 38916
rect 28718 38836 28724 38888
rect 28776 38876 28782 38888
rect 29104 38885 29132 38916
rect 33318 38904 33324 38956
rect 33376 38944 33382 38956
rect 34057 38947 34115 38953
rect 34057 38944 34069 38947
rect 33376 38916 34069 38944
rect 33376 38904 33382 38916
rect 34057 38913 34069 38916
rect 34103 38913 34115 38947
rect 35820 38944 35848 38984
rect 36078 38972 36084 38984
rect 36136 38972 36142 39024
rect 36372 39012 36400 39043
rect 37274 39040 37280 39092
rect 37332 39080 37338 39092
rect 37921 39083 37979 39089
rect 37921 39080 37933 39083
rect 37332 39052 37933 39080
rect 37332 39040 37338 39052
rect 37921 39049 37933 39052
rect 37967 39049 37979 39083
rect 37921 39043 37979 39049
rect 38473 39083 38531 39089
rect 38473 39049 38485 39083
rect 38519 39080 38531 39083
rect 38838 39080 38844 39092
rect 38519 39052 38844 39080
rect 38519 39049 38531 39052
rect 38473 39043 38531 39049
rect 38838 39040 38844 39052
rect 38896 39040 38902 39092
rect 39114 39040 39120 39092
rect 39172 39080 39178 39092
rect 39301 39083 39359 39089
rect 39301 39080 39313 39083
rect 39172 39052 39313 39080
rect 39172 39040 39178 39052
rect 39301 39049 39313 39052
rect 39347 39049 39359 39083
rect 39301 39043 39359 39049
rect 39761 39083 39819 39089
rect 39761 39049 39773 39083
rect 39807 39080 39819 39083
rect 40126 39080 40132 39092
rect 39807 39052 40132 39080
rect 39807 39049 39819 39052
rect 39761 39043 39819 39049
rect 40126 39040 40132 39052
rect 40184 39080 40190 39092
rect 40402 39080 40408 39092
rect 40184 39052 40408 39080
rect 40184 39040 40190 39052
rect 40402 39040 40408 39052
rect 40460 39040 40466 39092
rect 36446 39012 36452 39024
rect 36372 38984 36452 39012
rect 36446 38972 36452 38984
rect 36504 38972 36510 39024
rect 36725 39015 36783 39021
rect 36725 38981 36737 39015
rect 36771 39012 36783 39015
rect 38286 39012 38292 39024
rect 36771 38984 38292 39012
rect 36771 38981 36783 38984
rect 36725 38975 36783 38981
rect 38286 38972 38292 38984
rect 38344 38972 38350 39024
rect 38562 38972 38568 39024
rect 38620 39012 38626 39024
rect 43438 39012 43444 39024
rect 38620 38984 40172 39012
rect 41814 38984 43444 39012
rect 38620 38972 38626 38984
rect 34057 38907 34115 38913
rect 34164 38916 35848 38944
rect 28997 38879 29055 38885
rect 28997 38876 29009 38879
rect 28776 38848 29009 38876
rect 28776 38836 28782 38848
rect 28997 38845 29009 38848
rect 29043 38845 29055 38879
rect 28997 38839 29055 38845
rect 29089 38879 29147 38885
rect 29089 38845 29101 38879
rect 29135 38845 29147 38879
rect 29089 38839 29147 38845
rect 31021 38879 31079 38885
rect 31021 38845 31033 38879
rect 31067 38876 31079 38879
rect 32861 38879 32919 38885
rect 32861 38876 32873 38879
rect 31067 38848 32873 38876
rect 31067 38845 31079 38848
rect 31021 38839 31079 38845
rect 32861 38845 32873 38848
rect 32907 38845 32919 38879
rect 32861 38839 32919 38845
rect 32953 38879 33011 38885
rect 32953 38845 32965 38879
rect 32999 38845 33011 38879
rect 34164 38876 34192 38916
rect 36170 38904 36176 38956
rect 36228 38944 36234 38956
rect 36817 38947 36875 38953
rect 36817 38944 36829 38947
rect 36228 38916 36829 38944
rect 36228 38904 36234 38916
rect 36817 38913 36829 38916
rect 36863 38913 36875 38947
rect 36817 38907 36875 38913
rect 37274 38904 37280 38956
rect 37332 38944 37338 38956
rect 37829 38947 37887 38953
rect 37829 38944 37841 38947
rect 37332 38916 37841 38944
rect 37332 38904 37338 38916
rect 37829 38913 37841 38916
rect 37875 38913 37887 38947
rect 37829 38907 37887 38913
rect 38838 38904 38844 38956
rect 38896 38904 38902 38956
rect 39390 38904 39396 38956
rect 39448 38944 39454 38956
rect 39669 38947 39727 38953
rect 39669 38944 39681 38947
rect 39448 38916 39681 38944
rect 39448 38904 39454 38916
rect 39669 38913 39681 38916
rect 39715 38913 39727 38947
rect 39669 38907 39727 38913
rect 32953 38839 33011 38845
rect 33704 38848 34192 38876
rect 28074 38768 28080 38820
rect 28132 38808 28138 38820
rect 28350 38808 28356 38820
rect 28132 38780 28356 38808
rect 28132 38768 28138 38780
rect 28350 38768 28356 38780
rect 28408 38808 28414 38820
rect 31036 38808 31064 38839
rect 28408 38780 31064 38808
rect 28408 38768 28414 38780
rect 31938 38768 31944 38820
rect 31996 38808 32002 38820
rect 32968 38808 32996 38839
rect 33704 38817 33732 38848
rect 34238 38836 34244 38888
rect 34296 38836 34302 38888
rect 34882 38836 34888 38888
rect 34940 38876 34946 38888
rect 36081 38879 36139 38885
rect 36081 38876 36093 38879
rect 34940 38848 36093 38876
rect 34940 38836 34946 38848
rect 36081 38845 36093 38848
rect 36127 38845 36139 38879
rect 36081 38839 36139 38845
rect 36909 38879 36967 38885
rect 36909 38845 36921 38879
rect 36955 38876 36967 38879
rect 37182 38876 37188 38888
rect 36955 38848 37188 38876
rect 36955 38845 36967 38848
rect 36909 38839 36967 38845
rect 31996 38780 32996 38808
rect 33689 38811 33747 38817
rect 31996 38768 32002 38780
rect 33689 38777 33701 38811
rect 33735 38777 33747 38811
rect 33689 38771 33747 38777
rect 33778 38768 33784 38820
rect 33836 38808 33842 38820
rect 36924 38808 36952 38839
rect 37182 38836 37188 38848
rect 37240 38836 37246 38888
rect 37734 38836 37740 38888
rect 37792 38876 37798 38888
rect 38013 38879 38071 38885
rect 38013 38876 38025 38879
rect 37792 38848 38025 38876
rect 37792 38836 37798 38848
rect 38013 38845 38025 38848
rect 38059 38845 38071 38879
rect 38013 38839 38071 38845
rect 38930 38836 38936 38888
rect 38988 38836 38994 38888
rect 39022 38836 39028 38888
rect 39080 38836 39086 38888
rect 39853 38879 39911 38885
rect 39853 38845 39865 38879
rect 39899 38876 39911 38879
rect 39942 38876 39948 38888
rect 39899 38848 39948 38876
rect 39899 38845 39911 38848
rect 39853 38839 39911 38845
rect 33836 38780 36952 38808
rect 37384 38780 37596 38808
rect 33836 38768 33842 38780
rect 27632 38712 28028 38740
rect 28534 38700 28540 38752
rect 28592 38700 28598 38752
rect 32398 38700 32404 38752
rect 32456 38700 32462 38752
rect 34974 38700 34980 38752
rect 35032 38740 35038 38752
rect 37384 38740 37412 38780
rect 35032 38712 37412 38740
rect 35032 38700 35038 38712
rect 37458 38700 37464 38752
rect 37516 38700 37522 38752
rect 37568 38740 37596 38780
rect 37826 38768 37832 38820
rect 37884 38808 37890 38820
rect 38470 38808 38476 38820
rect 37884 38780 38476 38808
rect 37884 38768 37890 38780
rect 38470 38768 38476 38780
rect 38528 38808 38534 38820
rect 39868 38808 39896 38839
rect 39942 38836 39948 38848
rect 40000 38836 40006 38888
rect 40144 38876 40172 38984
rect 43438 38972 43444 38984
rect 43496 38972 43502 39024
rect 40310 38876 40316 38888
rect 40144 38848 40316 38876
rect 40310 38836 40316 38848
rect 40368 38836 40374 38888
rect 40589 38879 40647 38885
rect 40589 38845 40601 38879
rect 40635 38876 40647 38879
rect 41046 38876 41052 38888
rect 40635 38848 41052 38876
rect 40635 38845 40647 38848
rect 40589 38839 40647 38845
rect 41046 38836 41052 38848
rect 41104 38836 41110 38888
rect 41230 38836 41236 38888
rect 41288 38876 41294 38888
rect 43898 38876 43904 38888
rect 41288 38848 43904 38876
rect 41288 38836 41294 38848
rect 43898 38836 43904 38848
rect 43956 38836 43962 38888
rect 38528 38780 39896 38808
rect 38528 38768 38534 38780
rect 40954 38740 40960 38752
rect 37568 38712 40960 38740
rect 40954 38700 40960 38712
rect 41012 38700 41018 38752
rect 41782 38700 41788 38752
rect 41840 38740 41846 38752
rect 42061 38743 42119 38749
rect 42061 38740 42073 38743
rect 41840 38712 42073 38740
rect 41840 38700 41846 38712
rect 42061 38709 42073 38712
rect 42107 38709 42119 38743
rect 42061 38703 42119 38709
rect 1104 38650 49864 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 32950 38650
rect 33002 38598 33014 38650
rect 33066 38598 33078 38650
rect 33130 38598 33142 38650
rect 33194 38598 33206 38650
rect 33258 38598 42950 38650
rect 43002 38598 43014 38650
rect 43066 38598 43078 38650
rect 43130 38598 43142 38650
rect 43194 38598 43206 38650
rect 43258 38598 49864 38650
rect 1104 38576 49864 38598
rect 22094 38496 22100 38548
rect 22152 38536 22158 38548
rect 23293 38539 23351 38545
rect 23293 38536 23305 38539
rect 22152 38508 23305 38536
rect 22152 38496 22158 38508
rect 23293 38505 23305 38508
rect 23339 38505 23351 38539
rect 23293 38499 23351 38505
rect 26326 38496 26332 38548
rect 26384 38536 26390 38548
rect 27065 38539 27123 38545
rect 27065 38536 27077 38539
rect 26384 38508 27077 38536
rect 26384 38496 26390 38508
rect 27065 38505 27077 38508
rect 27111 38505 27123 38539
rect 27065 38499 27123 38505
rect 27246 38496 27252 38548
rect 27304 38536 27310 38548
rect 31570 38536 31576 38548
rect 27304 38508 31576 38536
rect 27304 38496 27310 38508
rect 31570 38496 31576 38508
rect 31628 38496 31634 38548
rect 34422 38536 34428 38548
rect 31726 38508 34428 38536
rect 22833 38471 22891 38477
rect 22833 38437 22845 38471
rect 22879 38468 22891 38471
rect 25038 38468 25044 38480
rect 22879 38440 25044 38468
rect 22879 38437 22891 38440
rect 22833 38431 22891 38437
rect 25038 38428 25044 38440
rect 25096 38428 25102 38480
rect 26970 38428 26976 38480
rect 27028 38468 27034 38480
rect 28445 38471 28503 38477
rect 28445 38468 28457 38471
rect 27028 38440 28457 38468
rect 27028 38428 27034 38440
rect 28445 38437 28457 38440
rect 28491 38437 28503 38471
rect 28445 38431 28503 38437
rect 28626 38428 28632 38480
rect 28684 38468 28690 38480
rect 28684 38440 29040 38468
rect 28684 38428 28690 38440
rect 20714 38360 20720 38412
rect 20772 38400 20778 38412
rect 21082 38400 21088 38412
rect 20772 38372 21088 38400
rect 20772 38360 20778 38372
rect 21082 38360 21088 38372
rect 21140 38360 21146 38412
rect 22370 38360 22376 38412
rect 22428 38400 22434 38412
rect 23845 38403 23903 38409
rect 23845 38400 23857 38403
rect 22428 38372 23857 38400
rect 22428 38360 22434 38372
rect 23845 38369 23857 38372
rect 23891 38369 23903 38403
rect 23845 38363 23903 38369
rect 27522 38360 27528 38412
rect 27580 38360 27586 38412
rect 27617 38403 27675 38409
rect 27617 38369 27629 38403
rect 27663 38369 27675 38403
rect 27617 38363 27675 38369
rect 24762 38292 24768 38344
rect 24820 38332 24826 38344
rect 25038 38332 25044 38344
rect 24820 38304 25044 38332
rect 24820 38292 24826 38304
rect 25038 38292 25044 38304
rect 25096 38292 25102 38344
rect 26694 38292 26700 38344
rect 26752 38332 26758 38344
rect 27632 38332 27660 38363
rect 28534 38360 28540 38412
rect 28592 38400 28598 38412
rect 29012 38409 29040 38440
rect 31018 38428 31024 38480
rect 31076 38468 31082 38480
rect 31726 38468 31754 38508
rect 34422 38496 34428 38508
rect 34480 38496 34486 38548
rect 36630 38496 36636 38548
rect 36688 38496 36694 38548
rect 39206 38496 39212 38548
rect 39264 38496 39270 38548
rect 40037 38539 40095 38545
rect 40037 38505 40049 38539
rect 40083 38536 40095 38539
rect 41138 38536 41144 38548
rect 40083 38508 41144 38536
rect 40083 38505 40095 38508
rect 40037 38499 40095 38505
rect 41138 38496 41144 38508
rect 41196 38496 41202 38548
rect 41230 38496 41236 38548
rect 41288 38536 41294 38548
rect 49145 38539 49203 38545
rect 49145 38536 49157 38539
rect 41288 38508 49157 38536
rect 41288 38496 41294 38508
rect 49145 38505 49157 38508
rect 49191 38505 49203 38539
rect 49145 38499 49203 38505
rect 31076 38440 31754 38468
rect 33689 38471 33747 38477
rect 31076 38428 31082 38440
rect 33689 38437 33701 38471
rect 33735 38468 33747 38471
rect 34790 38468 34796 38480
rect 33735 38440 34796 38468
rect 33735 38437 33747 38440
rect 33689 38431 33747 38437
rect 34790 38428 34796 38440
rect 34848 38428 34854 38480
rect 39224 38468 39252 38496
rect 39482 38468 39488 38480
rect 39224 38440 39488 38468
rect 39482 38428 39488 38440
rect 39540 38468 39546 38480
rect 41322 38468 41328 38480
rect 39540 38440 41328 38468
rect 39540 38428 39546 38440
rect 28905 38403 28963 38409
rect 28905 38400 28917 38403
rect 28592 38372 28917 38400
rect 28592 38360 28598 38372
rect 28905 38369 28917 38372
rect 28951 38369 28963 38403
rect 28905 38363 28963 38369
rect 28997 38403 29055 38409
rect 28997 38369 29009 38403
rect 29043 38369 29055 38403
rect 28997 38363 29055 38369
rect 29472 38372 32536 38400
rect 26752 38304 27660 38332
rect 26752 38292 26758 38304
rect 27706 38292 27712 38344
rect 27764 38332 27770 38344
rect 29472 38332 29500 38372
rect 27764 38304 29500 38332
rect 27764 38292 27770 38304
rect 29730 38292 29736 38344
rect 29788 38292 29794 38344
rect 31662 38292 31668 38344
rect 31720 38332 31726 38344
rect 31849 38335 31907 38341
rect 31849 38332 31861 38335
rect 31720 38304 31861 38332
rect 31720 38292 31726 38304
rect 31849 38301 31861 38304
rect 31895 38301 31907 38335
rect 32508 38332 32536 38372
rect 32582 38360 32588 38412
rect 32640 38360 32646 38412
rect 32766 38360 32772 38412
rect 32824 38400 32830 38412
rect 33413 38403 33471 38409
rect 33413 38400 33425 38403
rect 32824 38372 33425 38400
rect 32824 38360 32830 38372
rect 33413 38369 33425 38372
rect 33459 38369 33471 38403
rect 33413 38363 33471 38369
rect 34146 38360 34152 38412
rect 34204 38360 34210 38412
rect 34241 38403 34299 38409
rect 34241 38369 34253 38403
rect 34287 38369 34299 38403
rect 34241 38363 34299 38369
rect 33321 38335 33379 38341
rect 33321 38332 33333 38335
rect 32508 38304 33333 38332
rect 31849 38295 31907 38301
rect 33321 38301 33333 38304
rect 33367 38301 33379 38335
rect 33321 38295 33379 38301
rect 21358 38224 21364 38276
rect 21416 38224 21422 38276
rect 22094 38224 22100 38276
rect 22152 38224 22158 38276
rect 23661 38267 23719 38273
rect 23661 38233 23673 38267
rect 23707 38264 23719 38267
rect 25130 38264 25136 38276
rect 23707 38236 25136 38264
rect 23707 38233 23719 38236
rect 23661 38227 23719 38233
rect 25130 38224 25136 38236
rect 25188 38224 25194 38276
rect 26605 38267 26663 38273
rect 26605 38233 26617 38267
rect 26651 38264 26663 38267
rect 27433 38267 27491 38273
rect 27433 38264 27445 38267
rect 26651 38236 27445 38264
rect 26651 38233 26663 38236
rect 26605 38227 26663 38233
rect 27433 38233 27445 38236
rect 27479 38264 27491 38267
rect 28534 38264 28540 38276
rect 27479 38236 28540 38264
rect 27479 38233 27491 38236
rect 27433 38227 27491 38233
rect 28534 38224 28540 38236
rect 28592 38224 28598 38276
rect 28813 38267 28871 38273
rect 28813 38233 28825 38267
rect 28859 38264 28871 38267
rect 29086 38264 29092 38276
rect 28859 38236 29092 38264
rect 28859 38233 28871 38236
rect 28813 38227 28871 38233
rect 29086 38224 29092 38236
rect 29144 38224 29150 38276
rect 30006 38224 30012 38276
rect 30064 38224 30070 38276
rect 30466 38224 30472 38276
rect 30524 38224 30530 38276
rect 31570 38224 31576 38276
rect 31628 38264 31634 38276
rect 31757 38267 31815 38273
rect 31757 38264 31769 38267
rect 31628 38236 31769 38264
rect 31628 38224 31634 38236
rect 31757 38233 31769 38236
rect 31803 38264 31815 38267
rect 31938 38264 31944 38276
rect 31803 38236 31944 38264
rect 31803 38233 31815 38236
rect 31757 38227 31815 38233
rect 31938 38224 31944 38236
rect 31996 38224 32002 38276
rect 32030 38224 32036 38276
rect 32088 38264 32094 38276
rect 34256 38264 34284 38363
rect 34698 38360 34704 38412
rect 34756 38400 34762 38412
rect 34885 38403 34943 38409
rect 34885 38400 34897 38403
rect 34756 38372 34897 38400
rect 34756 38360 34762 38372
rect 34885 38369 34897 38372
rect 34931 38369 34943 38403
rect 34885 38363 34943 38369
rect 35802 38360 35808 38412
rect 35860 38400 35866 38412
rect 35860 38372 36400 38400
rect 35860 38360 35866 38372
rect 32088 38236 34284 38264
rect 35161 38267 35219 38273
rect 32088 38224 32094 38236
rect 35161 38233 35173 38267
rect 35207 38264 35219 38267
rect 35250 38264 35256 38276
rect 35207 38236 35256 38264
rect 35207 38233 35219 38236
rect 35161 38227 35219 38233
rect 35250 38224 35256 38236
rect 35308 38224 35314 38276
rect 36372 38264 36400 38372
rect 38286 38360 38292 38412
rect 38344 38400 38350 38412
rect 38344 38372 39988 38400
rect 38344 38360 38350 38372
rect 39960 38332 39988 38372
rect 40420 38341 40448 38440
rect 41322 38428 41328 38440
rect 41380 38428 41386 38480
rect 42794 38428 42800 38480
rect 42852 38468 42858 38480
rect 43257 38471 43315 38477
rect 43257 38468 43269 38471
rect 42852 38440 43269 38468
rect 42852 38428 42858 38440
rect 43257 38437 43269 38440
rect 43303 38468 43315 38471
rect 43346 38468 43352 38480
rect 43303 38440 43352 38468
rect 43303 38437 43315 38440
rect 43257 38431 43315 38437
rect 43346 38428 43352 38440
rect 43404 38428 43410 38480
rect 40494 38360 40500 38412
rect 40552 38400 40558 38412
rect 40681 38403 40739 38409
rect 40681 38400 40693 38403
rect 40552 38372 40693 38400
rect 40552 38360 40558 38372
rect 40681 38369 40693 38372
rect 40727 38400 40739 38403
rect 41046 38400 41052 38412
rect 40727 38372 41052 38400
rect 40727 38369 40739 38372
rect 40681 38363 40739 38369
rect 41046 38360 41052 38372
rect 41104 38360 41110 38412
rect 48682 38400 48688 38412
rect 41386 38372 48688 38400
rect 40405 38335 40463 38341
rect 39960 38304 40264 38332
rect 36998 38264 37004 38276
rect 36372 38250 37004 38264
rect 36386 38236 37004 38250
rect 36998 38224 37004 38236
rect 37056 38224 37062 38276
rect 37090 38224 37096 38276
rect 37148 38224 37154 38276
rect 37921 38267 37979 38273
rect 37921 38233 37933 38267
rect 37967 38264 37979 38267
rect 38470 38264 38476 38276
rect 37967 38236 38476 38264
rect 37967 38233 37979 38236
rect 37921 38227 37979 38233
rect 38470 38224 38476 38236
rect 38528 38224 38534 38276
rect 40126 38264 40132 38276
rect 38580 38236 40132 38264
rect 23753 38199 23811 38205
rect 23753 38165 23765 38199
rect 23799 38196 23811 38199
rect 25498 38196 25504 38208
rect 23799 38168 25504 38196
rect 23799 38165 23811 38168
rect 23753 38159 23811 38165
rect 25498 38156 25504 38168
rect 25556 38156 25562 38208
rect 32214 38156 32220 38208
rect 32272 38196 32278 38208
rect 32861 38199 32919 38205
rect 32861 38196 32873 38199
rect 32272 38168 32873 38196
rect 32272 38156 32278 38168
rect 32861 38165 32873 38168
rect 32907 38165 32919 38199
rect 32861 38159 32919 38165
rect 33229 38199 33287 38205
rect 33229 38165 33241 38199
rect 33275 38196 33287 38199
rect 33962 38196 33968 38208
rect 33275 38168 33968 38196
rect 33275 38165 33287 38168
rect 33229 38159 33287 38165
rect 33962 38156 33968 38168
rect 34020 38156 34026 38208
rect 34054 38156 34060 38208
rect 34112 38156 34118 38208
rect 35066 38156 35072 38208
rect 35124 38196 35130 38208
rect 38580 38196 38608 38236
rect 40126 38224 40132 38236
rect 40184 38224 40190 38276
rect 35124 38168 38608 38196
rect 35124 38156 35130 38168
rect 39022 38156 39028 38208
rect 39080 38196 39086 38208
rect 39850 38196 39856 38208
rect 39080 38168 39856 38196
rect 39080 38156 39086 38168
rect 39850 38156 39856 38168
rect 39908 38156 39914 38208
rect 40236 38196 40264 38304
rect 40405 38301 40417 38335
rect 40451 38301 40463 38335
rect 41386 38332 41414 38372
rect 48682 38360 48688 38372
rect 48740 38360 48746 38412
rect 40405 38295 40463 38301
rect 41156 38304 41414 38332
rect 40497 38199 40555 38205
rect 40497 38196 40509 38199
rect 40236 38168 40509 38196
rect 40497 38165 40509 38168
rect 40543 38196 40555 38199
rect 41156 38196 41184 38304
rect 41506 38292 41512 38344
rect 41564 38292 41570 38344
rect 49326 38292 49332 38344
rect 49384 38292 49390 38344
rect 41782 38224 41788 38276
rect 41840 38224 41846 38276
rect 43438 38264 43444 38276
rect 43010 38236 43444 38264
rect 43438 38224 43444 38236
rect 43496 38224 43502 38276
rect 41233 38199 41291 38205
rect 41233 38196 41245 38199
rect 40543 38168 41245 38196
rect 40543 38165 40555 38168
rect 40497 38159 40555 38165
rect 41233 38165 41245 38168
rect 41279 38165 41291 38199
rect 41233 38159 41291 38165
rect 41322 38156 41328 38208
rect 41380 38196 41386 38208
rect 48866 38196 48872 38208
rect 41380 38168 48872 38196
rect 41380 38156 41386 38168
rect 48866 38156 48872 38168
rect 48924 38156 48930 38208
rect 1104 38106 49864 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 27950 38106
rect 28002 38054 28014 38106
rect 28066 38054 28078 38106
rect 28130 38054 28142 38106
rect 28194 38054 28206 38106
rect 28258 38054 37950 38106
rect 38002 38054 38014 38106
rect 38066 38054 38078 38106
rect 38130 38054 38142 38106
rect 38194 38054 38206 38106
rect 38258 38054 47950 38106
rect 48002 38054 48014 38106
rect 48066 38054 48078 38106
rect 48130 38054 48142 38106
rect 48194 38054 48206 38106
rect 48258 38054 49864 38106
rect 1104 38032 49864 38054
rect 24118 37992 24124 38004
rect 23768 37964 24124 37992
rect 22094 37884 22100 37936
rect 22152 37924 22158 37936
rect 23768 37924 23796 37964
rect 24118 37952 24124 37964
rect 24176 37952 24182 38004
rect 25038 37952 25044 38004
rect 25096 37992 25102 38004
rect 25096 37964 29224 37992
rect 25096 37952 25102 37964
rect 22152 37896 23874 37924
rect 22152 37884 22158 37896
rect 28166 37884 28172 37936
rect 28224 37884 28230 37936
rect 29196 37933 29224 37964
rect 29730 37952 29736 38004
rect 29788 37992 29794 38004
rect 29788 37964 31524 37992
rect 29788 37952 29794 37964
rect 29181 37927 29239 37933
rect 29181 37893 29193 37927
rect 29227 37893 29239 37927
rect 29181 37887 29239 37893
rect 29196 37856 29224 37887
rect 30650 37884 30656 37936
rect 30708 37884 30714 37936
rect 31018 37856 31024 37868
rect 29196 37828 31024 37856
rect 31018 37816 31024 37828
rect 31076 37816 31082 37868
rect 31496 37865 31524 37964
rect 33502 37952 33508 38004
rect 33560 37952 33566 38004
rect 33962 37952 33968 38004
rect 34020 37992 34026 38004
rect 41230 37992 41236 38004
rect 34020 37964 41236 37992
rect 34020 37952 34026 37964
rect 41230 37952 41236 37964
rect 41288 37952 41294 38004
rect 43162 37992 43168 38004
rect 41386 37964 43168 37992
rect 31662 37884 31668 37936
rect 31720 37924 31726 37936
rect 35989 37927 36047 37933
rect 35989 37924 36001 37927
rect 31720 37896 36001 37924
rect 31720 37884 31726 37896
rect 35989 37893 36001 37896
rect 36035 37924 36047 37927
rect 37090 37924 37096 37936
rect 36035 37896 37096 37924
rect 36035 37893 36047 37896
rect 35989 37887 36047 37893
rect 37090 37884 37096 37896
rect 37148 37884 37154 37936
rect 39574 37884 39580 37936
rect 39632 37884 39638 37936
rect 40126 37884 40132 37936
rect 40184 37924 40190 37936
rect 41386 37924 41414 37964
rect 43162 37952 43168 37964
rect 43220 37952 43226 38004
rect 49145 37995 49203 38001
rect 49145 37992 49157 37995
rect 45526 37964 49157 37992
rect 40184 37896 41414 37924
rect 40184 37884 40190 37896
rect 41966 37884 41972 37936
rect 42024 37924 42030 37936
rect 42981 37927 43039 37933
rect 42981 37924 42993 37927
rect 42024 37896 42993 37924
rect 42024 37884 42030 37896
rect 42981 37893 42993 37896
rect 43027 37924 43039 37927
rect 45526 37924 45554 37964
rect 49145 37961 49157 37964
rect 49191 37961 49203 37995
rect 49145 37955 49203 37961
rect 43027 37896 45554 37924
rect 43027 37893 43039 37896
rect 42981 37887 43039 37893
rect 31481 37859 31539 37865
rect 31481 37825 31493 37859
rect 31527 37856 31539 37859
rect 32306 37856 32312 37868
rect 31527 37828 32312 37856
rect 31527 37825 31539 37828
rect 31481 37819 31539 37825
rect 32306 37816 32312 37828
rect 32364 37816 32370 37868
rect 32674 37816 32680 37868
rect 32732 37856 32738 37868
rect 33045 37859 33103 37865
rect 33045 37856 33057 37859
rect 32732 37828 33057 37856
rect 32732 37816 32738 37828
rect 33045 37825 33057 37828
rect 33091 37856 33103 37859
rect 33870 37856 33876 37868
rect 33091 37828 33876 37856
rect 33091 37825 33103 37828
rect 33045 37819 33103 37825
rect 33870 37816 33876 37828
rect 33928 37816 33934 37868
rect 33980 37828 34652 37856
rect 23109 37791 23167 37797
rect 23109 37757 23121 37791
rect 23155 37757 23167 37791
rect 23109 37751 23167 37757
rect 23385 37791 23443 37797
rect 23385 37757 23397 37791
rect 23431 37788 23443 37791
rect 26694 37788 26700 37800
rect 23431 37760 26700 37788
rect 23431 37757 23443 37760
rect 23385 37751 23443 37757
rect 22462 37612 22468 37664
rect 22520 37652 22526 37664
rect 22649 37655 22707 37661
rect 22649 37652 22661 37655
rect 22520 37624 22661 37652
rect 22520 37612 22526 37624
rect 22649 37621 22661 37624
rect 22695 37621 22707 37655
rect 23124 37652 23152 37751
rect 26694 37748 26700 37760
rect 26752 37748 26758 37800
rect 26786 37748 26792 37800
rect 26844 37788 26850 37800
rect 27157 37791 27215 37797
rect 27157 37788 27169 37791
rect 26844 37760 27169 37788
rect 26844 37748 26850 37760
rect 27157 37757 27169 37760
rect 27203 37757 27215 37791
rect 27157 37751 27215 37757
rect 27433 37791 27491 37797
rect 27433 37757 27445 37791
rect 27479 37788 27491 37791
rect 27798 37788 27804 37800
rect 27479 37760 27804 37788
rect 27479 37757 27491 37760
rect 27433 37751 27491 37757
rect 27798 37748 27804 37760
rect 27856 37748 27862 37800
rect 28902 37748 28908 37800
rect 28960 37788 28966 37800
rect 30834 37788 30840 37800
rect 28960 37760 30840 37788
rect 28960 37748 28966 37760
rect 30834 37748 30840 37760
rect 30892 37748 30898 37800
rect 33410 37748 33416 37800
rect 33468 37788 33474 37800
rect 33980 37788 34008 37828
rect 33468 37760 34008 37788
rect 34057 37791 34115 37797
rect 33468 37748 33474 37760
rect 34057 37757 34069 37791
rect 34103 37757 34115 37791
rect 34057 37751 34115 37757
rect 28534 37680 28540 37732
rect 28592 37720 28598 37732
rect 28592 37692 31524 37720
rect 28592 37680 28598 37692
rect 24670 37652 24676 37664
rect 23124 37624 24676 37652
rect 22649 37615 22707 37621
rect 24670 37612 24676 37624
rect 24728 37612 24734 37664
rect 24857 37655 24915 37661
rect 24857 37621 24869 37655
rect 24903 37652 24915 37655
rect 24946 37652 24952 37664
rect 24903 37624 24952 37652
rect 24903 37621 24915 37624
rect 24857 37615 24915 37621
rect 24946 37612 24952 37624
rect 25004 37612 25010 37664
rect 30193 37655 30251 37661
rect 30193 37621 30205 37655
rect 30239 37652 30251 37655
rect 31294 37652 31300 37664
rect 30239 37624 31300 37652
rect 30239 37621 30251 37624
rect 30193 37615 30251 37621
rect 31294 37612 31300 37624
rect 31352 37612 31358 37664
rect 31496 37652 31524 37692
rect 31754 37680 31760 37732
rect 31812 37720 31818 37732
rect 34072 37720 34100 37751
rect 31812 37692 34100 37720
rect 34624 37720 34652 37828
rect 34698 37816 34704 37868
rect 34756 37856 34762 37868
rect 36725 37859 36783 37865
rect 36725 37856 36737 37859
rect 34756 37828 36737 37856
rect 34756 37816 34762 37828
rect 36725 37825 36737 37828
rect 36771 37825 36783 37859
rect 36725 37819 36783 37825
rect 41141 37859 41199 37865
rect 41141 37825 41153 37859
rect 41187 37856 41199 37859
rect 41187 37828 42932 37856
rect 41187 37825 41199 37828
rect 41141 37819 41199 37825
rect 38470 37748 38476 37800
rect 38528 37788 38534 37800
rect 38565 37791 38623 37797
rect 38565 37788 38577 37791
rect 38528 37760 38577 37788
rect 38528 37748 38534 37760
rect 38565 37757 38577 37760
rect 38611 37757 38623 37791
rect 38565 37751 38623 37757
rect 38841 37791 38899 37797
rect 38841 37757 38853 37791
rect 38887 37788 38899 37791
rect 39206 37788 39212 37800
rect 38887 37760 39212 37788
rect 38887 37757 38899 37760
rect 38841 37751 38899 37757
rect 39206 37748 39212 37760
rect 39264 37748 39270 37800
rect 41233 37791 41291 37797
rect 41233 37788 41245 37791
rect 39868 37760 41245 37788
rect 34624 37692 38700 37720
rect 31812 37680 31818 37692
rect 37642 37652 37648 37664
rect 31496 37624 37648 37652
rect 37642 37612 37648 37624
rect 37700 37612 37706 37664
rect 38672 37652 38700 37692
rect 39868 37652 39896 37760
rect 41233 37757 41245 37760
rect 41279 37757 41291 37791
rect 41233 37751 41291 37757
rect 41322 37748 41328 37800
rect 41380 37748 41386 37800
rect 42904 37788 42932 37828
rect 49326 37816 49332 37868
rect 49384 37816 49390 37868
rect 43073 37791 43131 37797
rect 43073 37788 43085 37791
rect 42904 37760 43085 37788
rect 43073 37757 43085 37760
rect 43119 37757 43131 37791
rect 43073 37751 43131 37757
rect 40126 37680 40132 37732
rect 40184 37720 40190 37732
rect 42613 37723 42671 37729
rect 42613 37720 42625 37723
rect 40184 37692 42625 37720
rect 40184 37680 40190 37692
rect 42613 37689 42625 37692
rect 42659 37689 42671 37723
rect 43088 37720 43116 37751
rect 43162 37748 43168 37800
rect 43220 37748 43226 37800
rect 46934 37720 46940 37732
rect 43088 37692 46940 37720
rect 42613 37683 42671 37689
rect 46934 37680 46940 37692
rect 46992 37680 46998 37732
rect 38672 37624 39896 37652
rect 39942 37612 39948 37664
rect 40000 37652 40006 37664
rect 40310 37652 40316 37664
rect 40000 37624 40316 37652
rect 40000 37612 40006 37624
rect 40310 37612 40316 37624
rect 40368 37612 40374 37664
rect 40773 37655 40831 37661
rect 40773 37621 40785 37655
rect 40819 37652 40831 37655
rect 42150 37652 42156 37664
rect 40819 37624 42156 37652
rect 40819 37621 40831 37624
rect 40773 37615 40831 37621
rect 42150 37612 42156 37624
rect 42208 37612 42214 37664
rect 42242 37612 42248 37664
rect 42300 37652 42306 37664
rect 44358 37652 44364 37664
rect 42300 37624 44364 37652
rect 42300 37612 42306 37624
rect 44358 37612 44364 37624
rect 44416 37612 44422 37664
rect 1104 37562 49864 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 32950 37562
rect 33002 37510 33014 37562
rect 33066 37510 33078 37562
rect 33130 37510 33142 37562
rect 33194 37510 33206 37562
rect 33258 37510 42950 37562
rect 43002 37510 43014 37562
rect 43066 37510 43078 37562
rect 43130 37510 43142 37562
rect 43194 37510 43206 37562
rect 43258 37510 49864 37562
rect 1104 37488 49864 37510
rect 21542 37408 21548 37460
rect 21600 37408 21606 37460
rect 27246 37448 27252 37460
rect 23952 37420 27252 37448
rect 21560 37312 21588 37408
rect 22741 37315 22799 37321
rect 21560 37284 22600 37312
rect 22462 37204 22468 37256
rect 22520 37204 22526 37256
rect 22572 37253 22600 37284
rect 22741 37281 22753 37315
rect 22787 37312 22799 37315
rect 23566 37312 23572 37324
rect 22787 37284 23572 37312
rect 22787 37281 22799 37284
rect 22741 37275 22799 37281
rect 23566 37272 23572 37284
rect 23624 37272 23630 37324
rect 23952 37321 23980 37420
rect 27246 37408 27252 37420
rect 27304 37408 27310 37460
rect 27798 37408 27804 37460
rect 27856 37448 27862 37460
rect 28537 37451 28595 37457
rect 28537 37448 28549 37451
rect 27856 37420 28549 37448
rect 27856 37408 27862 37420
rect 28537 37417 28549 37420
rect 28583 37417 28595 37451
rect 28537 37411 28595 37417
rect 30650 37408 30656 37460
rect 30708 37448 30714 37460
rect 31662 37448 31668 37460
rect 30708 37420 31668 37448
rect 30708 37408 30714 37420
rect 31662 37408 31668 37420
rect 31720 37408 31726 37460
rect 33870 37408 33876 37460
rect 33928 37448 33934 37460
rect 42242 37448 42248 37460
rect 33928 37420 42248 37448
rect 33928 37408 33934 37420
rect 42242 37408 42248 37420
rect 42300 37408 42306 37460
rect 42416 37451 42474 37457
rect 42416 37417 42428 37451
rect 42462 37448 42474 37451
rect 43530 37448 43536 37460
rect 42462 37420 43536 37448
rect 42462 37417 42474 37420
rect 42416 37411 42474 37417
rect 43530 37408 43536 37420
rect 43588 37408 43594 37460
rect 24670 37340 24676 37392
rect 24728 37380 24734 37392
rect 24728 37352 26556 37380
rect 24728 37340 24734 37352
rect 23937 37315 23995 37321
rect 23937 37281 23949 37315
rect 23983 37281 23995 37315
rect 23937 37275 23995 37281
rect 24578 37272 24584 37324
rect 24636 37312 24642 37324
rect 26053 37315 26111 37321
rect 26053 37312 26065 37315
rect 24636 37284 26065 37312
rect 24636 37272 24642 37284
rect 26053 37281 26065 37284
rect 26099 37281 26111 37315
rect 26053 37275 26111 37281
rect 22557 37247 22615 37253
rect 22557 37213 22569 37247
rect 22603 37244 22615 37247
rect 23290 37244 23296 37256
rect 22603 37216 23296 37244
rect 22603 37213 22615 37216
rect 22557 37207 22615 37213
rect 23290 37204 23296 37216
rect 23348 37204 23354 37256
rect 23661 37247 23719 37253
rect 23661 37213 23673 37247
rect 23707 37244 23719 37247
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 23707 37216 24777 37244
rect 23707 37213 23719 37216
rect 23661 37207 23719 37213
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 25961 37247 26019 37253
rect 25961 37244 25973 37247
rect 24765 37207 24823 37213
rect 24872 37216 25973 37244
rect 14458 37136 14464 37188
rect 14516 37176 14522 37188
rect 14516 37148 23796 37176
rect 14516 37136 14522 37148
rect 22097 37111 22155 37117
rect 22097 37077 22109 37111
rect 22143 37108 22155 37111
rect 22186 37108 22192 37120
rect 22143 37080 22192 37108
rect 22143 37077 22155 37080
rect 22097 37071 22155 37077
rect 22186 37068 22192 37080
rect 22244 37068 22250 37120
rect 23293 37111 23351 37117
rect 23293 37077 23305 37111
rect 23339 37108 23351 37111
rect 23474 37108 23480 37120
rect 23339 37080 23480 37108
rect 23339 37077 23351 37080
rect 23293 37071 23351 37077
rect 23474 37068 23480 37080
rect 23532 37068 23538 37120
rect 23768 37117 23796 37148
rect 24394 37136 24400 37188
rect 24452 37176 24458 37188
rect 24872 37176 24900 37216
rect 25961 37213 25973 37216
rect 26007 37213 26019 37247
rect 26528 37244 26556 37352
rect 29270 37340 29276 37392
rect 29328 37380 29334 37392
rect 29822 37380 29828 37392
rect 29328 37352 29828 37380
rect 29328 37340 29334 37352
rect 29822 37340 29828 37352
rect 29880 37380 29886 37392
rect 38102 37380 38108 37392
rect 29880 37352 31754 37380
rect 29880 37340 29886 37352
rect 27062 37272 27068 37324
rect 27120 37272 27126 37324
rect 27614 37272 27620 37324
rect 27672 37312 27678 37324
rect 28534 37312 28540 37324
rect 27672 37284 28540 37312
rect 27672 37272 27678 37284
rect 28534 37272 28540 37284
rect 28592 37272 28598 37324
rect 30285 37315 30343 37321
rect 30285 37281 30297 37315
rect 30331 37312 30343 37315
rect 31202 37312 31208 37324
rect 30331 37284 31208 37312
rect 30331 37281 30343 37284
rect 30285 37275 30343 37281
rect 31202 37272 31208 37284
rect 31260 37272 31266 37324
rect 31478 37272 31484 37324
rect 31536 37272 31542 37324
rect 31726 37312 31754 37352
rect 37476 37352 38108 37380
rect 37476 37321 37504 37352
rect 38102 37340 38108 37352
rect 38160 37340 38166 37392
rect 38562 37340 38568 37392
rect 38620 37340 38626 37392
rect 39758 37340 39764 37392
rect 39816 37380 39822 37392
rect 39942 37380 39948 37392
rect 39816 37352 39948 37380
rect 39816 37340 39822 37352
rect 39942 37340 39948 37352
rect 40000 37340 40006 37392
rect 40034 37340 40040 37392
rect 40092 37340 40098 37392
rect 40678 37380 40684 37392
rect 40144 37352 40684 37380
rect 32677 37315 32735 37321
rect 32677 37312 32689 37315
rect 31726 37284 32689 37312
rect 32677 37281 32689 37284
rect 32723 37281 32735 37315
rect 32677 37275 32735 37281
rect 37461 37315 37519 37321
rect 37461 37281 37473 37315
rect 37507 37281 37519 37315
rect 37461 37275 37519 37281
rect 37550 37272 37556 37324
rect 37608 37272 37614 37324
rect 39206 37272 39212 37324
rect 39264 37312 39270 37324
rect 39264 37284 39712 37312
rect 39264 37272 39270 37284
rect 26786 37244 26792 37256
rect 26528 37216 26792 37244
rect 25961 37207 26019 37213
rect 26786 37204 26792 37216
rect 26844 37204 26850 37256
rect 28166 37204 28172 37256
rect 28224 37244 28230 37256
rect 28626 37244 28632 37256
rect 28224 37216 28632 37244
rect 28224 37204 28230 37216
rect 28626 37204 28632 37216
rect 28684 37204 28690 37256
rect 29181 37247 29239 37253
rect 29181 37213 29193 37247
rect 29227 37244 29239 37247
rect 30101 37247 30159 37253
rect 30101 37244 30113 37247
rect 29227 37216 30113 37244
rect 29227 37213 29239 37216
rect 29181 37207 29239 37213
rect 30101 37213 30113 37216
rect 30147 37213 30159 37247
rect 30101 37207 30159 37213
rect 31294 37204 31300 37256
rect 31352 37204 31358 37256
rect 32490 37204 32496 37256
rect 32548 37244 32554 37256
rect 32585 37247 32643 37253
rect 32585 37244 32597 37247
rect 32548 37216 32597 37244
rect 32548 37204 32554 37216
rect 32585 37213 32597 37216
rect 32631 37213 32643 37247
rect 32585 37207 32643 37213
rect 37090 37204 37096 37256
rect 37148 37244 37154 37256
rect 37369 37247 37427 37253
rect 37369 37244 37381 37247
rect 37148 37216 37381 37244
rect 37148 37204 37154 37216
rect 37369 37213 37381 37216
rect 37415 37213 37427 37247
rect 38933 37247 38991 37253
rect 38933 37244 38945 37247
rect 37369 37207 37427 37213
rect 37568 37216 38945 37244
rect 37568 37188 37596 37216
rect 38933 37213 38945 37216
rect 38979 37244 38991 37247
rect 39114 37244 39120 37256
rect 38979 37216 39120 37244
rect 38979 37213 38991 37216
rect 38933 37207 38991 37213
rect 39114 37204 39120 37216
rect 39172 37204 39178 37256
rect 39684 37244 39712 37284
rect 40144 37244 40172 37352
rect 40678 37340 40684 37352
rect 40736 37340 40742 37392
rect 40310 37272 40316 37324
rect 40368 37312 40374 37324
rect 40589 37315 40647 37321
rect 40589 37312 40601 37315
rect 40368 37284 40601 37312
rect 40368 37272 40374 37284
rect 40589 37281 40601 37284
rect 40635 37281 40647 37315
rect 40589 37275 40647 37281
rect 41506 37272 41512 37324
rect 41564 37312 41570 37324
rect 42153 37315 42211 37321
rect 42153 37312 42165 37315
rect 41564 37284 42165 37312
rect 41564 37272 41570 37284
rect 42153 37281 42165 37284
rect 42199 37312 42211 37315
rect 42518 37312 42524 37324
rect 42199 37284 42524 37312
rect 42199 37281 42211 37284
rect 42153 37275 42211 37281
rect 42518 37272 42524 37284
rect 42576 37272 42582 37324
rect 48041 37315 48099 37321
rect 48041 37281 48053 37315
rect 48087 37312 48099 37315
rect 48498 37312 48504 37324
rect 48087 37284 48504 37312
rect 48087 37281 48099 37284
rect 48041 37275 48099 37281
rect 48498 37272 48504 37284
rect 48556 37272 48562 37324
rect 39684 37216 40172 37244
rect 40218 37204 40224 37256
rect 40276 37244 40282 37256
rect 40497 37247 40555 37253
rect 40497 37244 40509 37247
rect 40276 37216 40509 37244
rect 40276 37204 40282 37216
rect 40497 37213 40509 37216
rect 40543 37213 40555 37247
rect 40497 37207 40555 37213
rect 41414 37204 41420 37256
rect 41472 37204 41478 37256
rect 48774 37204 48780 37256
rect 48832 37204 48838 37256
rect 24452 37148 24900 37176
rect 25869 37179 25927 37185
rect 24452 37136 24458 37148
rect 25869 37145 25881 37179
rect 25915 37176 25927 37179
rect 26970 37176 26976 37188
rect 25915 37148 26976 37176
rect 25915 37145 25927 37148
rect 25869 37139 25927 37145
rect 26970 37136 26976 37148
rect 27028 37136 27034 37188
rect 33318 37176 33324 37188
rect 29748 37148 33324 37176
rect 23753 37111 23811 37117
rect 23753 37077 23765 37111
rect 23799 37108 23811 37111
rect 25406 37108 25412 37120
rect 23799 37080 25412 37108
rect 23799 37077 23811 37080
rect 23753 37071 23811 37077
rect 25406 37068 25412 37080
rect 25464 37068 25470 37120
rect 25498 37068 25504 37120
rect 25556 37068 25562 37120
rect 29748 37117 29776 37148
rect 33318 37136 33324 37148
rect 33376 37136 33382 37188
rect 37550 37136 37556 37188
rect 37608 37136 37614 37188
rect 38562 37136 38568 37188
rect 38620 37176 38626 37188
rect 40405 37179 40463 37185
rect 40405 37176 40417 37179
rect 38620 37148 40417 37176
rect 38620 37136 38626 37148
rect 40405 37145 40417 37148
rect 40451 37145 40463 37179
rect 40405 37139 40463 37145
rect 40678 37136 40684 37188
rect 40736 37176 40742 37188
rect 40736 37148 41736 37176
rect 40736 37136 40742 37148
rect 29733 37111 29791 37117
rect 29733 37077 29745 37111
rect 29779 37077 29791 37111
rect 29733 37071 29791 37077
rect 29822 37068 29828 37120
rect 29880 37108 29886 37120
rect 30193 37111 30251 37117
rect 30193 37108 30205 37111
rect 29880 37080 30205 37108
rect 29880 37068 29886 37080
rect 30193 37077 30205 37080
rect 30239 37077 30251 37111
rect 30193 37071 30251 37077
rect 30742 37068 30748 37120
rect 30800 37108 30806 37120
rect 30929 37111 30987 37117
rect 30929 37108 30941 37111
rect 30800 37080 30941 37108
rect 30800 37068 30806 37080
rect 30929 37077 30941 37080
rect 30975 37077 30987 37111
rect 30929 37071 30987 37077
rect 31110 37068 31116 37120
rect 31168 37108 31174 37120
rect 31389 37111 31447 37117
rect 31389 37108 31401 37111
rect 31168 37080 31401 37108
rect 31168 37068 31174 37080
rect 31389 37077 31401 37080
rect 31435 37077 31447 37111
rect 31389 37071 31447 37077
rect 32122 37068 32128 37120
rect 32180 37068 32186 37120
rect 32490 37068 32496 37120
rect 32548 37068 32554 37120
rect 34238 37068 34244 37120
rect 34296 37108 34302 37120
rect 34422 37108 34428 37120
rect 34296 37080 34428 37108
rect 34296 37068 34302 37080
rect 34422 37068 34428 37080
rect 34480 37108 34486 37120
rect 36906 37108 36912 37120
rect 34480 37080 36912 37108
rect 34480 37068 34486 37080
rect 36906 37068 36912 37080
rect 36964 37068 36970 37120
rect 37001 37111 37059 37117
rect 37001 37077 37013 37111
rect 37047 37108 37059 37111
rect 37274 37108 37280 37120
rect 37047 37080 37280 37108
rect 37047 37077 37059 37080
rect 37001 37071 37059 37077
rect 37274 37068 37280 37080
rect 37332 37068 37338 37120
rect 38102 37068 38108 37120
rect 38160 37108 38166 37120
rect 39025 37111 39083 37117
rect 39025 37108 39037 37111
rect 38160 37080 39037 37108
rect 38160 37068 38166 37080
rect 39025 37077 39037 37080
rect 39071 37108 39083 37111
rect 41598 37108 41604 37120
rect 39071 37080 41604 37108
rect 39071 37077 39083 37080
rect 39025 37071 39083 37077
rect 41598 37068 41604 37080
rect 41656 37068 41662 37120
rect 41708 37108 41736 37148
rect 43438 37136 43444 37188
rect 43496 37136 43502 37188
rect 43901 37111 43959 37117
rect 43901 37108 43913 37111
rect 41708 37080 43913 37108
rect 43901 37077 43913 37080
rect 43947 37077 43959 37111
rect 43901 37071 43959 37077
rect 1104 37018 49864 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 27950 37018
rect 28002 36966 28014 37018
rect 28066 36966 28078 37018
rect 28130 36966 28142 37018
rect 28194 36966 28206 37018
rect 28258 36966 37950 37018
rect 38002 36966 38014 37018
rect 38066 36966 38078 37018
rect 38130 36966 38142 37018
rect 38194 36966 38206 37018
rect 38258 36966 47950 37018
rect 48002 36966 48014 37018
rect 48066 36966 48078 37018
rect 48130 36966 48142 37018
rect 48194 36966 48206 37018
rect 48258 36966 49864 37018
rect 1104 36944 49864 36966
rect 19426 36864 19432 36916
rect 19484 36864 19490 36916
rect 26237 36907 26295 36913
rect 26237 36873 26249 36907
rect 26283 36904 26295 36907
rect 32030 36904 32036 36916
rect 26283 36876 32036 36904
rect 26283 36873 26295 36876
rect 26237 36867 26295 36873
rect 32030 36864 32036 36876
rect 32088 36864 32094 36916
rect 32309 36907 32367 36913
rect 32309 36873 32321 36907
rect 32355 36873 32367 36907
rect 32309 36867 32367 36873
rect 21818 36796 21824 36848
rect 21876 36836 21882 36848
rect 22094 36836 22100 36848
rect 21876 36808 22100 36836
rect 21876 36796 21882 36808
rect 22094 36796 22100 36808
rect 22152 36796 22158 36848
rect 24118 36796 24124 36848
rect 24176 36796 24182 36848
rect 26329 36839 26387 36845
rect 26329 36805 26341 36839
rect 26375 36836 26387 36839
rect 26375 36808 30420 36836
rect 26375 36805 26387 36808
rect 26329 36799 26387 36805
rect 934 36728 940 36780
rect 992 36768 998 36780
rect 1765 36771 1823 36777
rect 1765 36768 1777 36771
rect 992 36740 1777 36768
rect 992 36728 998 36740
rect 1765 36737 1777 36740
rect 1811 36737 1823 36771
rect 1765 36731 1823 36737
rect 17218 36728 17224 36780
rect 17276 36768 17282 36780
rect 19797 36771 19855 36777
rect 19797 36768 19809 36771
rect 17276 36740 19809 36768
rect 17276 36728 17282 36740
rect 19797 36737 19809 36740
rect 19843 36737 19855 36771
rect 19797 36731 19855 36737
rect 19889 36771 19947 36777
rect 19889 36737 19901 36771
rect 19935 36768 19947 36771
rect 22002 36768 22008 36780
rect 19935 36740 22008 36768
rect 19935 36737 19947 36740
rect 19889 36731 19947 36737
rect 22002 36728 22008 36740
rect 22060 36728 22066 36780
rect 22646 36728 22652 36780
rect 22704 36768 22710 36780
rect 23385 36771 23443 36777
rect 23385 36768 23397 36771
rect 22704 36740 23397 36768
rect 22704 36728 22710 36740
rect 23385 36737 23397 36740
rect 23431 36737 23443 36771
rect 23385 36731 23443 36737
rect 25498 36728 25504 36780
rect 25556 36768 25562 36780
rect 25556 36740 26556 36768
rect 25556 36728 25562 36740
rect 20073 36703 20131 36709
rect 20073 36669 20085 36703
rect 20119 36700 20131 36703
rect 21358 36700 21364 36712
rect 20119 36672 21364 36700
rect 20119 36669 20131 36672
rect 20073 36663 20131 36669
rect 21358 36660 21364 36672
rect 21416 36660 21422 36712
rect 23661 36703 23719 36709
rect 23661 36669 23673 36703
rect 23707 36700 23719 36703
rect 24946 36700 24952 36712
rect 23707 36672 24952 36700
rect 23707 36669 23719 36672
rect 23661 36663 23719 36669
rect 24946 36660 24952 36672
rect 25004 36660 25010 36712
rect 25409 36703 25467 36709
rect 25409 36669 25421 36703
rect 25455 36700 25467 36703
rect 25590 36700 25596 36712
rect 25455 36672 25596 36700
rect 25455 36669 25467 36672
rect 25409 36663 25467 36669
rect 25590 36660 25596 36672
rect 25648 36660 25654 36712
rect 26418 36660 26424 36712
rect 26476 36660 26482 36712
rect 26528 36700 26556 36740
rect 27522 36728 27528 36780
rect 27580 36728 27586 36780
rect 28718 36728 28724 36780
rect 28776 36768 28782 36780
rect 30285 36771 30343 36777
rect 30285 36768 30297 36771
rect 28776 36740 30297 36768
rect 28776 36728 28782 36740
rect 30285 36737 30297 36740
rect 30331 36737 30343 36771
rect 30392 36768 30420 36808
rect 30466 36796 30472 36848
rect 30524 36836 30530 36848
rect 32324 36836 32352 36867
rect 32398 36864 32404 36916
rect 32456 36904 32462 36916
rect 32769 36907 32827 36913
rect 32769 36904 32781 36907
rect 32456 36876 32781 36904
rect 32456 36864 32462 36876
rect 32769 36873 32781 36876
rect 32815 36873 32827 36907
rect 32769 36867 32827 36873
rect 34882 36864 34888 36916
rect 34940 36864 34946 36916
rect 37366 36864 37372 36916
rect 37424 36904 37430 36916
rect 37829 36907 37887 36913
rect 37829 36904 37841 36907
rect 37424 36876 37841 36904
rect 37424 36864 37430 36876
rect 37829 36873 37841 36876
rect 37875 36873 37887 36907
rect 41506 36904 41512 36916
rect 37829 36867 37887 36873
rect 39776 36876 41512 36904
rect 30524 36808 32352 36836
rect 32677 36839 32735 36845
rect 30524 36796 30530 36808
rect 32677 36805 32689 36839
rect 32723 36836 32735 36839
rect 34900 36836 34928 36864
rect 32723 36808 34928 36836
rect 32723 36805 32735 36808
rect 32677 36799 32735 36805
rect 39114 36796 39120 36848
rect 39172 36836 39178 36848
rect 39666 36836 39672 36848
rect 39172 36808 39672 36836
rect 39172 36796 39178 36808
rect 39666 36796 39672 36808
rect 39724 36796 39730 36848
rect 32214 36768 32220 36780
rect 30392 36740 32220 36768
rect 30285 36731 30343 36737
rect 32214 36728 32220 36740
rect 32272 36728 32278 36780
rect 35802 36728 35808 36780
rect 35860 36728 35866 36780
rect 38838 36728 38844 36780
rect 38896 36768 38902 36780
rect 39209 36771 39267 36777
rect 39209 36768 39221 36771
rect 38896 36740 39221 36768
rect 38896 36728 38902 36740
rect 39209 36737 39221 36740
rect 39255 36737 39267 36771
rect 39209 36731 39267 36737
rect 27617 36703 27675 36709
rect 27617 36700 27629 36703
rect 26528 36672 27629 36700
rect 27617 36669 27629 36672
rect 27663 36669 27675 36703
rect 27617 36663 27675 36669
rect 27801 36703 27859 36709
rect 27801 36669 27813 36703
rect 27847 36700 27859 36703
rect 29362 36700 29368 36712
rect 27847 36672 29368 36700
rect 27847 36669 27859 36672
rect 27801 36663 27859 36669
rect 29362 36660 29368 36672
rect 29420 36660 29426 36712
rect 30377 36703 30435 36709
rect 30377 36669 30389 36703
rect 30423 36669 30435 36703
rect 30377 36663 30435 36669
rect 30561 36703 30619 36709
rect 30561 36669 30573 36703
rect 30607 36669 30619 36703
rect 30561 36663 30619 36669
rect 29178 36592 29184 36644
rect 29236 36632 29242 36644
rect 29917 36635 29975 36641
rect 29917 36632 29929 36635
rect 29236 36604 29929 36632
rect 29236 36592 29242 36604
rect 29917 36601 29929 36604
rect 29963 36601 29975 36635
rect 29917 36595 29975 36601
rect 1581 36567 1639 36573
rect 1581 36533 1593 36567
rect 1627 36564 1639 36567
rect 7558 36564 7564 36576
rect 1627 36536 7564 36564
rect 1627 36533 1639 36536
rect 1581 36527 1639 36533
rect 7558 36524 7564 36536
rect 7616 36524 7622 36576
rect 22925 36567 22983 36573
rect 22925 36533 22937 36567
rect 22971 36564 22983 36567
rect 23658 36564 23664 36576
rect 22971 36536 23664 36564
rect 22971 36533 22983 36536
rect 22925 36527 22983 36533
rect 23658 36524 23664 36536
rect 23716 36524 23722 36576
rect 25866 36524 25872 36576
rect 25924 36524 25930 36576
rect 27157 36567 27215 36573
rect 27157 36533 27169 36567
rect 27203 36564 27215 36567
rect 29454 36564 29460 36576
rect 27203 36536 29460 36564
rect 27203 36533 27215 36536
rect 27157 36527 27215 36533
rect 29454 36524 29460 36536
rect 29512 36524 29518 36576
rect 30392 36564 30420 36663
rect 30576 36632 30604 36663
rect 31662 36660 31668 36712
rect 31720 36700 31726 36712
rect 31757 36703 31815 36709
rect 31757 36700 31769 36703
rect 31720 36672 31769 36700
rect 31720 36660 31726 36672
rect 31757 36669 31769 36672
rect 31803 36669 31815 36703
rect 31757 36663 31815 36669
rect 32306 36660 32312 36712
rect 32364 36700 32370 36712
rect 32861 36703 32919 36709
rect 32861 36700 32873 36703
rect 32364 36672 32873 36700
rect 32364 36660 32370 36672
rect 32861 36669 32873 36672
rect 32907 36669 32919 36703
rect 32861 36663 32919 36669
rect 33962 36660 33968 36712
rect 34020 36700 34026 36712
rect 34425 36703 34483 36709
rect 34425 36700 34437 36703
rect 34020 36672 34437 36700
rect 34020 36660 34026 36672
rect 34425 36669 34437 36672
rect 34471 36669 34483 36703
rect 34425 36663 34483 36669
rect 34701 36703 34759 36709
rect 34701 36669 34713 36703
rect 34747 36700 34759 36703
rect 35066 36700 35072 36712
rect 34747 36672 35072 36700
rect 34747 36669 34759 36672
rect 34701 36663 34759 36669
rect 35066 36660 35072 36672
rect 35124 36660 35130 36712
rect 37366 36660 37372 36712
rect 37424 36700 37430 36712
rect 37921 36703 37979 36709
rect 37921 36700 37933 36703
rect 37424 36672 37933 36700
rect 37424 36660 37430 36672
rect 37921 36669 37933 36672
rect 37967 36669 37979 36703
rect 37921 36663 37979 36669
rect 38105 36703 38163 36709
rect 38105 36669 38117 36703
rect 38151 36669 38163 36703
rect 38105 36663 38163 36669
rect 33870 36632 33876 36644
rect 30576 36604 33876 36632
rect 33870 36592 33876 36604
rect 33928 36592 33934 36644
rect 37461 36635 37519 36641
rect 37461 36632 37473 36635
rect 35728 36604 37473 36632
rect 35066 36564 35072 36576
rect 30392 36536 35072 36564
rect 35066 36524 35072 36536
rect 35124 36524 35130 36576
rect 35158 36524 35164 36576
rect 35216 36564 35222 36576
rect 35728 36564 35756 36604
rect 37461 36601 37473 36604
rect 37507 36601 37519 36635
rect 38120 36632 38148 36663
rect 38470 36660 38476 36712
rect 38528 36700 38534 36712
rect 39776 36709 39804 36876
rect 41506 36864 41512 36876
rect 41564 36864 41570 36916
rect 41598 36864 41604 36916
rect 41656 36904 41662 36916
rect 48958 36904 48964 36916
rect 41656 36876 48964 36904
rect 41656 36864 41662 36876
rect 48958 36864 48964 36876
rect 49016 36864 49022 36916
rect 39942 36796 39948 36848
rect 40000 36836 40006 36848
rect 40037 36839 40095 36845
rect 40037 36836 40049 36839
rect 40000 36808 40049 36836
rect 40000 36796 40006 36808
rect 40037 36805 40049 36808
rect 40083 36805 40095 36839
rect 40037 36799 40095 36805
rect 42702 36796 42708 36848
rect 42760 36836 42766 36848
rect 43073 36839 43131 36845
rect 43073 36836 43085 36839
rect 42760 36808 43085 36836
rect 42760 36796 42766 36808
rect 43073 36805 43085 36808
rect 43119 36805 43131 36839
rect 43073 36799 43131 36805
rect 39761 36703 39819 36709
rect 39761 36700 39773 36703
rect 38528 36672 39773 36700
rect 38528 36660 38534 36672
rect 39761 36669 39773 36672
rect 39807 36669 39819 36703
rect 41156 36700 41184 36754
rect 41322 36728 41328 36780
rect 41380 36768 41386 36780
rect 42981 36771 43039 36777
rect 42981 36768 42993 36771
rect 41380 36740 42993 36768
rect 41380 36728 41386 36740
rect 42981 36737 42993 36740
rect 43027 36737 43039 36771
rect 42981 36731 43039 36737
rect 49326 36728 49332 36780
rect 49384 36728 49390 36780
rect 43257 36703 43315 36709
rect 39761 36663 39819 36669
rect 39868 36672 42840 36700
rect 38562 36632 38568 36644
rect 38120 36604 38568 36632
rect 37461 36595 37519 36601
rect 38562 36592 38568 36604
rect 38620 36592 38626 36644
rect 39666 36592 39672 36644
rect 39724 36632 39730 36644
rect 39868 36632 39896 36672
rect 39724 36604 39896 36632
rect 42812 36632 42840 36672
rect 43257 36669 43269 36703
rect 43303 36700 43315 36703
rect 43346 36700 43352 36712
rect 43303 36672 43352 36700
rect 43303 36669 43315 36672
rect 43257 36663 43315 36669
rect 43346 36660 43352 36672
rect 43404 36660 43410 36712
rect 43438 36632 43444 36644
rect 42812 36604 43444 36632
rect 39724 36592 39730 36604
rect 43438 36592 43444 36604
rect 43496 36592 43502 36644
rect 35216 36536 35756 36564
rect 36173 36567 36231 36573
rect 35216 36524 35222 36536
rect 36173 36533 36185 36567
rect 36219 36564 36231 36567
rect 36722 36564 36728 36576
rect 36219 36536 36728 36564
rect 36219 36533 36231 36536
rect 36173 36527 36231 36533
rect 36722 36524 36728 36536
rect 36780 36524 36786 36576
rect 36906 36524 36912 36576
rect 36964 36564 36970 36576
rect 38010 36564 38016 36576
rect 36964 36536 38016 36564
rect 36964 36524 36970 36536
rect 38010 36524 38016 36536
rect 38068 36524 38074 36576
rect 41046 36524 41052 36576
rect 41104 36564 41110 36576
rect 41509 36567 41567 36573
rect 41509 36564 41521 36567
rect 41104 36536 41521 36564
rect 41104 36524 41110 36536
rect 41509 36533 41521 36536
rect 41555 36533 41567 36567
rect 41509 36527 41567 36533
rect 42518 36524 42524 36576
rect 42576 36564 42582 36576
rect 42613 36567 42671 36573
rect 42613 36564 42625 36567
rect 42576 36536 42625 36564
rect 42576 36524 42582 36536
rect 42613 36533 42625 36536
rect 42659 36533 42671 36567
rect 42613 36527 42671 36533
rect 46934 36524 46940 36576
rect 46992 36564 46998 36576
rect 49145 36567 49203 36573
rect 49145 36564 49157 36567
rect 46992 36536 49157 36564
rect 46992 36524 46998 36536
rect 49145 36533 49157 36536
rect 49191 36533 49203 36567
rect 49145 36527 49203 36533
rect 1104 36474 49864 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 32950 36474
rect 33002 36422 33014 36474
rect 33066 36422 33078 36474
rect 33130 36422 33142 36474
rect 33194 36422 33206 36474
rect 33258 36422 42950 36474
rect 43002 36422 43014 36474
rect 43066 36422 43078 36474
rect 43130 36422 43142 36474
rect 43194 36422 43206 36474
rect 43258 36422 49864 36474
rect 1104 36400 49864 36422
rect 22281 36363 22339 36369
rect 22281 36329 22293 36363
rect 22327 36360 22339 36363
rect 22370 36360 22376 36372
rect 22327 36332 22376 36360
rect 22327 36329 22339 36332
rect 22281 36323 22339 36329
rect 22370 36320 22376 36332
rect 22428 36320 22434 36372
rect 23293 36363 23351 36369
rect 23293 36329 23305 36363
rect 23339 36360 23351 36363
rect 26234 36360 26240 36372
rect 23339 36332 26240 36360
rect 23339 36329 23351 36332
rect 23293 36323 23351 36329
rect 26234 36320 26240 36332
rect 26292 36320 26298 36372
rect 27522 36320 27528 36372
rect 27580 36360 27586 36372
rect 27617 36363 27675 36369
rect 27617 36360 27629 36363
rect 27580 36332 27629 36360
rect 27580 36320 27586 36332
rect 27617 36329 27629 36332
rect 27663 36329 27675 36363
rect 27617 36323 27675 36329
rect 29454 36320 29460 36372
rect 29512 36360 29518 36372
rect 29512 36332 31984 36360
rect 29512 36320 29518 36332
rect 21910 36252 21916 36304
rect 21968 36292 21974 36304
rect 23566 36292 23572 36304
rect 21968 36264 23572 36292
rect 21968 36252 21974 36264
rect 23566 36252 23572 36264
rect 23624 36252 23630 36304
rect 31846 36292 31852 36304
rect 28184 36264 31852 36292
rect 20530 36184 20536 36236
rect 20588 36184 20594 36236
rect 23382 36184 23388 36236
rect 23440 36224 23446 36236
rect 23937 36227 23995 36233
rect 23440 36196 23796 36224
rect 23440 36184 23446 36196
rect 23658 36116 23664 36168
rect 23716 36116 23722 36168
rect 23768 36156 23796 36196
rect 23937 36193 23949 36227
rect 23983 36224 23995 36227
rect 24302 36224 24308 36236
rect 23983 36196 24308 36224
rect 23983 36193 23995 36196
rect 23937 36187 23995 36193
rect 24302 36184 24308 36196
rect 24360 36184 24366 36236
rect 26602 36156 26608 36168
rect 23768 36128 26608 36156
rect 26602 36116 26608 36128
rect 26660 36116 26666 36168
rect 28184 36165 28212 36264
rect 31846 36252 31852 36264
rect 31904 36252 31910 36304
rect 31956 36292 31984 36332
rect 32030 36320 32036 36372
rect 32088 36320 32094 36372
rect 33502 36320 33508 36372
rect 33560 36360 33566 36372
rect 34146 36360 34152 36372
rect 33560 36332 34152 36360
rect 33560 36320 33566 36332
rect 34146 36320 34152 36332
rect 34204 36360 34210 36372
rect 37366 36360 37372 36372
rect 34204 36332 37372 36360
rect 34204 36320 34210 36332
rect 37366 36320 37372 36332
rect 37424 36320 37430 36372
rect 37461 36363 37519 36369
rect 37461 36329 37473 36363
rect 37507 36360 37519 36363
rect 37642 36360 37648 36372
rect 37507 36332 37648 36360
rect 37507 36329 37519 36332
rect 37461 36323 37519 36329
rect 37642 36320 37648 36332
rect 37700 36320 37706 36372
rect 40129 36363 40187 36369
rect 40129 36329 40141 36363
rect 40175 36360 40187 36363
rect 41322 36360 41328 36372
rect 40175 36332 41328 36360
rect 40175 36329 40187 36332
rect 40129 36323 40187 36329
rect 41322 36320 41328 36332
rect 41380 36320 41386 36372
rect 48774 36360 48780 36372
rect 41800 36332 48780 36360
rect 34054 36292 34060 36304
rect 31956 36264 34060 36292
rect 34054 36252 34060 36264
rect 34112 36252 34118 36304
rect 35069 36295 35127 36301
rect 35069 36261 35081 36295
rect 35115 36292 35127 36295
rect 36538 36292 36544 36304
rect 35115 36264 36544 36292
rect 35115 36261 35127 36264
rect 35069 36255 35127 36261
rect 36538 36252 36544 36264
rect 36596 36252 36602 36304
rect 40586 36292 40592 36304
rect 37936 36264 40592 36292
rect 28350 36184 28356 36236
rect 28408 36184 28414 36236
rect 28810 36184 28816 36236
rect 28868 36224 28874 36236
rect 30466 36224 30472 36236
rect 28868 36196 30472 36224
rect 28868 36184 28874 36196
rect 30466 36184 30472 36196
rect 30524 36184 30530 36236
rect 31754 36184 31760 36236
rect 31812 36224 31818 36236
rect 32585 36227 32643 36233
rect 31812 36196 32444 36224
rect 31812 36184 31818 36196
rect 27341 36159 27399 36165
rect 27341 36125 27353 36159
rect 27387 36156 27399 36159
rect 28169 36159 28227 36165
rect 28169 36156 28181 36159
rect 27387 36128 28181 36156
rect 27387 36125 27399 36128
rect 27341 36119 27399 36125
rect 28169 36125 28181 36128
rect 28215 36125 28227 36159
rect 28169 36119 28227 36125
rect 28258 36116 28264 36168
rect 28316 36116 28322 36168
rect 32416 36165 32444 36196
rect 32585 36193 32597 36227
rect 32631 36224 32643 36227
rect 32766 36224 32772 36236
rect 32631 36196 32772 36224
rect 32631 36193 32643 36196
rect 32585 36187 32643 36193
rect 32766 36184 32772 36196
rect 32824 36184 32830 36236
rect 35526 36184 35532 36236
rect 35584 36184 35590 36236
rect 35710 36184 35716 36236
rect 35768 36184 35774 36236
rect 36446 36184 36452 36236
rect 36504 36224 36510 36236
rect 36725 36227 36783 36233
rect 36725 36224 36737 36227
rect 36504 36196 36737 36224
rect 36504 36184 36510 36196
rect 36725 36193 36737 36196
rect 36771 36193 36783 36227
rect 36725 36187 36783 36193
rect 36814 36184 36820 36236
rect 36872 36184 36878 36236
rect 37936 36233 37964 36264
rect 40586 36252 40592 36264
rect 40644 36252 40650 36304
rect 41800 36292 41828 36332
rect 48774 36320 48780 36332
rect 48832 36320 48838 36372
rect 40696 36264 41828 36292
rect 41877 36295 41935 36301
rect 37921 36227 37979 36233
rect 37921 36193 37933 36227
rect 37967 36193 37979 36227
rect 37921 36187 37979 36193
rect 38010 36184 38016 36236
rect 38068 36184 38074 36236
rect 40696 36224 40724 36264
rect 41877 36261 41889 36295
rect 41923 36292 41935 36295
rect 42794 36292 42800 36304
rect 41923 36264 42800 36292
rect 41923 36261 41935 36264
rect 41877 36255 41935 36261
rect 42794 36252 42800 36264
rect 42852 36252 42858 36304
rect 40420 36196 40724 36224
rect 40773 36227 40831 36233
rect 32401 36159 32459 36165
rect 32401 36125 32413 36159
rect 32447 36125 32459 36159
rect 32401 36119 32459 36125
rect 32493 36159 32551 36165
rect 32493 36125 32505 36159
rect 32539 36156 32551 36159
rect 32674 36156 32680 36168
rect 32539 36128 32680 36156
rect 32539 36125 32551 36128
rect 32493 36119 32551 36125
rect 32674 36116 32680 36128
rect 32732 36116 32738 36168
rect 34606 36116 34612 36168
rect 34664 36156 34670 36168
rect 36633 36159 36691 36165
rect 36633 36156 36645 36159
rect 34664 36128 36645 36156
rect 34664 36116 34670 36128
rect 36633 36125 36645 36128
rect 36679 36125 36691 36159
rect 36633 36119 36691 36125
rect 37734 36116 37740 36168
rect 37792 36156 37798 36168
rect 40420 36156 40448 36196
rect 40773 36193 40785 36227
rect 40819 36224 40831 36227
rect 41782 36224 41788 36236
rect 40819 36196 41788 36224
rect 40819 36193 40831 36196
rect 40773 36187 40831 36193
rect 41782 36184 41788 36196
rect 41840 36184 41846 36236
rect 42334 36184 42340 36236
rect 42392 36184 42398 36236
rect 42521 36227 42579 36233
rect 42521 36193 42533 36227
rect 42567 36224 42579 36227
rect 42702 36224 42708 36236
rect 42567 36196 42708 36224
rect 42567 36193 42579 36196
rect 42521 36187 42579 36193
rect 42702 36184 42708 36196
rect 42760 36184 42766 36236
rect 37792 36128 40448 36156
rect 40497 36159 40555 36165
rect 37792 36116 37798 36128
rect 40497 36125 40509 36159
rect 40543 36156 40555 36159
rect 41414 36156 41420 36168
rect 40543 36128 41420 36156
rect 40543 36125 40555 36128
rect 40497 36119 40555 36125
rect 41414 36116 41420 36128
rect 41472 36116 41478 36168
rect 20809 36091 20867 36097
rect 20809 36057 20821 36091
rect 20855 36057 20867 36091
rect 20809 36051 20867 36057
rect 20824 36020 20852 36051
rect 21818 36048 21824 36100
rect 21876 36048 21882 36100
rect 24578 36088 24584 36100
rect 22756 36060 24584 36088
rect 22756 36020 22784 36060
rect 24578 36048 24584 36060
rect 24636 36048 24642 36100
rect 26970 36048 26976 36100
rect 27028 36088 27034 36100
rect 33042 36088 33048 36100
rect 27028 36060 33048 36088
rect 27028 36048 27034 36060
rect 33042 36048 33048 36060
rect 33100 36048 33106 36100
rect 33134 36048 33140 36100
rect 33192 36088 33198 36100
rect 35437 36091 35495 36097
rect 35437 36088 35449 36091
rect 33192 36060 35449 36088
rect 33192 36048 33198 36060
rect 35437 36057 35449 36060
rect 35483 36057 35495 36091
rect 37090 36088 37096 36100
rect 35437 36051 35495 36057
rect 36188 36060 37096 36088
rect 20824 35992 22784 36020
rect 22833 36023 22891 36029
rect 22833 35989 22845 36023
rect 22879 36020 22891 36023
rect 23566 36020 23572 36032
rect 22879 35992 23572 36020
rect 22879 35989 22891 35992
rect 22833 35983 22891 35989
rect 23566 35980 23572 35992
rect 23624 36020 23630 36032
rect 23753 36023 23811 36029
rect 23753 36020 23765 36023
rect 23624 35992 23765 36020
rect 23624 35980 23630 35992
rect 23753 35989 23765 35992
rect 23799 35989 23811 36023
rect 23753 35983 23811 35989
rect 26234 35980 26240 36032
rect 26292 36020 26298 36032
rect 27801 36023 27859 36029
rect 27801 36020 27813 36023
rect 26292 35992 27813 36020
rect 26292 35980 26298 35992
rect 27801 35989 27813 35992
rect 27847 35989 27859 36023
rect 27801 35983 27859 35989
rect 34054 35980 34060 36032
rect 34112 36020 34118 36032
rect 36188 36020 36216 36060
rect 37090 36048 37096 36060
rect 37148 36088 37154 36100
rect 37550 36088 37556 36100
rect 37148 36060 37556 36088
rect 37148 36048 37154 36060
rect 37550 36048 37556 36060
rect 37608 36048 37614 36100
rect 37829 36091 37887 36097
rect 37829 36057 37841 36091
rect 37875 36088 37887 36091
rect 40126 36088 40132 36100
rect 37875 36060 40132 36088
rect 37875 36057 37887 36060
rect 37829 36051 37887 36057
rect 40126 36048 40132 36060
rect 40184 36048 40190 36100
rect 34112 35992 36216 36020
rect 36265 36023 36323 36029
rect 34112 35980 34118 35992
rect 36265 35989 36277 36023
rect 36311 36020 36323 36023
rect 36446 36020 36452 36032
rect 36311 35992 36452 36020
rect 36311 35989 36323 35992
rect 36265 35983 36323 35989
rect 36446 35980 36452 35992
rect 36504 35980 36510 36032
rect 40586 35980 40592 36032
rect 40644 35980 40650 36032
rect 42242 35980 42248 36032
rect 42300 35980 42306 36032
rect 1104 35930 49864 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 27950 35930
rect 28002 35878 28014 35930
rect 28066 35878 28078 35930
rect 28130 35878 28142 35930
rect 28194 35878 28206 35930
rect 28258 35878 37950 35930
rect 38002 35878 38014 35930
rect 38066 35878 38078 35930
rect 38130 35878 38142 35930
rect 38194 35878 38206 35930
rect 38258 35878 47950 35930
rect 48002 35878 48014 35930
rect 48066 35878 48078 35930
rect 48130 35878 48142 35930
rect 48194 35878 48206 35930
rect 48258 35878 49864 35930
rect 1104 35856 49864 35878
rect 16114 35776 16120 35828
rect 16172 35816 16178 35828
rect 21174 35816 21180 35828
rect 16172 35788 21180 35816
rect 16172 35776 16178 35788
rect 21174 35776 21180 35788
rect 21232 35776 21238 35828
rect 21269 35819 21327 35825
rect 21269 35785 21281 35819
rect 21315 35816 21327 35819
rect 21358 35816 21364 35828
rect 21315 35788 21364 35816
rect 21315 35785 21327 35788
rect 21269 35779 21327 35785
rect 21358 35776 21364 35788
rect 21416 35776 21422 35828
rect 24762 35776 24768 35828
rect 24820 35816 24826 35828
rect 24820 35788 26280 35816
rect 24820 35776 24826 35788
rect 21910 35748 21916 35760
rect 21022 35720 21916 35748
rect 21910 35708 21916 35720
rect 21968 35708 21974 35760
rect 26252 35748 26280 35788
rect 26418 35776 26424 35828
rect 26476 35816 26482 35828
rect 26694 35816 26700 35828
rect 26476 35788 26700 35816
rect 26476 35776 26482 35788
rect 26694 35776 26700 35788
rect 26752 35776 26758 35828
rect 32214 35816 32220 35828
rect 29104 35788 32220 35816
rect 28626 35748 28632 35760
rect 26174 35720 28632 35748
rect 28626 35708 28632 35720
rect 28684 35708 28690 35760
rect 24670 35640 24676 35692
rect 24728 35640 24734 35692
rect 26786 35640 26792 35692
rect 26844 35680 26850 35692
rect 29104 35689 29132 35788
rect 32214 35776 32220 35788
rect 32272 35816 32278 35828
rect 32582 35816 32588 35828
rect 32272 35788 32588 35816
rect 32272 35776 32278 35788
rect 32582 35776 32588 35788
rect 32640 35776 32646 35828
rect 33042 35776 33048 35828
rect 33100 35816 33106 35828
rect 35621 35819 35679 35825
rect 35621 35816 35633 35819
rect 33100 35788 35633 35816
rect 33100 35776 33106 35788
rect 35621 35785 35633 35788
rect 35667 35785 35679 35819
rect 35621 35779 35679 35785
rect 35989 35819 36047 35825
rect 35989 35785 36001 35819
rect 36035 35816 36047 35819
rect 38746 35816 38752 35828
rect 36035 35788 38752 35816
rect 36035 35785 36047 35788
rect 35989 35779 36047 35785
rect 38746 35776 38752 35788
rect 38804 35776 38810 35828
rect 39390 35776 39396 35828
rect 39448 35816 39454 35828
rect 39853 35819 39911 35825
rect 39448 35788 39804 35816
rect 39448 35776 39454 35788
rect 30374 35708 30380 35760
rect 30432 35708 30438 35760
rect 30742 35708 30748 35760
rect 30800 35748 30806 35760
rect 30800 35720 32628 35748
rect 30800 35708 30806 35720
rect 29089 35683 29147 35689
rect 29089 35680 29101 35683
rect 26844 35652 29101 35680
rect 26844 35640 26850 35652
rect 29089 35649 29101 35652
rect 29135 35649 29147 35683
rect 31570 35680 31576 35692
rect 29089 35643 29147 35649
rect 30576 35652 31576 35680
rect 19521 35615 19579 35621
rect 19521 35581 19533 35615
rect 19567 35612 19579 35615
rect 19797 35615 19855 35621
rect 19567 35584 19656 35612
rect 19567 35581 19579 35584
rect 19521 35575 19579 35581
rect 19628 35476 19656 35584
rect 19797 35581 19809 35615
rect 19843 35612 19855 35615
rect 23290 35612 23296 35624
rect 19843 35584 23296 35612
rect 19843 35581 19855 35584
rect 19797 35575 19855 35581
rect 23290 35572 23296 35584
rect 23348 35572 23354 35624
rect 24949 35615 25007 35621
rect 24949 35581 24961 35615
rect 24995 35612 25007 35615
rect 25038 35612 25044 35624
rect 24995 35584 25044 35612
rect 24995 35581 25007 35584
rect 24949 35575 25007 35581
rect 25038 35572 25044 35584
rect 25096 35572 25102 35624
rect 27706 35612 27712 35624
rect 26804 35584 27712 35612
rect 20530 35476 20536 35488
rect 19628 35448 20536 35476
rect 20530 35436 20536 35448
rect 20588 35436 20594 35488
rect 21174 35436 21180 35488
rect 21232 35476 21238 35488
rect 26804 35476 26832 35584
rect 27706 35572 27712 35584
rect 27764 35572 27770 35624
rect 29362 35572 29368 35624
rect 29420 35612 29426 35624
rect 30576 35612 30604 35652
rect 31570 35640 31576 35652
rect 31628 35640 31634 35692
rect 32306 35612 32312 35624
rect 29420 35584 30604 35612
rect 30852 35584 32312 35612
rect 29420 35572 29426 35584
rect 27062 35504 27068 35556
rect 27120 35544 27126 35556
rect 27120 35516 29132 35544
rect 27120 35504 27126 35516
rect 21232 35448 26832 35476
rect 21232 35436 21238 35448
rect 26878 35436 26884 35488
rect 26936 35476 26942 35488
rect 27341 35479 27399 35485
rect 27341 35476 27353 35479
rect 26936 35448 27353 35476
rect 26936 35436 26942 35448
rect 27341 35445 27353 35448
rect 27387 35445 27399 35479
rect 29104 35476 29132 35516
rect 30852 35485 30880 35584
rect 32306 35572 32312 35584
rect 32364 35572 32370 35624
rect 32600 35544 32628 35720
rect 32766 35708 32772 35760
rect 32824 35748 32830 35760
rect 33505 35751 33563 35757
rect 33505 35748 33517 35751
rect 32824 35720 33517 35748
rect 32824 35708 32830 35720
rect 33505 35717 33517 35720
rect 33551 35717 33563 35751
rect 33505 35711 33563 35717
rect 36081 35751 36139 35757
rect 36081 35717 36093 35751
rect 36127 35748 36139 35751
rect 38470 35748 38476 35760
rect 36127 35720 36400 35748
rect 36127 35717 36139 35720
rect 36081 35711 36139 35717
rect 32677 35683 32735 35689
rect 32677 35649 32689 35683
rect 32723 35680 32735 35683
rect 33873 35683 33931 35689
rect 33873 35680 33885 35683
rect 32723 35652 33885 35680
rect 32723 35649 32735 35652
rect 32677 35643 32735 35649
rect 33873 35649 33885 35652
rect 33919 35649 33931 35683
rect 33873 35643 33931 35649
rect 34793 35683 34851 35689
rect 34793 35649 34805 35683
rect 34839 35680 34851 35683
rect 35250 35680 35256 35692
rect 34839 35652 35256 35680
rect 34839 35649 34851 35652
rect 34793 35643 34851 35649
rect 35250 35640 35256 35652
rect 35308 35640 35314 35692
rect 36372 35680 36400 35720
rect 38120 35720 38476 35748
rect 36814 35680 36820 35692
rect 35912 35652 36308 35680
rect 36372 35652 36820 35680
rect 32858 35572 32864 35624
rect 32916 35572 32922 35624
rect 34698 35572 34704 35624
rect 34756 35612 34762 35624
rect 34885 35615 34943 35621
rect 34885 35612 34897 35615
rect 34756 35584 34897 35612
rect 34756 35572 34762 35584
rect 34885 35581 34897 35584
rect 34931 35581 34943 35615
rect 34885 35575 34943 35581
rect 35069 35615 35127 35621
rect 35069 35581 35081 35615
rect 35115 35612 35127 35615
rect 35912 35612 35940 35652
rect 36173 35615 36231 35621
rect 36173 35612 36185 35615
rect 35115 35584 35940 35612
rect 36004 35584 36185 35612
rect 35115 35581 35127 35584
rect 35069 35575 35127 35581
rect 36004 35544 36032 35584
rect 36173 35581 36185 35584
rect 36219 35581 36231 35615
rect 36280 35612 36308 35652
rect 36814 35640 36820 35652
rect 36872 35640 36878 35692
rect 37642 35640 37648 35692
rect 37700 35680 37706 35692
rect 38120 35689 38148 35720
rect 38470 35708 38476 35720
rect 38528 35708 38534 35760
rect 39666 35748 39672 35760
rect 39606 35720 39672 35748
rect 39666 35708 39672 35720
rect 39724 35708 39730 35760
rect 38105 35683 38163 35689
rect 38105 35680 38117 35683
rect 37700 35652 38117 35680
rect 37700 35640 37706 35652
rect 38105 35649 38117 35652
rect 38151 35649 38163 35683
rect 39776 35680 39804 35788
rect 39853 35785 39865 35819
rect 39899 35816 39911 35819
rect 39942 35816 39948 35828
rect 39899 35788 39948 35816
rect 39899 35785 39911 35788
rect 39853 35779 39911 35785
rect 39942 35776 39948 35788
rect 40000 35776 40006 35828
rect 40126 35776 40132 35828
rect 40184 35816 40190 35828
rect 40770 35816 40776 35828
rect 40184 35788 40776 35816
rect 40184 35776 40190 35788
rect 40770 35776 40776 35788
rect 40828 35816 40834 35828
rect 49050 35816 49056 35828
rect 40828 35788 49056 35816
rect 40828 35776 40834 35788
rect 49050 35776 49056 35788
rect 49108 35776 49114 35828
rect 40218 35708 40224 35760
rect 40276 35748 40282 35760
rect 40276 35720 40816 35748
rect 40276 35708 40282 35720
rect 40681 35683 40739 35689
rect 40681 35680 40693 35683
rect 39776 35652 40693 35680
rect 38105 35643 38163 35649
rect 40681 35649 40693 35652
rect 40727 35649 40739 35683
rect 40788 35680 40816 35720
rect 41874 35708 41880 35760
rect 41932 35748 41938 35760
rect 42889 35751 42947 35757
rect 42889 35748 42901 35751
rect 41932 35720 42901 35748
rect 41932 35708 41938 35720
rect 42889 35717 42901 35720
rect 42935 35748 42947 35751
rect 43162 35748 43168 35760
rect 42935 35720 43168 35748
rect 42935 35717 42947 35720
rect 42889 35711 42947 35717
rect 43162 35708 43168 35720
rect 43220 35708 43226 35760
rect 43438 35708 43444 35760
rect 43496 35708 43502 35760
rect 40788 35652 40908 35680
rect 40681 35643 40739 35649
rect 37826 35612 37832 35624
rect 36280 35584 37832 35612
rect 36173 35575 36231 35581
rect 37826 35572 37832 35584
rect 37884 35572 37890 35624
rect 38378 35572 38384 35624
rect 38436 35612 38442 35624
rect 39758 35612 39764 35624
rect 38436 35584 39764 35612
rect 38436 35572 38442 35584
rect 39758 35572 39764 35584
rect 39816 35572 39822 35624
rect 40402 35572 40408 35624
rect 40460 35612 40466 35624
rect 40880 35621 40908 35652
rect 40773 35615 40831 35621
rect 40773 35612 40785 35615
rect 40460 35584 40785 35612
rect 40460 35572 40466 35584
rect 40773 35581 40785 35584
rect 40819 35581 40831 35615
rect 40773 35575 40831 35581
rect 40865 35615 40923 35621
rect 40865 35581 40877 35615
rect 40911 35612 40923 35615
rect 41892 35612 41920 35708
rect 42610 35640 42616 35692
rect 42668 35640 42674 35692
rect 49326 35640 49332 35692
rect 49384 35640 49390 35692
rect 40911 35584 41920 35612
rect 40911 35581 40923 35584
rect 40865 35575 40923 35581
rect 42334 35572 42340 35624
rect 42392 35612 42398 35624
rect 42392 35584 43944 35612
rect 42392 35572 42398 35584
rect 32600 35516 36032 35544
rect 40313 35547 40371 35553
rect 40313 35513 40325 35547
rect 40359 35544 40371 35547
rect 42242 35544 42248 35556
rect 40359 35516 42248 35544
rect 40359 35513 40371 35516
rect 40313 35507 40371 35513
rect 42242 35504 42248 35516
rect 42300 35504 42306 35556
rect 43916 35544 43944 35584
rect 49145 35547 49203 35553
rect 49145 35544 49157 35547
rect 43916 35516 49157 35544
rect 49145 35513 49157 35516
rect 49191 35513 49203 35547
rect 49145 35507 49203 35513
rect 30837 35479 30895 35485
rect 30837 35476 30849 35479
rect 29104 35448 30849 35476
rect 27341 35439 27399 35445
rect 30837 35445 30849 35448
rect 30883 35445 30895 35479
rect 30837 35439 30895 35445
rect 31754 35436 31760 35488
rect 31812 35436 31818 35488
rect 32309 35479 32367 35485
rect 32309 35445 32321 35479
rect 32355 35476 32367 35479
rect 33134 35476 33140 35488
rect 32355 35448 33140 35476
rect 32355 35445 32367 35448
rect 32309 35439 32367 35445
rect 33134 35436 33140 35448
rect 33192 35436 33198 35488
rect 34425 35479 34483 35485
rect 34425 35445 34437 35479
rect 34471 35476 34483 35479
rect 38930 35476 38936 35488
rect 34471 35448 38936 35476
rect 34471 35445 34483 35448
rect 34425 35439 34483 35445
rect 38930 35436 38936 35448
rect 38988 35436 38994 35488
rect 42702 35436 42708 35488
rect 42760 35476 42766 35488
rect 44361 35479 44419 35485
rect 44361 35476 44373 35479
rect 42760 35448 44373 35476
rect 42760 35436 42766 35448
rect 44361 35445 44373 35448
rect 44407 35445 44419 35479
rect 44361 35439 44419 35445
rect 1104 35386 49864 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 32950 35386
rect 33002 35334 33014 35386
rect 33066 35334 33078 35386
rect 33130 35334 33142 35386
rect 33194 35334 33206 35386
rect 33258 35334 42950 35386
rect 43002 35334 43014 35386
rect 43066 35334 43078 35386
rect 43130 35334 43142 35386
rect 43194 35334 43206 35386
rect 43258 35334 49864 35386
rect 1104 35312 49864 35334
rect 22002 35232 22008 35284
rect 22060 35272 22066 35284
rect 24581 35275 24639 35281
rect 24581 35272 24593 35275
rect 22060 35244 24593 35272
rect 22060 35232 22066 35244
rect 24581 35241 24593 35244
rect 24627 35241 24639 35275
rect 24581 35235 24639 35241
rect 25958 35232 25964 35284
rect 26016 35272 26022 35284
rect 26053 35275 26111 35281
rect 26053 35272 26065 35275
rect 26016 35244 26065 35272
rect 26016 35232 26022 35244
rect 26053 35241 26065 35244
rect 26099 35241 26111 35275
rect 26878 35272 26884 35284
rect 26053 35235 26111 35241
rect 26515 35244 26884 35272
rect 26515 35204 26543 35244
rect 26878 35232 26884 35244
rect 26936 35232 26942 35284
rect 27522 35232 27528 35284
rect 27580 35272 27586 35284
rect 28997 35275 29055 35281
rect 28997 35272 29009 35275
rect 27580 35244 29009 35272
rect 27580 35232 27586 35244
rect 28997 35241 29009 35244
rect 29043 35241 29055 35275
rect 28997 35235 29055 35241
rect 29178 35232 29184 35284
rect 29236 35272 29242 35284
rect 30742 35272 30748 35284
rect 29236 35244 30748 35272
rect 29236 35232 29242 35244
rect 30742 35232 30748 35244
rect 30800 35232 30806 35284
rect 33870 35232 33876 35284
rect 33928 35272 33934 35284
rect 33965 35275 34023 35281
rect 33965 35272 33977 35275
rect 33928 35244 33977 35272
rect 33928 35232 33934 35244
rect 33965 35241 33977 35244
rect 34011 35241 34023 35275
rect 33965 35235 34023 35241
rect 35066 35232 35072 35284
rect 35124 35272 35130 35284
rect 37369 35275 37427 35281
rect 37369 35272 37381 35275
rect 35124 35244 37381 35272
rect 35124 35232 35130 35244
rect 37369 35241 37381 35244
rect 37415 35241 37427 35275
rect 37369 35235 37427 35241
rect 38746 35232 38752 35284
rect 38804 35272 38810 35284
rect 49142 35272 49148 35284
rect 38804 35244 49148 35272
rect 38804 35232 38810 35244
rect 49142 35232 49148 35244
rect 49200 35232 49206 35284
rect 27062 35204 27068 35216
rect 26436 35176 26543 35204
rect 26712 35176 27068 35204
rect 22005 35139 22063 35145
rect 22005 35105 22017 35139
rect 22051 35136 22063 35139
rect 22094 35136 22100 35148
rect 22051 35108 22100 35136
rect 22051 35105 22063 35108
rect 22005 35099 22063 35105
rect 22094 35096 22100 35108
rect 22152 35136 22158 35148
rect 22152 35108 23244 35136
rect 22152 35096 22158 35108
rect 20530 35028 20536 35080
rect 20588 35068 20594 35080
rect 21726 35068 21732 35080
rect 20588 35040 21732 35068
rect 20588 35028 20594 35040
rect 21726 35028 21732 35040
rect 21784 35028 21790 35080
rect 23216 35068 23244 35108
rect 23290 35096 23296 35148
rect 23348 35136 23354 35148
rect 25133 35139 25191 35145
rect 25133 35136 25145 35139
rect 23348 35108 25145 35136
rect 23348 35096 23354 35108
rect 25133 35105 25145 35108
rect 25179 35105 25191 35139
rect 25133 35099 25191 35105
rect 25041 35071 25099 35077
rect 23216 35040 24992 35068
rect 24762 35000 24768 35012
rect 23230 34972 24768 35000
rect 21910 34892 21916 34944
rect 21968 34932 21974 34944
rect 23308 34932 23336 34972
rect 24762 34960 24768 34972
rect 24820 34960 24826 35012
rect 24964 35000 24992 35040
rect 25041 35037 25053 35071
rect 25087 35068 25099 35071
rect 26234 35068 26240 35080
rect 25087 35040 26240 35068
rect 25087 35037 25099 35040
rect 25041 35031 25099 35037
rect 26234 35028 26240 35040
rect 26292 35028 26298 35080
rect 26436 35077 26464 35176
rect 26712 35145 26740 35176
rect 27062 35164 27068 35176
rect 27120 35164 27126 35216
rect 28902 35164 28908 35216
rect 28960 35204 28966 35216
rect 29733 35207 29791 35213
rect 29733 35204 29745 35207
rect 28960 35176 29745 35204
rect 28960 35164 28966 35176
rect 29733 35173 29745 35176
rect 29779 35173 29791 35207
rect 29733 35167 29791 35173
rect 32140 35176 32352 35204
rect 26697 35139 26755 35145
rect 26697 35105 26709 35139
rect 26743 35105 26755 35139
rect 26697 35099 26755 35105
rect 26786 35096 26792 35148
rect 26844 35136 26850 35148
rect 27249 35139 27307 35145
rect 27249 35136 27261 35139
rect 26844 35108 27261 35136
rect 26844 35096 26850 35108
rect 27249 35105 27261 35108
rect 27295 35105 27307 35139
rect 27249 35099 27307 35105
rect 27525 35139 27583 35145
rect 27525 35105 27537 35139
rect 27571 35136 27583 35139
rect 30006 35136 30012 35148
rect 27571 35108 30012 35136
rect 27571 35105 27583 35108
rect 27525 35099 27583 35105
rect 30006 35096 30012 35108
rect 30064 35096 30070 35148
rect 30282 35096 30288 35148
rect 30340 35096 30346 35148
rect 31202 35096 31208 35148
rect 31260 35136 31266 35148
rect 31481 35139 31539 35145
rect 31481 35136 31493 35139
rect 31260 35108 31493 35136
rect 31260 35096 31266 35108
rect 31481 35105 31493 35108
rect 31527 35105 31539 35139
rect 31481 35099 31539 35105
rect 31662 35096 31668 35148
rect 31720 35096 31726 35148
rect 26421 35071 26479 35077
rect 26421 35037 26433 35071
rect 26467 35037 26479 35071
rect 26421 35031 26479 35037
rect 28626 35028 28632 35080
rect 28684 35068 28690 35080
rect 28810 35068 28816 35080
rect 28684 35040 28816 35068
rect 28684 35028 28690 35040
rect 28810 35028 28816 35040
rect 28868 35028 28874 35080
rect 30098 35028 30104 35080
rect 30156 35028 30162 35080
rect 31386 35028 31392 35080
rect 31444 35028 31450 35080
rect 25590 35000 25596 35012
rect 24964 34972 25596 35000
rect 25590 34960 25596 34972
rect 25648 34960 25654 35012
rect 26326 34960 26332 35012
rect 26384 35000 26390 35012
rect 26513 35003 26571 35009
rect 26513 35000 26525 35003
rect 26384 34972 26525 35000
rect 26384 34960 26390 34972
rect 26513 34969 26525 34972
rect 26559 34969 26571 35003
rect 26513 34963 26571 34969
rect 26602 34960 26608 35012
rect 26660 35000 26666 35012
rect 26660 34972 27936 35000
rect 26660 34960 26666 34972
rect 21968 34904 23336 34932
rect 23477 34935 23535 34941
rect 21968 34892 21974 34904
rect 23477 34901 23489 34935
rect 23523 34932 23535 34935
rect 24578 34932 24584 34944
rect 23523 34904 24584 34932
rect 23523 34901 23535 34904
rect 23477 34895 23535 34901
rect 24578 34892 24584 34904
rect 24636 34892 24642 34944
rect 24949 34935 25007 34941
rect 24949 34901 24961 34935
rect 24995 34932 25007 34935
rect 27798 34932 27804 34944
rect 24995 34904 27804 34932
rect 24995 34901 25007 34904
rect 24949 34895 25007 34901
rect 27798 34892 27804 34904
rect 27856 34892 27862 34944
rect 27908 34932 27936 34972
rect 30558 34960 30564 35012
rect 30616 35000 30622 35012
rect 32140 35000 32168 35176
rect 32214 35096 32220 35148
rect 32272 35096 32278 35148
rect 32324 35136 32352 35176
rect 34624 35176 36768 35204
rect 32493 35139 32551 35145
rect 32493 35136 32505 35139
rect 32324 35108 32505 35136
rect 32493 35105 32505 35108
rect 32539 35136 32551 35139
rect 34624 35136 34652 35176
rect 36740 35148 36768 35176
rect 36814 35164 36820 35216
rect 36872 35204 36878 35216
rect 39022 35204 39028 35216
rect 36872 35176 39028 35204
rect 36872 35164 36878 35176
rect 39022 35164 39028 35176
rect 39080 35164 39086 35216
rect 32539 35108 34652 35136
rect 32539 35105 32551 35108
rect 32493 35099 32551 35105
rect 36630 35096 36636 35148
rect 36688 35096 36694 35148
rect 36722 35096 36728 35148
rect 36780 35136 36786 35148
rect 37921 35139 37979 35145
rect 37921 35136 37933 35139
rect 36780 35108 37933 35136
rect 36780 35096 36786 35108
rect 37921 35105 37933 35108
rect 37967 35105 37979 35139
rect 37921 35099 37979 35105
rect 38654 35096 38660 35148
rect 38712 35136 38718 35148
rect 39117 35139 39175 35145
rect 39117 35136 39129 35139
rect 38712 35108 39129 35136
rect 38712 35096 38718 35108
rect 39117 35105 39129 35108
rect 39163 35105 39175 35139
rect 39117 35099 39175 35105
rect 42610 35096 42616 35148
rect 42668 35136 42674 35148
rect 42705 35139 42763 35145
rect 42705 35136 42717 35139
rect 42668 35108 42717 35136
rect 42668 35096 42674 35108
rect 42705 35105 42717 35108
rect 42751 35105 42763 35139
rect 42705 35099 42763 35105
rect 43530 35096 43536 35148
rect 43588 35136 43594 35148
rect 44453 35139 44511 35145
rect 44453 35136 44465 35139
rect 43588 35108 44465 35136
rect 43588 35096 43594 35108
rect 44453 35105 44465 35108
rect 44499 35105 44511 35139
rect 44453 35099 44511 35105
rect 34974 35068 34980 35080
rect 33626 35054 34980 35068
rect 30616 34972 32168 35000
rect 33612 35040 34980 35054
rect 30616 34960 30622 34972
rect 30193 34935 30251 34941
rect 30193 34932 30205 34935
rect 27908 34904 30205 34932
rect 30193 34901 30205 34904
rect 30239 34901 30251 34935
rect 30193 34895 30251 34901
rect 31018 34892 31024 34944
rect 31076 34892 31082 34944
rect 31202 34892 31208 34944
rect 31260 34932 31266 34944
rect 32766 34932 32772 34944
rect 31260 34904 32772 34932
rect 31260 34892 31266 34904
rect 32766 34892 32772 34904
rect 32824 34892 32830 34944
rect 33410 34892 33416 34944
rect 33468 34932 33474 34944
rect 33612 34932 33640 35040
rect 34974 35028 34980 35040
rect 35032 35068 35038 35080
rect 35802 35068 35808 35080
rect 35032 35040 35808 35068
rect 35032 35028 35038 35040
rect 35802 35028 35808 35040
rect 35860 35028 35866 35080
rect 36449 35071 36507 35077
rect 36449 35037 36461 35071
rect 36495 35068 36507 35071
rect 37458 35068 37464 35080
rect 36495 35040 37464 35068
rect 36495 35037 36507 35040
rect 36449 35031 36507 35037
rect 37458 35028 37464 35040
rect 37516 35028 37522 35080
rect 37829 35071 37887 35077
rect 37829 35037 37841 35071
rect 37875 35068 37887 35071
rect 39850 35068 39856 35080
rect 37875 35040 39856 35068
rect 37875 35037 37887 35040
rect 37829 35031 37887 35037
rect 39850 35028 39856 35040
rect 39908 35028 39914 35080
rect 41690 35028 41696 35080
rect 41748 35068 41754 35080
rect 41969 35071 42027 35077
rect 41969 35068 41981 35071
rect 41748 35040 41981 35068
rect 41748 35028 41754 35040
rect 41969 35037 41981 35040
rect 42015 35037 42027 35071
rect 48406 35068 48412 35080
rect 41969 35031 42027 35037
rect 44468 35040 48412 35068
rect 34514 34960 34520 35012
rect 34572 35000 34578 35012
rect 37737 35003 37795 35009
rect 34572 34972 36492 35000
rect 34572 34960 34578 34972
rect 33468 34904 33640 34932
rect 35989 34935 36047 34941
rect 33468 34892 33474 34904
rect 35989 34901 36001 34935
rect 36035 34932 36047 34935
rect 36170 34932 36176 34944
rect 36035 34904 36176 34932
rect 36035 34901 36047 34904
rect 35989 34895 36047 34901
rect 36170 34892 36176 34904
rect 36228 34892 36234 34944
rect 36354 34892 36360 34944
rect 36412 34892 36418 34944
rect 36464 34932 36492 34972
rect 37737 34969 37749 35003
rect 37783 35000 37795 35003
rect 42426 35000 42432 35012
rect 37783 34972 42432 35000
rect 37783 34969 37795 34972
rect 37737 34963 37795 34969
rect 42426 34960 42432 34972
rect 42484 34960 42490 35012
rect 42702 34960 42708 35012
rect 42760 35000 42766 35012
rect 42981 35003 43039 35009
rect 42981 35000 42993 35003
rect 42760 34972 42993 35000
rect 42760 34960 42766 34972
rect 42981 34969 42993 34972
rect 43027 34969 43039 35003
rect 42981 34963 43039 34969
rect 43438 34960 43444 35012
rect 43496 34960 43502 35012
rect 38565 34935 38623 34941
rect 38565 34932 38577 34935
rect 36464 34904 38577 34932
rect 38565 34901 38577 34904
rect 38611 34901 38623 34935
rect 38565 34895 38623 34901
rect 38930 34892 38936 34944
rect 38988 34892 38994 34944
rect 39025 34935 39083 34941
rect 39025 34901 39037 34935
rect 39071 34932 39083 34935
rect 40494 34932 40500 34944
rect 39071 34904 40500 34932
rect 39071 34901 39083 34904
rect 39025 34895 39083 34901
rect 40494 34892 40500 34904
rect 40552 34892 40558 34944
rect 40862 34892 40868 34944
rect 40920 34932 40926 34944
rect 44468 34932 44496 35040
rect 48406 35028 48412 35040
rect 48464 35028 48470 35080
rect 49326 35028 49332 35080
rect 49384 35028 49390 35080
rect 40920 34904 44496 34932
rect 40920 34892 40926 34904
rect 44542 34892 44548 34944
rect 44600 34932 44606 34944
rect 46934 34932 46940 34944
rect 44600 34904 46940 34932
rect 44600 34892 44606 34904
rect 46934 34892 46940 34904
rect 46992 34892 46998 34944
rect 49050 34892 49056 34944
rect 49108 34932 49114 34944
rect 49145 34935 49203 34941
rect 49145 34932 49157 34935
rect 49108 34904 49157 34932
rect 49108 34892 49114 34904
rect 49145 34901 49157 34904
rect 49191 34901 49203 34935
rect 49145 34895 49203 34901
rect 1104 34842 49864 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 27950 34842
rect 28002 34790 28014 34842
rect 28066 34790 28078 34842
rect 28130 34790 28142 34842
rect 28194 34790 28206 34842
rect 28258 34790 37950 34842
rect 38002 34790 38014 34842
rect 38066 34790 38078 34842
rect 38130 34790 38142 34842
rect 38194 34790 38206 34842
rect 38258 34790 47950 34842
rect 48002 34790 48014 34842
rect 48066 34790 48078 34842
rect 48130 34790 48142 34842
rect 48194 34790 48206 34842
rect 48258 34790 49864 34842
rect 1104 34768 49864 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 7834 34728 7840 34740
rect 1627 34700 7840 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 7834 34688 7840 34700
rect 7892 34688 7898 34740
rect 24854 34688 24860 34740
rect 24912 34728 24918 34740
rect 25317 34731 25375 34737
rect 25317 34728 25329 34731
rect 24912 34700 25329 34728
rect 24912 34688 24918 34700
rect 25317 34697 25329 34700
rect 25363 34697 25375 34731
rect 25317 34691 25375 34697
rect 25590 34688 25596 34740
rect 25648 34728 25654 34740
rect 28258 34728 28264 34740
rect 25648 34700 28264 34728
rect 25648 34688 25654 34700
rect 28258 34688 28264 34700
rect 28316 34728 28322 34740
rect 29178 34728 29184 34740
rect 28316 34700 29184 34728
rect 28316 34688 28322 34700
rect 29178 34688 29184 34700
rect 29236 34688 29242 34740
rect 31021 34731 31079 34737
rect 31021 34728 31033 34731
rect 30484 34700 31033 34728
rect 24762 34660 24768 34672
rect 24518 34632 24768 34660
rect 24762 34620 24768 34632
rect 24820 34620 24826 34672
rect 25777 34663 25835 34669
rect 25777 34629 25789 34663
rect 25823 34660 25835 34663
rect 28626 34660 28632 34672
rect 25823 34632 28632 34660
rect 25823 34629 25835 34632
rect 25777 34623 25835 34629
rect 28626 34620 28632 34632
rect 28684 34620 28690 34672
rect 30374 34660 30380 34672
rect 29762 34632 30380 34660
rect 30374 34620 30380 34632
rect 30432 34620 30438 34672
rect 1762 34552 1768 34604
rect 1820 34552 1826 34604
rect 22646 34552 22652 34604
rect 22704 34592 22710 34604
rect 23017 34595 23075 34601
rect 23017 34592 23029 34595
rect 22704 34564 23029 34592
rect 22704 34552 22710 34564
rect 23017 34561 23029 34564
rect 23063 34561 23075 34595
rect 23017 34555 23075 34561
rect 25682 34552 25688 34604
rect 25740 34552 25746 34604
rect 26786 34552 26792 34604
rect 26844 34592 26850 34604
rect 28261 34595 28319 34601
rect 28261 34592 28273 34595
rect 26844 34564 28273 34592
rect 26844 34552 26850 34564
rect 28261 34561 28273 34564
rect 28307 34561 28319 34595
rect 28261 34555 28319 34561
rect 29914 34552 29920 34604
rect 29972 34592 29978 34604
rect 30484 34592 30512 34700
rect 31021 34697 31033 34700
rect 31067 34697 31079 34731
rect 31021 34691 31079 34697
rect 31294 34688 31300 34740
rect 31352 34728 31358 34740
rect 31389 34731 31447 34737
rect 31389 34728 31401 34731
rect 31352 34700 31401 34728
rect 31352 34688 31358 34700
rect 31389 34697 31401 34700
rect 31435 34697 31447 34731
rect 31389 34691 31447 34697
rect 31754 34688 31760 34740
rect 31812 34728 31818 34740
rect 32677 34731 32735 34737
rect 32677 34728 32689 34731
rect 31812 34700 32689 34728
rect 31812 34688 31818 34700
rect 32677 34697 32689 34700
rect 32723 34697 32735 34731
rect 32677 34691 32735 34697
rect 32766 34688 32772 34740
rect 32824 34728 32830 34740
rect 33505 34731 33563 34737
rect 33505 34728 33517 34731
rect 32824 34700 33517 34728
rect 32824 34688 32830 34700
rect 33505 34697 33517 34700
rect 33551 34697 33563 34731
rect 35805 34731 35863 34737
rect 35805 34728 35817 34731
rect 33505 34691 33563 34697
rect 33612 34700 35817 34728
rect 33612 34660 33640 34700
rect 35805 34697 35817 34700
rect 35851 34697 35863 34731
rect 35805 34691 35863 34697
rect 38933 34731 38991 34737
rect 38933 34697 38945 34731
rect 38979 34697 38991 34731
rect 38933 34691 38991 34697
rect 39393 34731 39451 34737
rect 39393 34697 39405 34731
rect 39439 34728 39451 34731
rect 40034 34728 40040 34740
rect 39439 34700 40040 34728
rect 39439 34697 39451 34700
rect 39393 34691 39451 34697
rect 34606 34660 34612 34672
rect 32692 34632 33640 34660
rect 34072 34632 34612 34660
rect 32692 34604 32720 34632
rect 29972 34564 30512 34592
rect 31481 34595 31539 34601
rect 29972 34552 29978 34564
rect 31481 34561 31493 34595
rect 31527 34592 31539 34595
rect 32582 34592 32588 34604
rect 31527 34564 32588 34592
rect 31527 34561 31539 34564
rect 31481 34555 31539 34561
rect 32582 34552 32588 34564
rect 32640 34552 32646 34604
rect 32674 34552 32680 34604
rect 32732 34552 32738 34604
rect 34072 34592 34100 34632
rect 34606 34620 34612 34632
rect 34664 34620 34670 34672
rect 34974 34620 34980 34672
rect 35032 34620 35038 34672
rect 37642 34660 37648 34672
rect 37016 34632 37648 34660
rect 32784 34564 34100 34592
rect 24765 34527 24823 34533
rect 24765 34493 24777 34527
rect 24811 34524 24823 34527
rect 24854 34524 24860 34536
rect 24811 34496 24860 34524
rect 24811 34493 24823 34496
rect 24765 34487 24823 34493
rect 24854 34484 24860 34496
rect 24912 34484 24918 34536
rect 25961 34527 26019 34533
rect 25961 34493 25973 34527
rect 26007 34524 26019 34527
rect 26418 34524 26424 34536
rect 26007 34496 26424 34524
rect 26007 34493 26019 34496
rect 25961 34487 26019 34493
rect 26418 34484 26424 34496
rect 26476 34484 26482 34536
rect 31573 34527 31631 34533
rect 28368 34496 29592 34524
rect 24302 34416 24308 34468
rect 24360 34456 24366 34468
rect 28368 34456 28396 34496
rect 24360 34428 28396 34456
rect 29564 34456 29592 34496
rect 31573 34493 31585 34527
rect 31619 34493 31631 34527
rect 32784 34524 32812 34564
rect 31573 34487 31631 34493
rect 32324 34496 32812 34524
rect 32953 34527 33011 34533
rect 30926 34456 30932 34468
rect 29564 34428 30932 34456
rect 24360 34416 24366 34428
rect 30926 34416 30932 34428
rect 30984 34456 30990 34468
rect 31588 34456 31616 34487
rect 32324 34465 32352 34496
rect 32953 34493 32965 34527
rect 32999 34493 33011 34527
rect 32953 34487 33011 34493
rect 30984 34428 31616 34456
rect 32309 34459 32367 34465
rect 30984 34416 30990 34428
rect 32309 34425 32321 34459
rect 32355 34425 32367 34459
rect 32968 34456 32996 34487
rect 33962 34484 33968 34536
rect 34020 34524 34026 34536
rect 34057 34527 34115 34533
rect 34057 34524 34069 34527
rect 34020 34496 34069 34524
rect 34020 34484 34026 34496
rect 34057 34493 34069 34496
rect 34103 34524 34115 34527
rect 37016 34524 37044 34632
rect 37642 34620 37648 34632
rect 37700 34620 37706 34672
rect 38948 34660 38976 34691
rect 40034 34688 40040 34700
rect 40092 34688 40098 34740
rect 40494 34688 40500 34740
rect 40552 34688 40558 34740
rect 40589 34731 40647 34737
rect 40589 34697 40601 34731
rect 40635 34728 40647 34731
rect 40954 34728 40960 34740
rect 40635 34700 40960 34728
rect 40635 34697 40647 34700
rect 40589 34691 40647 34697
rect 40954 34688 40960 34700
rect 41012 34688 41018 34740
rect 41325 34731 41383 34737
rect 41325 34697 41337 34731
rect 41371 34697 41383 34731
rect 41325 34691 41383 34697
rect 41230 34660 41236 34672
rect 38948 34632 41236 34660
rect 41230 34620 41236 34632
rect 41288 34620 41294 34672
rect 41340 34660 41368 34691
rect 41690 34688 41696 34740
rect 41748 34688 41754 34740
rect 42794 34688 42800 34740
rect 42852 34728 42858 34740
rect 43441 34731 43499 34737
rect 43441 34728 43453 34731
rect 42852 34700 43453 34728
rect 42852 34688 42858 34700
rect 43441 34697 43453 34700
rect 43487 34697 43499 34731
rect 43441 34691 43499 34697
rect 49142 34688 49148 34740
rect 49200 34688 49206 34740
rect 43349 34663 43407 34669
rect 43349 34660 43361 34663
rect 41340 34632 43361 34660
rect 43349 34629 43361 34632
rect 43395 34629 43407 34663
rect 43349 34623 43407 34629
rect 37274 34552 37280 34604
rect 37332 34592 37338 34604
rect 39301 34595 39359 34601
rect 39301 34592 39313 34595
rect 37332 34564 39313 34592
rect 37332 34552 37338 34564
rect 39301 34561 39313 34564
rect 39347 34561 39359 34595
rect 39301 34555 39359 34561
rect 39408 34564 40172 34592
rect 34103 34496 37044 34524
rect 34103 34493 34115 34496
rect 34057 34487 34115 34493
rect 37090 34484 37096 34536
rect 37148 34524 37154 34536
rect 39408 34524 39436 34564
rect 37148 34496 39436 34524
rect 39577 34527 39635 34533
rect 37148 34484 37154 34496
rect 39577 34493 39589 34527
rect 39623 34524 39635 34527
rect 39942 34524 39948 34536
rect 39623 34496 39948 34524
rect 39623 34493 39635 34496
rect 39577 34487 39635 34493
rect 39942 34484 39948 34496
rect 40000 34484 40006 34536
rect 33778 34456 33784 34468
rect 32968 34428 33784 34456
rect 32309 34419 32367 34425
rect 33778 34416 33784 34428
rect 33836 34416 33842 34468
rect 37734 34416 37740 34468
rect 37792 34456 37798 34468
rect 38562 34456 38568 34468
rect 37792 34428 38568 34456
rect 37792 34416 37798 34428
rect 38562 34416 38568 34428
rect 38620 34416 38626 34468
rect 40144 34465 40172 34564
rect 40494 34552 40500 34604
rect 40552 34592 40558 34604
rect 44542 34592 44548 34604
rect 40552 34564 44548 34592
rect 40552 34552 40558 34564
rect 44542 34552 44548 34564
rect 44600 34552 44606 34604
rect 49326 34552 49332 34604
rect 49384 34552 49390 34604
rect 40773 34527 40831 34533
rect 40773 34493 40785 34527
rect 40819 34493 40831 34527
rect 40773 34487 40831 34493
rect 40129 34459 40187 34465
rect 40129 34425 40141 34459
rect 40175 34425 40187 34459
rect 40788 34456 40816 34487
rect 40862 34484 40868 34536
rect 40920 34524 40926 34536
rect 41785 34527 41843 34533
rect 41785 34524 41797 34527
rect 40920 34496 41797 34524
rect 40920 34484 40926 34496
rect 41785 34493 41797 34496
rect 41831 34493 41843 34527
rect 41785 34487 41843 34493
rect 41969 34527 42027 34533
rect 41969 34493 41981 34527
rect 42015 34524 42027 34527
rect 42702 34524 42708 34536
rect 42015 34496 42708 34524
rect 42015 34493 42027 34496
rect 41969 34487 42027 34493
rect 42702 34484 42708 34496
rect 42760 34484 42766 34536
rect 43530 34484 43536 34536
rect 43588 34484 43594 34536
rect 44266 34524 44272 34536
rect 43640 34496 44272 34524
rect 41598 34456 41604 34468
rect 40788 34428 41604 34456
rect 40129 34419 40187 34425
rect 41598 34416 41604 34428
rect 41656 34416 41662 34468
rect 42981 34459 43039 34465
rect 42981 34425 42993 34459
rect 43027 34456 43039 34459
rect 43640 34456 43668 34496
rect 44266 34484 44272 34496
rect 44324 34484 44330 34536
rect 43027 34428 43668 34456
rect 43027 34425 43039 34428
rect 42981 34419 43039 34425
rect 22370 34348 22376 34400
rect 22428 34388 22434 34400
rect 23274 34391 23332 34397
rect 23274 34388 23286 34391
rect 22428 34360 23286 34388
rect 22428 34348 22434 34360
rect 23274 34357 23286 34360
rect 23320 34357 23332 34391
rect 23274 34351 23332 34357
rect 27706 34348 27712 34400
rect 27764 34388 27770 34400
rect 28518 34391 28576 34397
rect 28518 34388 28530 34391
rect 27764 34360 28530 34388
rect 27764 34348 27770 34360
rect 28518 34357 28530 34360
rect 28564 34388 28576 34391
rect 29270 34388 29276 34400
rect 28564 34360 29276 34388
rect 28564 34357 28576 34360
rect 28518 34351 28576 34357
rect 29270 34348 29276 34360
rect 29328 34348 29334 34400
rect 30006 34348 30012 34400
rect 30064 34388 30070 34400
rect 31478 34388 31484 34400
rect 30064 34360 31484 34388
rect 30064 34348 30070 34360
rect 31478 34348 31484 34360
rect 31536 34348 31542 34400
rect 34320 34391 34378 34397
rect 34320 34357 34332 34391
rect 34366 34388 34378 34391
rect 39758 34388 39764 34400
rect 34366 34360 39764 34388
rect 34366 34357 34378 34360
rect 34320 34351 34378 34357
rect 39758 34348 39764 34360
rect 39816 34348 39822 34400
rect 1104 34298 49864 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 32950 34298
rect 33002 34246 33014 34298
rect 33066 34246 33078 34298
rect 33130 34246 33142 34298
rect 33194 34246 33206 34298
rect 33258 34246 42950 34298
rect 43002 34246 43014 34298
rect 43066 34246 43078 34298
rect 43130 34246 43142 34298
rect 43194 34246 43206 34298
rect 43258 34246 49864 34298
rect 1104 34224 49864 34246
rect 20990 34144 20996 34196
rect 21048 34184 21054 34196
rect 23293 34187 23351 34193
rect 23293 34184 23305 34187
rect 21048 34156 23305 34184
rect 21048 34144 21054 34156
rect 23293 34153 23305 34156
rect 23339 34153 23351 34187
rect 23293 34147 23351 34153
rect 26500 34187 26558 34193
rect 26500 34153 26512 34187
rect 26546 34184 26558 34187
rect 27522 34184 27528 34196
rect 26546 34156 27528 34184
rect 26546 34153 26558 34156
rect 26500 34147 26558 34153
rect 27522 34144 27528 34156
rect 27580 34144 27586 34196
rect 29086 34144 29092 34196
rect 29144 34184 29150 34196
rect 35986 34184 35992 34196
rect 29144 34156 35992 34184
rect 29144 34144 29150 34156
rect 35986 34144 35992 34156
rect 36044 34144 36050 34196
rect 36265 34187 36323 34193
rect 36265 34153 36277 34187
rect 36311 34184 36323 34187
rect 40586 34184 40592 34196
rect 36311 34156 40592 34184
rect 36311 34153 36323 34156
rect 36265 34147 36323 34153
rect 40586 34144 40592 34156
rect 40644 34144 40650 34196
rect 48958 34184 48964 34196
rect 41386 34156 48964 34184
rect 22554 34076 22560 34128
rect 22612 34116 22618 34128
rect 24581 34119 24639 34125
rect 24581 34116 24593 34119
rect 22612 34088 24593 34116
rect 22612 34076 22618 34088
rect 24581 34085 24593 34088
rect 24627 34085 24639 34119
rect 24581 34079 24639 34085
rect 30745 34119 30803 34125
rect 30745 34085 30757 34119
rect 30791 34116 30803 34119
rect 36354 34116 36360 34128
rect 30791 34088 36360 34116
rect 30791 34085 30803 34088
rect 30745 34079 30803 34085
rect 36354 34076 36360 34088
rect 36412 34076 36418 34128
rect 37366 34116 37372 34128
rect 36740 34088 37372 34116
rect 23937 34051 23995 34057
rect 23937 34017 23949 34051
rect 23983 34048 23995 34051
rect 24026 34048 24032 34060
rect 23983 34020 24032 34048
rect 23983 34017 23995 34020
rect 23937 34011 23995 34017
rect 24026 34008 24032 34020
rect 24084 34008 24090 34060
rect 25225 34051 25283 34057
rect 25225 34017 25237 34051
rect 25271 34048 25283 34051
rect 25590 34048 25596 34060
rect 25271 34020 25596 34048
rect 25271 34017 25283 34020
rect 25225 34011 25283 34017
rect 25590 34008 25596 34020
rect 25648 34008 25654 34060
rect 27522 34008 27528 34060
rect 27580 34048 27586 34060
rect 27985 34051 28043 34057
rect 27985 34048 27997 34051
rect 27580 34020 27997 34048
rect 27580 34008 27586 34020
rect 27985 34017 27997 34020
rect 28031 34048 28043 34051
rect 30374 34048 30380 34060
rect 28031 34020 30380 34048
rect 28031 34017 28043 34020
rect 27985 34011 28043 34017
rect 30374 34008 30380 34020
rect 30432 34008 30438 34060
rect 31389 34051 31447 34057
rect 31389 34017 31401 34051
rect 31435 34048 31447 34051
rect 35342 34048 35348 34060
rect 31435 34020 35348 34048
rect 31435 34017 31447 34020
rect 31389 34011 31447 34017
rect 35342 34008 35348 34020
rect 35400 34008 35406 34060
rect 36740 34057 36768 34088
rect 37366 34076 37372 34088
rect 37424 34116 37430 34128
rect 41386 34116 41414 34156
rect 48958 34144 48964 34156
rect 49016 34144 49022 34196
rect 37424 34088 41414 34116
rect 37424 34076 37430 34088
rect 42058 34076 42064 34128
rect 42116 34116 42122 34128
rect 42116 34088 42288 34116
rect 42116 34076 42122 34088
rect 36725 34051 36783 34057
rect 36725 34017 36737 34051
rect 36771 34017 36783 34051
rect 36725 34011 36783 34017
rect 36909 34051 36967 34057
rect 36909 34017 36921 34051
rect 36955 34017 36967 34051
rect 36909 34011 36967 34017
rect 26237 33983 26295 33989
rect 26237 33949 26249 33983
rect 26283 33949 26295 33983
rect 26237 33943 26295 33949
rect 23753 33915 23811 33921
rect 23753 33881 23765 33915
rect 23799 33912 23811 33915
rect 26050 33912 26056 33924
rect 23799 33884 26056 33912
rect 23799 33881 23811 33884
rect 23753 33875 23811 33881
rect 26050 33872 26056 33884
rect 26108 33872 26114 33924
rect 26252 33912 26280 33943
rect 29086 33940 29092 33992
rect 29144 33980 29150 33992
rect 29917 33983 29975 33989
rect 29917 33980 29929 33983
rect 29144 33952 29929 33980
rect 29144 33940 29150 33952
rect 29917 33949 29929 33952
rect 29963 33949 29975 33983
rect 29917 33943 29975 33949
rect 31113 33983 31171 33989
rect 31113 33949 31125 33983
rect 31159 33980 31171 33983
rect 32125 33983 32183 33989
rect 32125 33980 32137 33983
rect 31159 33952 32137 33980
rect 31159 33949 31171 33952
rect 31113 33943 31171 33949
rect 32125 33949 32137 33952
rect 32171 33949 32183 33983
rect 32125 33943 32183 33949
rect 26786 33912 26792 33924
rect 26252 33884 26792 33912
rect 26786 33872 26792 33884
rect 26844 33872 26850 33924
rect 28810 33912 28816 33924
rect 27738 33884 28816 33912
rect 28810 33872 28816 33884
rect 28868 33872 28874 33924
rect 32582 33872 32588 33924
rect 32640 33912 32646 33924
rect 36924 33912 36952 34011
rect 38470 34008 38476 34060
rect 38528 34048 38534 34060
rect 38749 34051 38807 34057
rect 38749 34048 38761 34051
rect 38528 34020 38761 34048
rect 38528 34008 38534 34020
rect 38749 34017 38761 34020
rect 38795 34017 38807 34051
rect 38749 34011 38807 34017
rect 42150 34008 42156 34060
rect 42208 34008 42214 34060
rect 42260 34057 42288 34088
rect 42245 34051 42303 34057
rect 42245 34017 42257 34051
rect 42291 34017 42303 34051
rect 42245 34011 42303 34017
rect 37458 33940 37464 33992
rect 37516 33980 37522 33992
rect 38562 33980 38568 33992
rect 37516 33952 38568 33980
rect 37516 33940 37522 33952
rect 38562 33940 38568 33952
rect 38620 33940 38626 33992
rect 38654 33940 38660 33992
rect 38712 33940 38718 33992
rect 41046 33980 41052 33992
rect 39316 33952 41052 33980
rect 39316 33912 39344 33952
rect 41046 33940 41052 33952
rect 41104 33940 41110 33992
rect 41966 33940 41972 33992
rect 42024 33980 42030 33992
rect 42061 33983 42119 33989
rect 42061 33980 42073 33983
rect 42024 33952 42073 33980
rect 42024 33940 42030 33952
rect 42061 33949 42073 33952
rect 42107 33949 42119 33983
rect 42061 33943 42119 33949
rect 49326 33940 49332 33992
rect 49384 33940 49390 33992
rect 49234 33912 49240 33924
rect 32640 33884 36768 33912
rect 36924 33884 39344 33912
rect 39408 33884 49240 33912
rect 32640 33872 32646 33884
rect 22738 33804 22744 33856
rect 22796 33844 22802 33856
rect 23661 33847 23719 33853
rect 23661 33844 23673 33847
rect 22796 33816 23673 33844
rect 22796 33804 22802 33816
rect 23661 33813 23673 33816
rect 23707 33813 23719 33847
rect 23661 33807 23719 33813
rect 24670 33804 24676 33856
rect 24728 33844 24734 33856
rect 24949 33847 25007 33853
rect 24949 33844 24961 33847
rect 24728 33816 24961 33844
rect 24728 33804 24734 33816
rect 24949 33813 24961 33816
rect 24995 33813 25007 33847
rect 24949 33807 25007 33813
rect 25041 33847 25099 33853
rect 25041 33813 25053 33847
rect 25087 33844 25099 33847
rect 27522 33844 27528 33856
rect 25087 33816 27528 33844
rect 25087 33813 25099 33816
rect 25041 33807 25099 33813
rect 27522 33804 27528 33816
rect 27580 33804 27586 33856
rect 31202 33804 31208 33856
rect 31260 33804 31266 33856
rect 33686 33804 33692 33856
rect 33744 33844 33750 33856
rect 35713 33847 35771 33853
rect 35713 33844 35725 33847
rect 33744 33816 35725 33844
rect 33744 33804 33750 33816
rect 35713 33813 35725 33816
rect 35759 33844 35771 33847
rect 36633 33847 36691 33853
rect 36633 33844 36645 33847
rect 35759 33816 36645 33844
rect 35759 33813 35771 33816
rect 35713 33807 35771 33813
rect 36633 33813 36645 33816
rect 36679 33813 36691 33847
rect 36740 33844 36768 33884
rect 37458 33844 37464 33856
rect 36740 33816 37464 33844
rect 36633 33807 36691 33813
rect 37458 33804 37464 33816
rect 37516 33844 37522 33856
rect 37645 33847 37703 33853
rect 37645 33844 37657 33847
rect 37516 33816 37657 33844
rect 37516 33804 37522 33816
rect 37645 33813 37657 33816
rect 37691 33813 37703 33847
rect 37645 33807 37703 33813
rect 37734 33804 37740 33856
rect 37792 33844 37798 33856
rect 38197 33847 38255 33853
rect 38197 33844 38209 33847
rect 37792 33816 38209 33844
rect 37792 33804 37798 33816
rect 38197 33813 38209 33816
rect 38243 33813 38255 33847
rect 38197 33807 38255 33813
rect 38838 33804 38844 33856
rect 38896 33844 38902 33856
rect 39408 33853 39436 33884
rect 49234 33872 49240 33884
rect 49292 33872 49298 33924
rect 39393 33847 39451 33853
rect 39393 33844 39405 33847
rect 38896 33816 39405 33844
rect 38896 33804 38902 33816
rect 39393 33813 39405 33816
rect 39439 33813 39451 33847
rect 39393 33807 39451 33813
rect 41414 33804 41420 33856
rect 41472 33844 41478 33856
rect 41693 33847 41751 33853
rect 41693 33844 41705 33847
rect 41472 33816 41705 33844
rect 41472 33804 41478 33816
rect 41693 33813 41705 33816
rect 41739 33813 41751 33847
rect 41693 33807 41751 33813
rect 41874 33804 41880 33856
rect 41932 33844 41938 33856
rect 49145 33847 49203 33853
rect 49145 33844 49157 33847
rect 41932 33816 49157 33844
rect 41932 33804 41938 33816
rect 49145 33813 49157 33816
rect 49191 33813 49203 33847
rect 49145 33807 49203 33813
rect 1104 33754 49864 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 27950 33754
rect 28002 33702 28014 33754
rect 28066 33702 28078 33754
rect 28130 33702 28142 33754
rect 28194 33702 28206 33754
rect 28258 33702 37950 33754
rect 38002 33702 38014 33754
rect 38066 33702 38078 33754
rect 38130 33702 38142 33754
rect 38194 33702 38206 33754
rect 38258 33702 47950 33754
rect 48002 33702 48014 33754
rect 48066 33702 48078 33754
rect 48130 33702 48142 33754
rect 48194 33702 48206 33754
rect 48258 33702 49864 33754
rect 1104 33680 49864 33702
rect 24026 33640 24032 33652
rect 23124 33612 24032 33640
rect 23124 33581 23152 33612
rect 24026 33600 24032 33612
rect 24084 33600 24090 33652
rect 25041 33643 25099 33649
rect 25041 33609 25053 33643
rect 25087 33640 25099 33643
rect 25130 33640 25136 33652
rect 25087 33612 25136 33640
rect 25087 33609 25099 33612
rect 25041 33603 25099 33609
rect 25130 33600 25136 33612
rect 25188 33600 25194 33652
rect 28718 33600 28724 33652
rect 28776 33600 28782 33652
rect 29086 33600 29092 33652
rect 29144 33600 29150 33652
rect 34054 33640 34060 33652
rect 30300 33612 34060 33640
rect 23109 33575 23167 33581
rect 23109 33541 23121 33575
rect 23155 33541 23167 33575
rect 24762 33572 24768 33584
rect 24334 33544 24768 33572
rect 23109 33535 23167 33541
rect 24762 33532 24768 33544
rect 24820 33532 24826 33584
rect 25130 33464 25136 33516
rect 25188 33504 25194 33516
rect 25409 33507 25467 33513
rect 25409 33504 25421 33507
rect 25188 33476 25421 33504
rect 25188 33464 25194 33476
rect 25409 33473 25421 33476
rect 25455 33473 25467 33507
rect 25409 33467 25467 33473
rect 25501 33507 25559 33513
rect 25501 33473 25513 33507
rect 25547 33504 25559 33507
rect 27430 33504 27436 33516
rect 25547 33476 27436 33504
rect 25547 33473 25559 33476
rect 25501 33467 25559 33473
rect 27430 33464 27436 33476
rect 27488 33464 27494 33516
rect 28552 33476 29500 33504
rect 21082 33396 21088 33448
rect 21140 33436 21146 33448
rect 21726 33436 21732 33448
rect 21140 33408 21732 33436
rect 21140 33396 21146 33408
rect 21726 33396 21732 33408
rect 21784 33436 21790 33448
rect 22833 33439 22891 33445
rect 22833 33436 22845 33439
rect 21784 33408 22845 33436
rect 21784 33396 21790 33408
rect 22833 33405 22845 33408
rect 22879 33405 22891 33439
rect 22833 33399 22891 33405
rect 24578 33396 24584 33448
rect 24636 33436 24642 33448
rect 25593 33439 25651 33445
rect 25593 33436 25605 33439
rect 24636 33408 25605 33436
rect 24636 33396 24642 33408
rect 25593 33405 25605 33408
rect 25639 33405 25651 33439
rect 25593 33399 25651 33405
rect 27062 33396 27068 33448
rect 27120 33436 27126 33448
rect 28552 33436 28580 33476
rect 27120 33408 28580 33436
rect 27120 33396 27126 33408
rect 29178 33396 29184 33448
rect 29236 33396 29242 33448
rect 29365 33439 29423 33445
rect 29365 33405 29377 33439
rect 29411 33405 29423 33439
rect 29472 33436 29500 33476
rect 29638 33464 29644 33516
rect 29696 33504 29702 33516
rect 30300 33513 30328 33612
rect 34054 33600 34060 33612
rect 34112 33600 34118 33652
rect 34882 33600 34888 33652
rect 34940 33640 34946 33652
rect 38841 33643 38899 33649
rect 38841 33640 38853 33643
rect 34940 33612 38853 33640
rect 34940 33600 34946 33612
rect 38841 33609 38853 33612
rect 38887 33609 38899 33643
rect 38841 33603 38899 33609
rect 39301 33643 39359 33649
rect 39301 33609 39313 33643
rect 39347 33640 39359 33643
rect 42334 33640 42340 33652
rect 39347 33612 42340 33640
rect 39347 33609 39359 33612
rect 39301 33603 39359 33609
rect 42334 33600 42340 33612
rect 42392 33600 42398 33652
rect 30374 33532 30380 33584
rect 30432 33532 30438 33584
rect 33870 33532 33876 33584
rect 33928 33572 33934 33584
rect 34241 33575 34299 33581
rect 34241 33572 34253 33575
rect 33928 33544 34253 33572
rect 33928 33532 33934 33544
rect 34241 33541 34253 33544
rect 34287 33541 34299 33575
rect 34241 33535 34299 33541
rect 34974 33532 34980 33584
rect 35032 33532 35038 33584
rect 37458 33532 37464 33584
rect 37516 33572 37522 33584
rect 40862 33572 40868 33584
rect 37516 33544 40868 33572
rect 37516 33532 37522 33544
rect 40862 33532 40868 33544
rect 40920 33532 40926 33584
rect 42610 33572 42616 33584
rect 41814 33544 42616 33572
rect 42610 33532 42616 33544
rect 42668 33572 42674 33584
rect 43438 33572 43444 33584
rect 42668 33544 43444 33572
rect 42668 33532 42674 33544
rect 43438 33532 43444 33544
rect 43496 33532 43502 33584
rect 30285 33507 30343 33513
rect 30285 33504 30297 33507
rect 29696 33476 30297 33504
rect 29696 33464 29702 33476
rect 30285 33473 30297 33476
rect 30331 33473 30343 33507
rect 30392 33504 30420 33532
rect 30392 33476 30512 33504
rect 30285 33467 30343 33473
rect 30484 33445 30512 33476
rect 33962 33464 33968 33516
rect 34020 33464 34026 33516
rect 35636 33476 37044 33504
rect 30377 33439 30435 33445
rect 30377 33436 30389 33439
rect 29472 33408 30389 33436
rect 29365 33399 29423 33405
rect 30377 33405 30389 33408
rect 30423 33405 30435 33439
rect 30377 33399 30435 33405
rect 30469 33439 30527 33445
rect 30469 33405 30481 33439
rect 30515 33405 30527 33439
rect 30469 33399 30527 33405
rect 29380 33368 29408 33399
rect 34238 33396 34244 33448
rect 34296 33436 34302 33448
rect 34698 33436 34704 33448
rect 34296 33408 34704 33436
rect 34296 33396 34302 33408
rect 34698 33396 34704 33408
rect 34756 33436 34762 33448
rect 35636 33436 35664 33476
rect 34756 33408 35664 33436
rect 35713 33439 35771 33445
rect 34756 33396 34762 33408
rect 35713 33405 35725 33439
rect 35759 33436 35771 33439
rect 36906 33436 36912 33448
rect 35759 33408 36912 33436
rect 35759 33405 35771 33408
rect 35713 33399 35771 33405
rect 36906 33396 36912 33408
rect 36964 33396 36970 33448
rect 37016 33436 37044 33476
rect 37826 33464 37832 33516
rect 37884 33504 37890 33516
rect 38657 33507 38715 33513
rect 38657 33504 38669 33507
rect 37884 33476 38669 33504
rect 37884 33464 37890 33476
rect 38657 33473 38669 33476
rect 38703 33473 38715 33507
rect 38657 33467 38715 33473
rect 39206 33464 39212 33516
rect 39264 33464 39270 33516
rect 40218 33504 40224 33516
rect 39316 33476 40224 33504
rect 37921 33439 37979 33445
rect 37921 33436 37933 33439
rect 37016 33408 37933 33436
rect 37921 33405 37933 33408
rect 37967 33405 37979 33439
rect 37921 33399 37979 33405
rect 38105 33439 38163 33445
rect 38105 33405 38117 33439
rect 38151 33436 38163 33439
rect 39316 33436 39344 33476
rect 40218 33464 40224 33476
rect 40276 33464 40282 33516
rect 38151 33408 39344 33436
rect 39393 33439 39451 33445
rect 38151 33405 38163 33408
rect 38105 33399 38163 33405
rect 39393 33405 39405 33439
rect 39439 33405 39451 33439
rect 39393 33399 39451 33405
rect 30558 33368 30564 33380
rect 29380 33340 30564 33368
rect 30558 33328 30564 33340
rect 30616 33328 30622 33380
rect 36998 33368 37004 33380
rect 35268 33340 37004 33368
rect 22370 33260 22376 33312
rect 22428 33300 22434 33312
rect 24581 33303 24639 33309
rect 24581 33300 24593 33303
rect 22428 33272 24593 33300
rect 22428 33260 22434 33272
rect 24581 33269 24593 33272
rect 24627 33300 24639 33303
rect 28350 33300 28356 33312
rect 24627 33272 28356 33300
rect 24627 33269 24639 33272
rect 24581 33263 24639 33269
rect 28350 33260 28356 33272
rect 28408 33260 28414 33312
rect 29914 33260 29920 33312
rect 29972 33260 29978 33312
rect 31570 33260 31576 33312
rect 31628 33300 31634 33312
rect 35268 33300 35296 33340
rect 36998 33328 37004 33340
rect 37056 33328 37062 33380
rect 37458 33328 37464 33380
rect 37516 33328 37522 33380
rect 31628 33272 35296 33300
rect 31628 33260 31634 33272
rect 35894 33260 35900 33312
rect 35952 33300 35958 33312
rect 36173 33303 36231 33309
rect 36173 33300 36185 33303
rect 35952 33272 36185 33300
rect 35952 33260 35958 33272
rect 36173 33269 36185 33272
rect 36219 33269 36231 33303
rect 37936 33300 37964 33399
rect 38194 33328 38200 33380
rect 38252 33368 38258 33380
rect 39408 33368 39436 33399
rect 40310 33396 40316 33448
rect 40368 33396 40374 33448
rect 40586 33396 40592 33448
rect 40644 33436 40650 33448
rect 41138 33436 41144 33448
rect 40644 33408 41144 33436
rect 40644 33396 40650 33408
rect 41138 33396 41144 33408
rect 41196 33396 41202 33448
rect 38252 33340 39436 33368
rect 38252 33328 38258 33340
rect 38838 33300 38844 33312
rect 37936 33272 38844 33300
rect 36173 33263 36231 33269
rect 38838 33260 38844 33272
rect 38896 33260 38902 33312
rect 42058 33260 42064 33312
rect 42116 33260 42122 33312
rect 1104 33210 49864 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 32950 33210
rect 33002 33158 33014 33210
rect 33066 33158 33078 33210
rect 33130 33158 33142 33210
rect 33194 33158 33206 33210
rect 33258 33158 42950 33210
rect 43002 33158 43014 33210
rect 43066 33158 43078 33210
rect 43130 33158 43142 33210
rect 43194 33158 43206 33210
rect 43258 33158 49864 33210
rect 1104 33136 49864 33158
rect 22830 33056 22836 33108
rect 22888 33096 22894 33108
rect 23290 33096 23296 33108
rect 22888 33068 23296 33096
rect 22888 33056 22894 33068
rect 23290 33056 23296 33068
rect 23348 33056 23354 33108
rect 27522 33056 27528 33108
rect 27580 33096 27586 33108
rect 28445 33099 28503 33105
rect 28445 33096 28457 33099
rect 27580 33068 28457 33096
rect 27580 33056 27586 33068
rect 28445 33065 28457 33068
rect 28491 33065 28503 33099
rect 28445 33059 28503 33065
rect 28902 33056 28908 33108
rect 28960 33096 28966 33108
rect 30929 33099 30987 33105
rect 28960 33068 29040 33096
rect 28960 33056 28966 33068
rect 26050 32988 26056 33040
rect 26108 33028 26114 33040
rect 26108 33000 27384 33028
rect 26108 32988 26114 33000
rect 21361 32963 21419 32969
rect 21361 32929 21373 32963
rect 21407 32960 21419 32963
rect 22370 32960 22376 32972
rect 21407 32932 22376 32960
rect 21407 32929 21419 32932
rect 21361 32923 21419 32929
rect 22370 32920 22376 32932
rect 22428 32920 22434 32972
rect 23658 32960 23664 32972
rect 22480 32932 23664 32960
rect 21082 32852 21088 32904
rect 21140 32852 21146 32904
rect 22480 32878 22508 32932
rect 23658 32920 23664 32932
rect 23716 32920 23722 32972
rect 26786 32920 26792 32972
rect 26844 32960 26850 32972
rect 27065 32963 27123 32969
rect 27065 32960 27077 32963
rect 26844 32932 27077 32960
rect 26844 32920 26850 32932
rect 27065 32929 27077 32932
rect 27111 32929 27123 32963
rect 27065 32923 27123 32929
rect 27249 32963 27307 32969
rect 27249 32929 27261 32963
rect 27295 32929 27307 32963
rect 27249 32923 27307 32929
rect 26053 32895 26111 32901
rect 26053 32892 26065 32895
rect 22756 32864 26065 32892
rect 12066 32716 12072 32768
rect 12124 32756 12130 32768
rect 22756 32756 22784 32864
rect 26053 32861 26065 32864
rect 26099 32892 26111 32895
rect 26878 32892 26884 32904
rect 26099 32864 26884 32892
rect 26099 32861 26111 32864
rect 26053 32855 26111 32861
rect 26878 32852 26884 32864
rect 26936 32892 26942 32904
rect 26973 32895 27031 32901
rect 26973 32892 26985 32895
rect 26936 32864 26985 32892
rect 26936 32852 26942 32864
rect 26973 32861 26985 32864
rect 27019 32861 27031 32895
rect 26973 32855 27031 32861
rect 12124 32728 22784 32756
rect 12124 32716 12130 32728
rect 23658 32716 23664 32768
rect 23716 32756 23722 32768
rect 24762 32756 24768 32768
rect 23716 32728 24768 32756
rect 23716 32716 23722 32728
rect 24762 32716 24768 32728
rect 24820 32716 24826 32768
rect 26602 32716 26608 32768
rect 26660 32716 26666 32768
rect 27264 32756 27292 32923
rect 27356 32824 27384 33000
rect 28350 32920 28356 32972
rect 28408 32960 28414 32972
rect 28718 32960 28724 32972
rect 28408 32932 28724 32960
rect 28408 32920 28414 32932
rect 28718 32920 28724 32932
rect 28776 32920 28782 32972
rect 28905 32963 28963 32969
rect 28905 32929 28917 32963
rect 28951 32960 28963 32963
rect 29012 32960 29040 33068
rect 30929 33065 30941 33099
rect 30975 33096 30987 33099
rect 31846 33096 31852 33108
rect 30975 33068 31852 33096
rect 30975 33065 30987 33068
rect 30929 33059 30987 33065
rect 31846 33056 31852 33068
rect 31904 33056 31910 33108
rect 32582 33056 32588 33108
rect 32640 33096 32646 33108
rect 36522 33099 36580 33105
rect 36522 33096 36534 33099
rect 32640 33068 36534 33096
rect 32640 33056 32646 33068
rect 36522 33065 36534 33068
rect 36568 33065 36580 33099
rect 36522 33059 36580 33065
rect 36906 33056 36912 33108
rect 36964 33096 36970 33108
rect 38381 33099 38439 33105
rect 38381 33096 38393 33099
rect 36964 33068 38393 33096
rect 36964 33056 36970 33068
rect 38381 33065 38393 33068
rect 38427 33065 38439 33099
rect 38381 33059 38439 33065
rect 34885 33031 34943 33037
rect 34885 32997 34897 33031
rect 34931 33028 34943 33031
rect 38013 33031 38071 33037
rect 34931 33000 36400 33028
rect 34931 32997 34943 33000
rect 34885 32991 34943 32997
rect 28951 32932 29040 32960
rect 29089 32963 29147 32969
rect 28951 32929 28963 32932
rect 28905 32923 28963 32929
rect 29089 32929 29101 32963
rect 29135 32960 29147 32963
rect 29270 32960 29276 32972
rect 29135 32932 29276 32960
rect 29135 32929 29147 32932
rect 29089 32923 29147 32929
rect 29270 32920 29276 32932
rect 29328 32920 29334 32972
rect 30374 32920 30380 32972
rect 30432 32920 30438 32972
rect 31478 32920 31484 32972
rect 31536 32920 31542 32972
rect 35529 32963 35587 32969
rect 35529 32929 35541 32963
rect 35575 32929 35587 32963
rect 36372 32960 36400 33000
rect 38013 32997 38025 33031
rect 38059 33028 38071 33031
rect 40586 33028 40592 33040
rect 38059 33000 40592 33028
rect 38059 32997 38071 33000
rect 38013 32991 38071 32997
rect 40586 32988 40592 33000
rect 40644 32988 40650 33040
rect 48774 33028 48780 33040
rect 41386 33000 48780 33028
rect 37274 32960 37280 32972
rect 36372 32932 37280 32960
rect 35529 32923 35587 32929
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32892 28871 32895
rect 31018 32892 31024 32904
rect 28859 32864 31024 32892
rect 28859 32861 28871 32864
rect 28813 32855 28871 32861
rect 31018 32852 31024 32864
rect 31076 32852 31082 32904
rect 31389 32895 31447 32901
rect 31389 32861 31401 32895
rect 31435 32892 31447 32895
rect 32122 32892 32128 32904
rect 31435 32864 32128 32892
rect 31435 32861 31447 32864
rect 31389 32855 31447 32861
rect 32122 32852 32128 32864
rect 32180 32852 32186 32904
rect 34517 32895 34575 32901
rect 34517 32861 34529 32895
rect 34563 32892 34575 32895
rect 35253 32895 35311 32901
rect 35253 32892 35265 32895
rect 34563 32864 35265 32892
rect 34563 32861 34575 32864
rect 34517 32855 34575 32861
rect 35253 32861 35265 32864
rect 35299 32861 35311 32895
rect 35253 32855 35311 32861
rect 30101 32827 30159 32833
rect 27356 32796 29776 32824
rect 28994 32756 29000 32768
rect 27264 32728 29000 32756
rect 28994 32716 29000 32728
rect 29052 32716 29058 32768
rect 29748 32765 29776 32796
rect 30101 32793 30113 32827
rect 30147 32824 30159 32827
rect 34606 32824 34612 32836
rect 30147 32796 34612 32824
rect 30147 32793 30159 32796
rect 30101 32787 30159 32793
rect 34606 32784 34612 32796
rect 34664 32784 34670 32836
rect 35544 32824 35572 32923
rect 37274 32920 37280 32932
rect 37332 32920 37338 32972
rect 37550 32920 37556 32972
rect 37608 32960 37614 32972
rect 38933 32963 38991 32969
rect 38933 32960 38945 32963
rect 37608 32932 38945 32960
rect 37608 32920 37614 32932
rect 38933 32929 38945 32932
rect 38979 32929 38991 32963
rect 38933 32923 38991 32929
rect 40678 32920 40684 32972
rect 40736 32960 40742 32972
rect 40865 32963 40923 32969
rect 40865 32960 40877 32963
rect 40736 32932 40877 32960
rect 40736 32920 40742 32932
rect 40865 32929 40877 32932
rect 40911 32929 40923 32963
rect 40865 32923 40923 32929
rect 41049 32963 41107 32969
rect 41049 32929 41061 32963
rect 41095 32960 41107 32963
rect 41230 32960 41236 32972
rect 41095 32932 41236 32960
rect 41095 32929 41107 32932
rect 41049 32923 41107 32929
rect 41230 32920 41236 32932
rect 41288 32920 41294 32972
rect 36262 32852 36268 32904
rect 36320 32852 36326 32904
rect 38746 32852 38752 32904
rect 38804 32852 38810 32904
rect 38841 32895 38899 32901
rect 38841 32861 38853 32895
rect 38887 32892 38899 32895
rect 39022 32892 39028 32904
rect 38887 32864 39028 32892
rect 38887 32861 38899 32864
rect 38841 32855 38899 32861
rect 39022 32852 39028 32864
rect 39080 32852 39086 32904
rect 40770 32852 40776 32904
rect 40828 32852 40834 32904
rect 35544 32796 36216 32824
rect 29733 32759 29791 32765
rect 29733 32725 29745 32759
rect 29779 32725 29791 32759
rect 29733 32719 29791 32725
rect 30193 32759 30251 32765
rect 30193 32725 30205 32759
rect 30239 32756 30251 32759
rect 30926 32756 30932 32768
rect 30239 32728 30932 32756
rect 30239 32725 30251 32728
rect 30193 32719 30251 32725
rect 30926 32716 30932 32728
rect 30984 32716 30990 32768
rect 31294 32716 31300 32768
rect 31352 32716 31358 32768
rect 34054 32716 34060 32768
rect 34112 32756 34118 32768
rect 34974 32756 34980 32768
rect 34112 32728 34980 32756
rect 34112 32716 34118 32728
rect 34974 32716 34980 32728
rect 35032 32716 35038 32768
rect 35345 32759 35403 32765
rect 35345 32725 35357 32759
rect 35391 32756 35403 32759
rect 35894 32756 35900 32768
rect 35391 32728 35900 32756
rect 35391 32725 35403 32728
rect 35345 32719 35403 32725
rect 35894 32716 35900 32728
rect 35952 32756 35958 32768
rect 36081 32759 36139 32765
rect 36081 32756 36093 32759
rect 35952 32728 36093 32756
rect 35952 32716 35958 32728
rect 36081 32725 36093 32728
rect 36127 32725 36139 32759
rect 36188 32756 36216 32796
rect 37274 32784 37280 32836
rect 37332 32784 37338 32836
rect 37826 32784 37832 32836
rect 37884 32824 37890 32836
rect 41386 32824 41414 33000
rect 48774 32988 48780 33000
rect 48832 32988 48838 33040
rect 41782 32920 41788 32972
rect 41840 32960 41846 32972
rect 42061 32963 42119 32969
rect 42061 32960 42073 32963
rect 41840 32932 42073 32960
rect 41840 32920 41846 32932
rect 42061 32929 42073 32932
rect 42107 32929 42119 32963
rect 42061 32923 42119 32929
rect 42242 32920 42248 32972
rect 42300 32920 42306 32972
rect 41969 32895 42027 32901
rect 41969 32861 41981 32895
rect 42015 32892 42027 32895
rect 42334 32892 42340 32904
rect 42015 32864 42340 32892
rect 42015 32861 42027 32864
rect 41969 32855 42027 32861
rect 42334 32852 42340 32864
rect 42392 32852 42398 32904
rect 43806 32852 43812 32904
rect 43864 32852 43870 32904
rect 49326 32852 49332 32904
rect 49384 32852 49390 32904
rect 37884 32796 41414 32824
rect 37884 32784 37890 32796
rect 38286 32756 38292 32768
rect 36188 32728 38292 32756
rect 36081 32719 36139 32725
rect 38286 32716 38292 32728
rect 38344 32716 38350 32768
rect 38746 32716 38752 32768
rect 38804 32756 38810 32768
rect 39298 32756 39304 32768
rect 38804 32728 39304 32756
rect 38804 32716 38810 32728
rect 39298 32716 39304 32728
rect 39356 32716 39362 32768
rect 40218 32716 40224 32768
rect 40276 32756 40282 32768
rect 40405 32759 40463 32765
rect 40405 32756 40417 32759
rect 40276 32728 40417 32756
rect 40276 32716 40282 32728
rect 40405 32725 40417 32728
rect 40451 32725 40463 32759
rect 40405 32719 40463 32725
rect 41046 32716 41052 32768
rect 41104 32756 41110 32768
rect 41601 32759 41659 32765
rect 41601 32756 41613 32759
rect 41104 32728 41613 32756
rect 41104 32716 41110 32728
rect 41601 32725 41613 32728
rect 41647 32725 41659 32759
rect 41601 32719 41659 32725
rect 43625 32759 43683 32765
rect 43625 32725 43637 32759
rect 43671 32756 43683 32759
rect 47210 32756 47216 32768
rect 43671 32728 47216 32756
rect 43671 32725 43683 32728
rect 43625 32719 43683 32725
rect 47210 32716 47216 32728
rect 47268 32716 47274 32768
rect 49142 32716 49148 32768
rect 49200 32716 49206 32768
rect 1104 32666 49864 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 27950 32666
rect 28002 32614 28014 32666
rect 28066 32614 28078 32666
rect 28130 32614 28142 32666
rect 28194 32614 28206 32666
rect 28258 32614 37950 32666
rect 38002 32614 38014 32666
rect 38066 32614 38078 32666
rect 38130 32614 38142 32666
rect 38194 32614 38206 32666
rect 38258 32614 47950 32666
rect 48002 32614 48014 32666
rect 48066 32614 48078 32666
rect 48130 32614 48142 32666
rect 48194 32614 48206 32666
rect 48258 32614 49864 32666
rect 1104 32592 49864 32614
rect 17218 32512 17224 32564
rect 17276 32512 17282 32564
rect 17678 32512 17684 32564
rect 17736 32512 17742 32564
rect 23768 32524 25544 32552
rect 23768 32496 23796 32524
rect 13446 32444 13452 32496
rect 13504 32484 13510 32496
rect 23750 32484 23756 32496
rect 13504 32456 23756 32484
rect 13504 32444 13510 32456
rect 23750 32444 23756 32456
rect 23808 32444 23814 32496
rect 24762 32444 24768 32496
rect 24820 32444 24826 32496
rect 934 32376 940 32428
rect 992 32416 998 32428
rect 1765 32419 1823 32425
rect 1765 32416 1777 32419
rect 992 32388 1777 32416
rect 992 32376 998 32388
rect 1765 32385 1777 32388
rect 1811 32385 1823 32419
rect 1765 32379 1823 32385
rect 17589 32419 17647 32425
rect 17589 32385 17601 32419
rect 17635 32416 17647 32419
rect 18601 32419 18659 32425
rect 18601 32416 18613 32419
rect 17635 32388 18613 32416
rect 17635 32385 17647 32388
rect 17589 32379 17647 32385
rect 18601 32385 18613 32388
rect 18647 32385 18659 32419
rect 18601 32379 18659 32385
rect 22646 32376 22652 32428
rect 22704 32416 22710 32428
rect 23474 32416 23480 32428
rect 22704 32388 23480 32416
rect 22704 32376 22710 32388
rect 23474 32376 23480 32388
rect 23532 32416 23538 32428
rect 23845 32419 23903 32425
rect 23845 32416 23857 32419
rect 23532 32388 23857 32416
rect 23532 32376 23538 32388
rect 23845 32385 23857 32388
rect 23891 32385 23903 32419
rect 23845 32379 23903 32385
rect 17865 32351 17923 32357
rect 17865 32317 17877 32351
rect 17911 32348 17923 32351
rect 22830 32348 22836 32360
rect 17911 32320 22836 32348
rect 17911 32317 17923 32320
rect 17865 32311 17923 32317
rect 22830 32308 22836 32320
rect 22888 32308 22894 32360
rect 24118 32308 24124 32360
rect 24176 32308 24182 32360
rect 24762 32308 24768 32360
rect 24820 32348 24826 32360
rect 25516 32348 25544 32524
rect 25590 32512 25596 32564
rect 25648 32552 25654 32564
rect 26050 32552 26056 32564
rect 25648 32524 26056 32552
rect 25648 32512 25654 32524
rect 26050 32512 26056 32524
rect 26108 32512 26114 32564
rect 27249 32555 27307 32561
rect 27249 32521 27261 32555
rect 27295 32552 27307 32555
rect 31294 32552 31300 32564
rect 27295 32524 31300 32552
rect 27295 32521 27307 32524
rect 27249 32515 27307 32521
rect 31294 32512 31300 32524
rect 31352 32512 31358 32564
rect 31570 32512 31576 32564
rect 31628 32552 31634 32564
rect 34241 32555 34299 32561
rect 34241 32552 34253 32555
rect 31628 32524 34253 32552
rect 31628 32512 31634 32524
rect 34241 32521 34253 32524
rect 34287 32552 34299 32555
rect 35069 32555 35127 32561
rect 34287 32524 35020 32552
rect 34287 32521 34299 32524
rect 34241 32515 34299 32521
rect 26602 32444 26608 32496
rect 26660 32484 26666 32496
rect 31110 32484 31116 32496
rect 26660 32456 31116 32484
rect 26660 32444 26666 32456
rect 31110 32444 31116 32456
rect 31168 32444 31174 32496
rect 34054 32484 34060 32496
rect 33994 32456 34060 32484
rect 34054 32444 34060 32456
rect 34112 32444 34118 32496
rect 34992 32484 35020 32524
rect 35069 32521 35081 32555
rect 35115 32552 35127 32555
rect 37734 32552 37740 32564
rect 35115 32524 37740 32552
rect 35115 32521 35127 32524
rect 35069 32515 35127 32521
rect 37734 32512 37740 32524
rect 37792 32512 37798 32564
rect 40310 32552 40316 32564
rect 39316 32524 40316 32552
rect 34992 32456 35296 32484
rect 27617 32419 27675 32425
rect 27617 32385 27629 32419
rect 27663 32416 27675 32419
rect 28813 32419 28871 32425
rect 28813 32416 28825 32419
rect 27663 32388 28825 32416
rect 27663 32385 27675 32388
rect 27617 32379 27675 32385
rect 28813 32385 28825 32388
rect 28859 32385 28871 32419
rect 28813 32379 28871 32385
rect 29086 32376 29092 32428
rect 29144 32416 29150 32428
rect 30374 32416 30380 32428
rect 29144 32388 30380 32416
rect 29144 32376 29150 32388
rect 30374 32376 30380 32388
rect 30432 32376 30438 32428
rect 35066 32416 35072 32428
rect 34072 32388 35072 32416
rect 27709 32351 27767 32357
rect 27709 32348 27721 32351
rect 24820 32320 25452 32348
rect 25516 32320 27721 32348
rect 24820 32308 24826 32320
rect 25424 32280 25452 32320
rect 27709 32317 27721 32320
rect 27755 32317 27767 32351
rect 27709 32311 27767 32317
rect 26418 32280 26424 32292
rect 25424 32252 26424 32280
rect 26418 32240 26424 32252
rect 26476 32240 26482 32292
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 7466 32212 7472 32224
rect 1627 32184 7472 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 7466 32172 7472 32184
rect 7524 32172 7530 32224
rect 20254 32172 20260 32224
rect 20312 32212 20318 32224
rect 25958 32212 25964 32224
rect 20312 32184 25964 32212
rect 20312 32172 20318 32184
rect 25958 32172 25964 32184
rect 26016 32212 26022 32224
rect 27154 32212 27160 32224
rect 26016 32184 27160 32212
rect 26016 32172 26022 32184
rect 27154 32172 27160 32184
rect 27212 32172 27218 32224
rect 27724 32212 27752 32311
rect 27890 32308 27896 32360
rect 27948 32308 27954 32360
rect 28258 32308 28264 32360
rect 28316 32348 28322 32360
rect 28442 32348 28448 32360
rect 28316 32320 28448 32348
rect 28316 32308 28322 32320
rect 28442 32308 28448 32320
rect 28500 32308 28506 32360
rect 29270 32348 29276 32360
rect 28552 32320 29276 32348
rect 28350 32240 28356 32292
rect 28408 32280 28414 32292
rect 28552 32280 28580 32320
rect 29270 32308 29276 32320
rect 29328 32308 29334 32360
rect 32122 32308 32128 32360
rect 32180 32348 32186 32360
rect 32493 32351 32551 32357
rect 32493 32348 32505 32351
rect 32180 32320 32505 32348
rect 32180 32308 32186 32320
rect 32493 32317 32505 32320
rect 32539 32317 32551 32351
rect 32493 32311 32551 32317
rect 32769 32351 32827 32357
rect 32769 32317 32781 32351
rect 32815 32348 32827 32351
rect 34072 32348 34100 32388
rect 35066 32376 35072 32388
rect 35124 32376 35130 32428
rect 35158 32376 35164 32428
rect 35216 32376 35222 32428
rect 35268 32357 35296 32456
rect 37642 32444 37648 32496
rect 37700 32484 37706 32496
rect 37918 32484 37924 32496
rect 37700 32456 37924 32484
rect 37700 32444 37706 32456
rect 37918 32444 37924 32456
rect 37976 32444 37982 32496
rect 36262 32376 36268 32428
rect 36320 32416 36326 32428
rect 39316 32425 39344 32524
rect 40310 32512 40316 32524
rect 40368 32512 40374 32564
rect 41322 32512 41328 32564
rect 41380 32552 41386 32564
rect 49142 32552 49148 32564
rect 41380 32524 49148 32552
rect 41380 32512 41386 32524
rect 49142 32512 49148 32524
rect 49200 32512 49206 32564
rect 39666 32444 39672 32496
rect 39724 32484 39730 32496
rect 39724 32456 40066 32484
rect 39724 32444 39730 32456
rect 39301 32419 39359 32425
rect 39301 32416 39313 32419
rect 36320 32388 39313 32416
rect 36320 32376 36326 32388
rect 39301 32385 39313 32388
rect 39347 32385 39359 32419
rect 39301 32379 39359 32385
rect 42518 32376 42524 32428
rect 42576 32416 42582 32428
rect 45005 32419 45063 32425
rect 45005 32416 45017 32419
rect 42576 32388 45017 32416
rect 42576 32376 42582 32388
rect 45005 32385 45017 32388
rect 45051 32385 45063 32419
rect 45005 32379 45063 32385
rect 48774 32376 48780 32428
rect 48832 32376 48838 32428
rect 32815 32320 34100 32348
rect 35253 32351 35311 32357
rect 32815 32317 32827 32320
rect 32769 32311 32827 32317
rect 35253 32317 35265 32351
rect 35299 32317 35311 32351
rect 35253 32311 35311 32317
rect 36078 32308 36084 32360
rect 36136 32348 36142 32360
rect 39577 32351 39635 32357
rect 36136 32320 39344 32348
rect 36136 32308 36142 32320
rect 39316 32292 39344 32320
rect 39577 32317 39589 32351
rect 39623 32348 39635 32351
rect 42058 32348 42064 32360
rect 39623 32320 42064 32348
rect 39623 32317 39635 32320
rect 39577 32311 39635 32317
rect 42058 32308 42064 32320
rect 42116 32308 42122 32360
rect 48498 32308 48504 32360
rect 48556 32308 48562 32360
rect 29178 32280 29184 32292
rect 28408 32252 28580 32280
rect 28828 32252 29184 32280
rect 28408 32240 28414 32252
rect 28445 32215 28503 32221
rect 28445 32212 28457 32215
rect 27724 32184 28457 32212
rect 28445 32181 28457 32184
rect 28491 32212 28503 32215
rect 28828 32212 28856 32252
rect 29178 32240 29184 32252
rect 29236 32240 29242 32292
rect 34440 32252 35112 32280
rect 28491 32184 28856 32212
rect 28491 32181 28503 32184
rect 28445 32175 28503 32181
rect 32214 32172 32220 32224
rect 32272 32212 32278 32224
rect 34440 32212 34468 32252
rect 32272 32184 34468 32212
rect 32272 32172 32278 32184
rect 34514 32172 34520 32224
rect 34572 32212 34578 32224
rect 34701 32215 34759 32221
rect 34701 32212 34713 32215
rect 34572 32184 34713 32212
rect 34572 32172 34578 32184
rect 34701 32181 34713 32184
rect 34747 32181 34759 32215
rect 35084 32212 35112 32252
rect 39298 32240 39304 32292
rect 39356 32240 39362 32292
rect 45278 32280 45284 32292
rect 40604 32252 45284 32280
rect 37826 32212 37832 32224
rect 35084 32184 37832 32212
rect 34701 32175 34759 32181
rect 37826 32172 37832 32184
rect 37884 32172 37890 32224
rect 39666 32172 39672 32224
rect 39724 32212 39730 32224
rect 40604 32212 40632 32252
rect 45278 32240 45284 32252
rect 45336 32240 45342 32292
rect 39724 32184 40632 32212
rect 39724 32172 39730 32184
rect 40954 32172 40960 32224
rect 41012 32212 41018 32224
rect 41049 32215 41107 32221
rect 41049 32212 41061 32215
rect 41012 32184 41061 32212
rect 41012 32172 41018 32184
rect 41049 32181 41061 32184
rect 41095 32181 41107 32215
rect 41049 32175 41107 32181
rect 42794 32172 42800 32224
rect 42852 32172 42858 32224
rect 44818 32172 44824 32224
rect 44876 32172 44882 32224
rect 1104 32122 49864 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 32950 32122
rect 33002 32070 33014 32122
rect 33066 32070 33078 32122
rect 33130 32070 33142 32122
rect 33194 32070 33206 32122
rect 33258 32070 42950 32122
rect 43002 32070 43014 32122
rect 43066 32070 43078 32122
rect 43130 32070 43142 32122
rect 43194 32070 43206 32122
rect 43258 32070 49864 32122
rect 1104 32048 49864 32070
rect 22646 32008 22652 32020
rect 22388 31980 22652 32008
rect 22281 31875 22339 31881
rect 22281 31841 22293 31875
rect 22327 31872 22339 31875
rect 22388 31872 22416 31980
rect 22646 31968 22652 31980
rect 22704 31968 22710 32020
rect 24026 31968 24032 32020
rect 24084 31968 24090 32020
rect 27062 32008 27068 32020
rect 25792 31980 27068 32008
rect 23750 31900 23756 31952
rect 23808 31940 23814 31952
rect 23808 31912 24072 31940
rect 23808 31900 23814 31912
rect 24044 31884 24072 31912
rect 22327 31844 22416 31872
rect 22557 31875 22615 31881
rect 22327 31841 22339 31844
rect 22281 31835 22339 31841
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 23934 31872 23940 31884
rect 22603 31844 23940 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 23934 31832 23940 31844
rect 23992 31832 23998 31884
rect 24026 31832 24032 31884
rect 24084 31832 24090 31884
rect 25792 31881 25820 31980
rect 27062 31968 27068 31980
rect 27120 31968 27126 32020
rect 27522 31968 27528 32020
rect 27580 31968 27586 32020
rect 27798 31968 27804 32020
rect 27856 32008 27862 32020
rect 28445 32011 28503 32017
rect 28445 32008 28457 32011
rect 27856 31980 28457 32008
rect 27856 31968 27862 31980
rect 28445 31977 28457 31980
rect 28491 31977 28503 32011
rect 35894 32008 35900 32020
rect 28445 31971 28503 31977
rect 28552 31980 35900 32008
rect 27154 31900 27160 31952
rect 27212 31940 27218 31952
rect 28552 31940 28580 31980
rect 35894 31968 35900 31980
rect 35952 31968 35958 32020
rect 38470 32008 38476 32020
rect 36372 31980 38476 32008
rect 36372 31952 36400 31980
rect 38470 31968 38476 31980
rect 38528 31968 38534 32020
rect 39758 31968 39764 32020
rect 39816 32008 39822 32020
rect 40954 32008 40960 32020
rect 39816 31980 40960 32008
rect 39816 31968 39822 31980
rect 40954 31968 40960 31980
rect 41012 31968 41018 32020
rect 41386 31980 45554 32008
rect 32214 31940 32220 31952
rect 27212 31912 28580 31940
rect 28920 31912 32220 31940
rect 27212 31900 27218 31912
rect 25777 31875 25835 31881
rect 25777 31841 25789 31875
rect 25823 31841 25835 31875
rect 25777 31835 25835 31841
rect 26050 31832 26056 31884
rect 26108 31832 26114 31884
rect 28920 31881 28948 31912
rect 32214 31900 32220 31912
rect 32272 31900 32278 31952
rect 32309 31943 32367 31949
rect 32309 31909 32321 31943
rect 32355 31940 32367 31943
rect 32355 31912 34192 31940
rect 32355 31909 32367 31912
rect 32309 31903 32367 31909
rect 28905 31875 28963 31881
rect 28905 31841 28917 31875
rect 28951 31841 28963 31875
rect 28905 31835 28963 31841
rect 28994 31832 29000 31884
rect 29052 31832 29058 31884
rect 32766 31832 32772 31884
rect 32824 31832 32830 31884
rect 32953 31875 33011 31881
rect 32953 31841 32965 31875
rect 32999 31841 33011 31875
rect 34164 31872 34192 31912
rect 35066 31900 35072 31952
rect 35124 31940 35130 31952
rect 36354 31940 36360 31952
rect 35124 31912 36360 31940
rect 35124 31900 35130 31912
rect 36354 31900 36360 31912
rect 36412 31900 36418 31952
rect 37921 31943 37979 31949
rect 37921 31909 37933 31943
rect 37967 31940 37979 31943
rect 40494 31940 40500 31952
rect 37967 31912 40500 31940
rect 37967 31909 37979 31912
rect 37921 31903 37979 31909
rect 40494 31900 40500 31912
rect 40552 31900 40558 31952
rect 40586 31900 40592 31952
rect 40644 31940 40650 31952
rect 41386 31940 41414 31980
rect 40644 31912 41414 31940
rect 40644 31900 40650 31912
rect 43346 31900 43352 31952
rect 43404 31940 43410 31952
rect 43625 31943 43683 31949
rect 43625 31940 43637 31943
rect 43404 31912 43637 31940
rect 43404 31900 43410 31912
rect 43625 31909 43637 31912
rect 43671 31909 43683 31943
rect 43625 31903 43683 31909
rect 35897 31875 35955 31881
rect 35897 31872 35909 31875
rect 34164 31844 35909 31872
rect 32953 31835 33011 31841
rect 35897 31841 35909 31844
rect 35943 31841 35955 31875
rect 35897 31835 35955 31841
rect 23658 31764 23664 31816
rect 23716 31764 23722 31816
rect 23842 31764 23848 31816
rect 23900 31804 23906 31816
rect 24765 31807 24823 31813
rect 24765 31804 24777 31807
rect 23900 31776 24777 31804
rect 23900 31764 23906 31776
rect 24765 31773 24777 31776
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 27522 31764 27528 31816
rect 27580 31804 27586 31816
rect 31662 31804 31668 31816
rect 27580 31776 31668 31804
rect 27580 31764 27586 31776
rect 31662 31764 31668 31776
rect 31720 31764 31726 31816
rect 32968 31804 32996 31835
rect 36078 31832 36084 31884
rect 36136 31832 36142 31884
rect 37274 31872 37280 31884
rect 36280 31844 37280 31872
rect 34698 31804 34704 31816
rect 32968 31776 34704 31804
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 34974 31764 34980 31816
rect 35032 31804 35038 31816
rect 35710 31804 35716 31816
rect 35032 31776 35716 31804
rect 35032 31764 35038 31776
rect 35710 31764 35716 31776
rect 35768 31804 35774 31816
rect 36280 31804 36308 31844
rect 37274 31832 37280 31844
rect 37332 31832 37338 31884
rect 37458 31832 37464 31884
rect 37516 31872 37522 31884
rect 38470 31872 38476 31884
rect 37516 31844 38476 31872
rect 37516 31832 37522 31844
rect 38470 31832 38476 31844
rect 38528 31832 38534 31884
rect 38580 31844 39804 31872
rect 38580 31804 38608 31844
rect 35768 31776 36308 31804
rect 36372 31776 38608 31804
rect 35768 31764 35774 31776
rect 24854 31696 24860 31748
rect 24912 31736 24918 31748
rect 24912 31708 26464 31736
rect 24912 31696 24918 31708
rect 23198 31628 23204 31680
rect 23256 31668 23262 31680
rect 25682 31668 25688 31680
rect 23256 31640 25688 31668
rect 23256 31628 23262 31640
rect 25682 31628 25688 31640
rect 25740 31628 25746 31680
rect 26436 31668 26464 31708
rect 26510 31696 26516 31748
rect 26568 31696 26574 31748
rect 30282 31736 30288 31748
rect 27632 31708 30288 31736
rect 27632 31668 27660 31708
rect 30282 31696 30288 31708
rect 30340 31696 30346 31748
rect 30374 31696 30380 31748
rect 30432 31736 30438 31748
rect 32677 31739 32735 31745
rect 32677 31736 32689 31739
rect 30432 31708 32689 31736
rect 30432 31696 30438 31708
rect 32677 31705 32689 31708
rect 32723 31705 32735 31739
rect 32677 31699 32735 31705
rect 35618 31696 35624 31748
rect 35676 31736 35682 31748
rect 36372 31736 36400 31776
rect 39298 31764 39304 31816
rect 39356 31804 39362 31816
rect 39485 31807 39543 31813
rect 39485 31804 39497 31807
rect 39356 31776 39497 31804
rect 39356 31764 39362 31776
rect 39485 31773 39497 31776
rect 39531 31773 39543 31807
rect 39485 31767 39543 31773
rect 35676 31708 36400 31736
rect 38381 31739 38439 31745
rect 35676 31696 35682 31708
rect 38381 31705 38393 31739
rect 38427 31736 38439 31739
rect 38654 31736 38660 31748
rect 38427 31708 38660 31736
rect 38427 31705 38439 31708
rect 38381 31699 38439 31705
rect 38654 31696 38660 31708
rect 38712 31696 38718 31748
rect 26436 31640 27660 31668
rect 27706 31628 27712 31680
rect 27764 31668 27770 31680
rect 28718 31668 28724 31680
rect 27764 31640 28724 31668
rect 27764 31628 27770 31640
rect 28718 31628 28724 31640
rect 28776 31668 28782 31680
rect 28813 31671 28871 31677
rect 28813 31668 28825 31671
rect 28776 31640 28825 31668
rect 28776 31628 28782 31640
rect 28813 31637 28825 31640
rect 28859 31637 28871 31671
rect 28813 31631 28871 31637
rect 35434 31628 35440 31680
rect 35492 31628 35498 31680
rect 35805 31671 35863 31677
rect 35805 31637 35817 31671
rect 35851 31668 35863 31671
rect 37090 31668 37096 31680
rect 35851 31640 37096 31668
rect 35851 31637 35863 31640
rect 35805 31631 35863 31637
rect 37090 31628 37096 31640
rect 37148 31628 37154 31680
rect 37366 31628 37372 31680
rect 37424 31668 37430 31680
rect 37918 31668 37924 31680
rect 37424 31640 37924 31668
rect 37424 31628 37430 31640
rect 37918 31628 37924 31640
rect 37976 31668 37982 31680
rect 38289 31671 38347 31677
rect 38289 31668 38301 31671
rect 37976 31640 38301 31668
rect 37976 31628 37982 31640
rect 38289 31637 38301 31640
rect 38335 31637 38347 31671
rect 38289 31631 38347 31637
rect 39301 31671 39359 31677
rect 39301 31637 39313 31671
rect 39347 31668 39359 31671
rect 39666 31668 39672 31680
rect 39347 31640 39672 31668
rect 39347 31637 39359 31640
rect 39301 31631 39359 31637
rect 39666 31628 39672 31640
rect 39724 31628 39730 31680
rect 39776 31668 39804 31844
rect 40310 31832 40316 31884
rect 40368 31872 40374 31884
rect 41877 31875 41935 31881
rect 41877 31872 41889 31875
rect 40368 31844 41889 31872
rect 40368 31832 40374 31844
rect 41877 31841 41889 31844
rect 41923 31841 41935 31875
rect 41877 31835 41935 31841
rect 42153 31875 42211 31881
rect 42153 31841 42165 31875
rect 42199 31872 42211 31875
rect 42702 31872 42708 31884
rect 42199 31844 42708 31872
rect 42199 31841 42211 31844
rect 42153 31835 42211 31841
rect 42702 31832 42708 31844
rect 42760 31832 42766 31884
rect 45526 31872 45554 31980
rect 48777 31875 48835 31881
rect 48777 31872 48789 31875
rect 45526 31844 48789 31872
rect 48777 31841 48789 31844
rect 48823 31841 48835 31875
rect 48777 31835 48835 31841
rect 48041 31807 48099 31813
rect 48041 31773 48053 31807
rect 48087 31804 48099 31807
rect 48498 31804 48504 31816
rect 48087 31776 48504 31804
rect 48087 31773 48099 31776
rect 48041 31767 48099 31773
rect 48498 31764 48504 31776
rect 48556 31764 48562 31816
rect 42610 31696 42616 31748
rect 42668 31696 42674 31748
rect 41782 31668 41788 31680
rect 39776 31640 41788 31668
rect 41782 31628 41788 31640
rect 41840 31668 41846 31680
rect 42242 31668 42248 31680
rect 41840 31640 42248 31668
rect 41840 31628 41846 31640
rect 42242 31628 42248 31640
rect 42300 31628 42306 31680
rect 1104 31578 49864 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 27950 31578
rect 28002 31526 28014 31578
rect 28066 31526 28078 31578
rect 28130 31526 28142 31578
rect 28194 31526 28206 31578
rect 28258 31526 37950 31578
rect 38002 31526 38014 31578
rect 38066 31526 38078 31578
rect 38130 31526 38142 31578
rect 38194 31526 38206 31578
rect 38258 31526 47950 31578
rect 48002 31526 48014 31578
rect 48066 31526 48078 31578
rect 48130 31526 48142 31578
rect 48194 31526 48206 31578
rect 48258 31526 49864 31578
rect 1104 31504 49864 31526
rect 23842 31424 23848 31476
rect 23900 31424 23906 31476
rect 23934 31424 23940 31476
rect 23992 31464 23998 31476
rect 26605 31467 26663 31473
rect 26605 31464 26617 31467
rect 23992 31436 26617 31464
rect 23992 31424 23998 31436
rect 26605 31433 26617 31436
rect 26651 31464 26663 31467
rect 28902 31464 28908 31476
rect 26651 31436 28908 31464
rect 26651 31433 26663 31436
rect 26605 31427 26663 31433
rect 28902 31424 28908 31436
rect 28960 31424 28966 31476
rect 36262 31464 36268 31476
rect 34532 31436 36268 31464
rect 23474 31356 23480 31408
rect 23532 31396 23538 31408
rect 24762 31396 24768 31408
rect 23532 31368 24768 31396
rect 23532 31356 23538 31368
rect 24762 31356 24768 31368
rect 24820 31396 24826 31408
rect 24820 31368 24900 31396
rect 24820 31356 24826 31368
rect 22373 31331 22431 31337
rect 22373 31297 22385 31331
rect 22419 31328 22431 31331
rect 22830 31328 22836 31340
rect 22419 31300 22836 31328
rect 22419 31297 22431 31300
rect 22373 31291 22431 31297
rect 22830 31288 22836 31300
rect 22888 31288 22894 31340
rect 23290 31288 23296 31340
rect 23348 31328 23354 31340
rect 24872 31337 24900 31368
rect 23937 31331 23995 31337
rect 23937 31328 23949 31331
rect 23348 31300 23949 31328
rect 23348 31288 23354 31300
rect 23937 31297 23949 31300
rect 23983 31297 23995 31331
rect 23937 31291 23995 31297
rect 24857 31331 24915 31337
rect 24857 31297 24869 31331
rect 24903 31297 24915 31331
rect 24857 31291 24915 31297
rect 26234 31288 26240 31340
rect 26292 31328 26298 31340
rect 26510 31328 26516 31340
rect 26292 31300 26516 31328
rect 26292 31288 26298 31300
rect 26510 31288 26516 31300
rect 26568 31288 26574 31340
rect 27154 31288 27160 31340
rect 27212 31328 27218 31340
rect 33321 31331 33379 31337
rect 33321 31328 33333 31331
rect 27212 31300 33333 31328
rect 27212 31288 27218 31300
rect 33321 31297 33333 31300
rect 33367 31297 33379 31331
rect 33321 31291 33379 31297
rect 33413 31331 33471 31337
rect 33413 31297 33425 31331
rect 33459 31328 33471 31331
rect 33870 31328 33876 31340
rect 33459 31300 33876 31328
rect 33459 31297 33471 31300
rect 33413 31291 33471 31297
rect 33870 31288 33876 31300
rect 33928 31288 33934 31340
rect 34532 31337 34560 31436
rect 36262 31424 36268 31436
rect 36320 31424 36326 31476
rect 39298 31464 39304 31476
rect 38764 31436 39304 31464
rect 35802 31356 35808 31408
rect 35860 31356 35866 31408
rect 36538 31356 36544 31408
rect 36596 31396 36602 31408
rect 38194 31396 38200 31408
rect 36596 31368 38200 31396
rect 36596 31356 36602 31368
rect 38194 31356 38200 31368
rect 38252 31356 38258 31408
rect 38657 31399 38715 31405
rect 38657 31365 38669 31399
rect 38703 31396 38715 31399
rect 38764 31396 38792 31436
rect 39298 31424 39304 31436
rect 39356 31464 39362 31476
rect 39482 31464 39488 31476
rect 39356 31436 39488 31464
rect 39356 31424 39362 31436
rect 39482 31424 39488 31436
rect 39540 31424 39546 31476
rect 42794 31424 42800 31476
rect 42852 31464 42858 31476
rect 42981 31467 43039 31473
rect 42981 31464 42993 31467
rect 42852 31436 42993 31464
rect 42852 31424 42858 31436
rect 42981 31433 42993 31436
rect 43027 31433 43039 31467
rect 42981 31427 43039 31433
rect 47854 31424 47860 31476
rect 47912 31464 47918 31476
rect 47949 31467 48007 31473
rect 47949 31464 47961 31467
rect 47912 31436 47961 31464
rect 47912 31424 47918 31436
rect 47949 31433 47961 31436
rect 47995 31433 48007 31467
rect 47949 31427 48007 31433
rect 38703 31368 38792 31396
rect 38703 31365 38715 31368
rect 38657 31359 38715 31365
rect 42426 31356 42432 31408
rect 42484 31396 42490 31408
rect 43073 31399 43131 31405
rect 43073 31396 43085 31399
rect 42484 31368 43085 31396
rect 42484 31356 42490 31368
rect 43073 31365 43085 31368
rect 43119 31396 43131 31399
rect 45738 31396 45744 31408
rect 43119 31368 45744 31396
rect 43119 31365 43131 31368
rect 43073 31359 43131 31365
rect 45738 31356 45744 31368
rect 45796 31356 45802 31408
rect 34517 31331 34575 31337
rect 34517 31297 34529 31331
rect 34563 31297 34575 31331
rect 34517 31291 34575 31297
rect 37734 31288 37740 31340
rect 37792 31288 37798 31340
rect 38378 31288 38384 31340
rect 38436 31328 38442 31340
rect 38565 31331 38623 31337
rect 38565 31328 38577 31331
rect 38436 31300 38577 31328
rect 38436 31288 38442 31300
rect 38565 31297 38577 31300
rect 38611 31297 38623 31331
rect 38565 31291 38623 31297
rect 38764 31300 38976 31328
rect 22462 31220 22468 31272
rect 22520 31220 22526 31272
rect 22649 31263 22707 31269
rect 22649 31229 22661 31263
rect 22695 31260 22707 31263
rect 22695 31232 23428 31260
rect 22695 31229 22707 31232
rect 22649 31223 22707 31229
rect 21453 31127 21511 31133
rect 21453 31093 21465 31127
rect 21499 31124 21511 31127
rect 21818 31124 21824 31136
rect 21499 31096 21824 31124
rect 21499 31093 21511 31096
rect 21453 31087 21511 31093
rect 21818 31084 21824 31096
rect 21876 31084 21882 31136
rect 22005 31127 22063 31133
rect 22005 31093 22017 31127
rect 22051 31124 22063 31127
rect 23198 31124 23204 31136
rect 22051 31096 23204 31124
rect 22051 31093 22063 31096
rect 22005 31087 22063 31093
rect 23198 31084 23204 31096
rect 23256 31084 23262 31136
rect 23400 31124 23428 31232
rect 24118 31220 24124 31272
rect 24176 31220 24182 31272
rect 24578 31220 24584 31272
rect 24636 31260 24642 31272
rect 25133 31263 25191 31269
rect 25133 31260 25145 31263
rect 24636 31232 25145 31260
rect 24636 31220 24642 31232
rect 25133 31229 25145 31232
rect 25179 31260 25191 31263
rect 27522 31260 27528 31272
rect 25179 31232 27528 31260
rect 25179 31229 25191 31232
rect 25133 31223 25191 31229
rect 27522 31220 27528 31232
rect 27580 31220 27586 31272
rect 31662 31220 31668 31272
rect 31720 31260 31726 31272
rect 33597 31263 33655 31269
rect 33597 31260 33609 31263
rect 31720 31232 33364 31260
rect 31720 31220 31726 31232
rect 23477 31195 23535 31201
rect 23477 31161 23489 31195
rect 23523 31192 23535 31195
rect 24670 31192 24676 31204
rect 23523 31164 24676 31192
rect 23523 31161 23535 31164
rect 23477 31155 23535 31161
rect 24670 31152 24676 31164
rect 24728 31152 24734 31204
rect 24946 31124 24952 31136
rect 23400 31096 24952 31124
rect 24946 31084 24952 31096
rect 25004 31084 25010 31136
rect 25774 31084 25780 31136
rect 25832 31124 25838 31136
rect 30374 31124 30380 31136
rect 25832 31096 30380 31124
rect 25832 31084 25838 31096
rect 30374 31084 30380 31096
rect 30432 31084 30438 31136
rect 32858 31084 32864 31136
rect 32916 31124 32922 31136
rect 32953 31127 33011 31133
rect 32953 31124 32965 31127
rect 32916 31096 32965 31124
rect 32916 31084 32922 31096
rect 32953 31093 32965 31096
rect 32999 31093 33011 31127
rect 33336 31124 33364 31232
rect 33428 31232 33609 31260
rect 33428 31204 33456 31232
rect 33597 31229 33609 31232
rect 33643 31260 33655 31263
rect 34054 31260 34060 31272
rect 33643 31232 34060 31260
rect 33643 31229 33655 31232
rect 33597 31223 33655 31229
rect 34054 31220 34060 31232
rect 34112 31220 34118 31272
rect 34793 31263 34851 31269
rect 34793 31229 34805 31263
rect 34839 31260 34851 31263
rect 35526 31260 35532 31272
rect 34839 31232 35532 31260
rect 34839 31229 34851 31232
rect 34793 31223 34851 31229
rect 35526 31220 35532 31232
rect 35584 31220 35590 31272
rect 36265 31263 36323 31269
rect 36265 31229 36277 31263
rect 36311 31260 36323 31263
rect 36354 31260 36360 31272
rect 36311 31232 36360 31260
rect 36311 31229 36323 31232
rect 36265 31223 36323 31229
rect 36354 31220 36360 31232
rect 36412 31220 36418 31272
rect 36446 31220 36452 31272
rect 36504 31260 36510 31272
rect 38764 31260 38792 31300
rect 36504 31232 38792 31260
rect 38841 31263 38899 31269
rect 36504 31220 36510 31232
rect 38841 31229 38853 31263
rect 38887 31229 38899 31263
rect 38948 31260 38976 31300
rect 39022 31288 39028 31340
rect 39080 31328 39086 31340
rect 40865 31331 40923 31337
rect 40865 31328 40877 31331
rect 39080 31300 40877 31328
rect 39080 31288 39086 31300
rect 40865 31297 40877 31300
rect 40911 31297 40923 31331
rect 40865 31291 40923 31297
rect 42058 31288 42064 31340
rect 42116 31328 42122 31340
rect 42116 31300 43208 31328
rect 42116 31288 42122 31300
rect 42150 31260 42156 31272
rect 38948 31232 42156 31260
rect 38841 31223 38899 31229
rect 33410 31152 33416 31204
rect 33468 31152 33474 31204
rect 38470 31152 38476 31204
rect 38528 31192 38534 31204
rect 38856 31192 38884 31223
rect 42150 31220 42156 31232
rect 42208 31220 42214 31272
rect 43180 31269 43208 31300
rect 44266 31288 44272 31340
rect 44324 31328 44330 31340
rect 45649 31331 45707 31337
rect 45649 31328 45661 31331
rect 44324 31300 45661 31328
rect 44324 31288 44330 31300
rect 45649 31297 45661 31300
rect 45695 31297 45707 31331
rect 45649 31291 45707 31297
rect 47394 31288 47400 31340
rect 47452 31328 47458 31340
rect 47857 31331 47915 31337
rect 47857 31328 47869 31331
rect 47452 31300 47869 31328
rect 47452 31288 47458 31300
rect 47857 31297 47869 31300
rect 47903 31297 47915 31331
rect 48777 31331 48835 31337
rect 48777 31328 48789 31331
rect 47857 31291 47915 31297
rect 47964 31300 48789 31328
rect 43165 31263 43223 31269
rect 43165 31229 43177 31263
rect 43211 31229 43223 31263
rect 43165 31223 43223 31229
rect 44358 31220 44364 31272
rect 44416 31260 44422 31272
rect 47964 31260 47992 31300
rect 48777 31297 48789 31300
rect 48823 31297 48835 31331
rect 48777 31291 48835 31297
rect 44416 31232 47992 31260
rect 44416 31220 44422 31232
rect 48498 31220 48504 31272
rect 48556 31220 48562 31272
rect 38528 31164 38884 31192
rect 40681 31195 40739 31201
rect 38528 31152 38534 31164
rect 40681 31161 40693 31195
rect 40727 31192 40739 31195
rect 46014 31192 46020 31204
rect 40727 31164 46020 31192
rect 40727 31161 40739 31164
rect 40681 31155 40739 31161
rect 46014 31152 46020 31164
rect 46072 31152 46078 31204
rect 36998 31124 37004 31136
rect 33336 31096 37004 31124
rect 32953 31087 33011 31093
rect 36998 31084 37004 31096
rect 37056 31084 37062 31136
rect 37550 31084 37556 31136
rect 37608 31084 37614 31136
rect 38197 31127 38255 31133
rect 38197 31093 38209 31127
rect 38243 31124 38255 31127
rect 40402 31124 40408 31136
rect 38243 31096 40408 31124
rect 38243 31093 38255 31096
rect 38197 31087 38255 31093
rect 40402 31084 40408 31096
rect 40460 31084 40466 31136
rect 40770 31084 40776 31136
rect 40828 31124 40834 31136
rect 42613 31127 42671 31133
rect 42613 31124 42625 31127
rect 40828 31096 42625 31124
rect 40828 31084 40834 31096
rect 42613 31093 42625 31096
rect 42659 31093 42671 31127
rect 42613 31087 42671 31093
rect 45465 31127 45523 31133
rect 45465 31093 45477 31127
rect 45511 31124 45523 31127
rect 46934 31124 46940 31136
rect 45511 31096 46940 31124
rect 45511 31093 45523 31096
rect 45465 31087 45523 31093
rect 46934 31084 46940 31096
rect 46992 31084 46998 31136
rect 1104 31034 49864 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 32950 31034
rect 33002 30982 33014 31034
rect 33066 30982 33078 31034
rect 33130 30982 33142 31034
rect 33194 30982 33206 31034
rect 33258 30982 42950 31034
rect 43002 30982 43014 31034
rect 43066 30982 43078 31034
rect 43130 30982 43142 31034
rect 43194 30982 43206 31034
rect 43258 30982 49864 31034
rect 1104 30960 49864 30982
rect 22738 30880 22744 30932
rect 22796 30920 22802 30932
rect 23293 30923 23351 30929
rect 23293 30920 23305 30923
rect 22796 30892 23305 30920
rect 22796 30880 22802 30892
rect 23293 30889 23305 30892
rect 23339 30889 23351 30923
rect 25130 30920 25136 30932
rect 23293 30883 23351 30889
rect 23584 30892 25136 30920
rect 21453 30855 21511 30861
rect 21453 30821 21465 30855
rect 21499 30852 21511 30855
rect 21499 30824 22784 30852
rect 21499 30821 21511 30824
rect 21453 30815 21511 30821
rect 22094 30744 22100 30796
rect 22152 30744 22158 30796
rect 22756 30784 22784 30824
rect 22830 30812 22836 30864
rect 22888 30812 22894 30864
rect 23584 30784 23612 30892
rect 25130 30880 25136 30892
rect 25188 30880 25194 30932
rect 26605 30923 26663 30929
rect 26605 30889 26617 30923
rect 26651 30920 26663 30923
rect 28350 30920 28356 30932
rect 26651 30892 28356 30920
rect 26651 30889 26663 30892
rect 26605 30883 26663 30889
rect 24118 30812 24124 30864
rect 24176 30852 24182 30864
rect 24176 30824 24992 30852
rect 24176 30812 24182 30824
rect 22756 30756 23612 30784
rect 23934 30744 23940 30796
rect 23992 30744 23998 30796
rect 24762 30744 24768 30796
rect 24820 30784 24826 30796
rect 24857 30787 24915 30793
rect 24857 30784 24869 30787
rect 24820 30756 24869 30784
rect 24820 30744 24826 30756
rect 24857 30753 24869 30756
rect 24903 30753 24915 30787
rect 24964 30784 24992 30824
rect 26620 30784 26648 30883
rect 28350 30880 28356 30892
rect 28408 30880 28414 30932
rect 30944 30892 34560 30920
rect 30944 30861 30972 30892
rect 30929 30855 30987 30861
rect 30929 30852 30941 30855
rect 24964 30756 26648 30784
rect 26988 30824 27200 30852
rect 24857 30747 24915 30753
rect 21818 30676 21824 30728
rect 21876 30676 21882 30728
rect 23382 30676 23388 30728
rect 23440 30716 23446 30728
rect 24578 30716 24584 30728
rect 23440 30688 24584 30716
rect 23440 30676 23446 30688
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 26234 30676 26240 30728
rect 26292 30716 26298 30728
rect 26988 30716 27016 30824
rect 27062 30744 27068 30796
rect 27120 30744 27126 30796
rect 27172 30784 27200 30824
rect 30208 30824 30941 30852
rect 27172 30756 28488 30784
rect 26292 30688 27016 30716
rect 28460 30702 28488 30756
rect 30208 30725 30236 30824
rect 30929 30821 30941 30824
rect 30975 30821 30987 30855
rect 30929 30815 30987 30821
rect 30282 30744 30288 30796
rect 30340 30744 30346 30796
rect 32122 30784 32128 30796
rect 31312 30756 32128 30784
rect 31312 30728 31340 30756
rect 32122 30744 32128 30756
rect 32180 30784 32186 30796
rect 32306 30784 32312 30796
rect 32180 30756 32312 30784
rect 32180 30744 32186 30756
rect 32306 30744 32312 30756
rect 32364 30744 32370 30796
rect 34532 30784 34560 30892
rect 36170 30880 36176 30932
rect 36228 30920 36234 30932
rect 36228 30892 39436 30920
rect 36228 30880 36234 30892
rect 35894 30852 35900 30864
rect 35544 30824 35900 30852
rect 35437 30787 35495 30793
rect 34532 30756 35388 30784
rect 30193 30719 30251 30725
rect 30193 30716 30205 30719
rect 28736 30688 30205 30716
rect 26292 30676 26298 30688
rect 22186 30608 22192 30660
rect 22244 30648 22250 30660
rect 23753 30651 23811 30657
rect 23753 30648 23765 30651
rect 22244 30620 23765 30648
rect 22244 30608 22250 30620
rect 23753 30617 23765 30620
rect 23799 30617 23811 30651
rect 23753 30611 23811 30617
rect 24854 30608 24860 30660
rect 24912 30648 24918 30660
rect 25130 30648 25136 30660
rect 24912 30620 25136 30648
rect 24912 30608 24918 30620
rect 25130 30608 25136 30620
rect 25188 30608 25194 30660
rect 27338 30608 27344 30660
rect 27396 30608 27402 30660
rect 9214 30540 9220 30592
rect 9272 30580 9278 30592
rect 20901 30583 20959 30589
rect 20901 30580 20913 30583
rect 9272 30552 20913 30580
rect 9272 30540 9278 30552
rect 20901 30549 20913 30552
rect 20947 30580 20959 30583
rect 21818 30580 21824 30592
rect 20947 30552 21824 30580
rect 20947 30549 20959 30552
rect 20901 30543 20959 30549
rect 21818 30540 21824 30552
rect 21876 30580 21882 30592
rect 21913 30583 21971 30589
rect 21913 30580 21925 30583
rect 21876 30552 21925 30580
rect 21876 30540 21882 30552
rect 21913 30549 21925 30552
rect 21959 30549 21971 30583
rect 21913 30543 21971 30549
rect 23566 30540 23572 30592
rect 23624 30580 23630 30592
rect 23661 30583 23719 30589
rect 23661 30580 23673 30583
rect 23624 30552 23673 30580
rect 23624 30540 23630 30552
rect 23661 30549 23673 30552
rect 23707 30549 23719 30583
rect 23661 30543 23719 30549
rect 25406 30540 25412 30592
rect 25464 30580 25470 30592
rect 28736 30580 28764 30688
rect 30193 30685 30205 30688
rect 30239 30685 30251 30719
rect 30193 30679 30251 30685
rect 30374 30676 30380 30728
rect 30432 30716 30438 30728
rect 30432 30688 31156 30716
rect 30432 30676 30438 30688
rect 30101 30651 30159 30657
rect 30101 30617 30113 30651
rect 30147 30648 30159 30651
rect 31128 30648 31156 30688
rect 31294 30676 31300 30728
rect 31352 30676 31358 30728
rect 34790 30676 34796 30728
rect 34848 30716 34854 30728
rect 34974 30716 34980 30728
rect 34848 30688 34980 30716
rect 34848 30676 34854 30688
rect 34974 30676 34980 30688
rect 35032 30676 35038 30728
rect 35360 30725 35388 30756
rect 35437 30753 35449 30787
rect 35483 30784 35495 30787
rect 35544 30784 35572 30824
rect 35894 30812 35900 30824
rect 35952 30812 35958 30864
rect 35986 30812 35992 30864
rect 36044 30852 36050 30864
rect 36357 30855 36415 30861
rect 36357 30852 36369 30855
rect 36044 30824 36369 30852
rect 36044 30812 36050 30824
rect 36357 30821 36369 30824
rect 36403 30821 36415 30855
rect 36357 30815 36415 30821
rect 36538 30812 36544 30864
rect 36596 30852 36602 30864
rect 38930 30852 38936 30864
rect 36596 30824 38936 30852
rect 36596 30812 36602 30824
rect 38930 30812 38936 30824
rect 38988 30812 38994 30864
rect 39408 30852 39436 30892
rect 39482 30880 39488 30932
rect 39540 30920 39546 30932
rect 41874 30920 41880 30932
rect 39540 30892 41880 30920
rect 39540 30880 39546 30892
rect 41874 30880 41880 30892
rect 41932 30880 41938 30932
rect 47670 30880 47676 30932
rect 47728 30920 47734 30932
rect 48777 30923 48835 30929
rect 48777 30920 48789 30923
rect 47728 30892 48789 30920
rect 47728 30880 47734 30892
rect 48777 30889 48789 30892
rect 48823 30889 48835 30923
rect 48777 30883 48835 30889
rect 39408 30824 40724 30852
rect 35483 30756 35572 30784
rect 35621 30787 35679 30793
rect 35483 30753 35495 30756
rect 35437 30747 35495 30753
rect 35621 30753 35633 30787
rect 35667 30784 35679 30787
rect 35710 30784 35716 30796
rect 35667 30756 35716 30784
rect 35667 30753 35679 30756
rect 35621 30747 35679 30753
rect 35710 30744 35716 30756
rect 35768 30744 35774 30796
rect 36906 30744 36912 30796
rect 36964 30744 36970 30796
rect 36998 30744 37004 30796
rect 37056 30784 37062 30796
rect 37921 30787 37979 30793
rect 37921 30784 37933 30787
rect 37056 30756 37933 30784
rect 37056 30744 37062 30756
rect 37921 30753 37933 30756
rect 37967 30753 37979 30787
rect 37921 30747 37979 30753
rect 38746 30744 38752 30796
rect 38804 30784 38810 30796
rect 39117 30787 39175 30793
rect 39117 30784 39129 30787
rect 38804 30756 39129 30784
rect 38804 30744 38810 30756
rect 39117 30753 39129 30756
rect 39163 30753 39175 30787
rect 39117 30747 39175 30753
rect 39209 30787 39267 30793
rect 39209 30753 39221 30787
rect 39255 30784 39267 30787
rect 39390 30784 39396 30796
rect 39255 30756 39396 30784
rect 39255 30753 39267 30756
rect 39209 30747 39267 30753
rect 39390 30744 39396 30756
rect 39448 30744 39454 30796
rect 40494 30744 40500 30796
rect 40552 30744 40558 30796
rect 40586 30744 40592 30796
rect 40644 30744 40650 30796
rect 35345 30719 35403 30725
rect 35345 30685 35357 30719
rect 35391 30716 35403 30719
rect 36173 30719 36231 30725
rect 36173 30716 36185 30719
rect 35391 30688 36185 30716
rect 35391 30685 35403 30688
rect 35345 30679 35403 30685
rect 36173 30685 36185 30688
rect 36219 30685 36231 30719
rect 36173 30679 36231 30685
rect 36817 30719 36875 30725
rect 36817 30685 36829 30719
rect 36863 30716 36875 30719
rect 39025 30719 39083 30725
rect 39025 30716 39037 30719
rect 36863 30688 39037 30716
rect 36863 30685 36875 30688
rect 36817 30679 36875 30685
rect 39025 30685 39037 30688
rect 39071 30716 39083 30719
rect 39482 30716 39488 30728
rect 39071 30688 39488 30716
rect 39071 30685 39083 30688
rect 39025 30679 39083 30685
rect 39482 30676 39488 30688
rect 39540 30676 39546 30728
rect 40402 30676 40408 30728
rect 40460 30676 40466 30728
rect 40696 30716 40724 30824
rect 41506 30812 41512 30864
rect 41564 30812 41570 30864
rect 41524 30784 41552 30812
rect 41524 30756 43300 30784
rect 41509 30719 41567 30725
rect 41509 30716 41521 30719
rect 40696 30688 41521 30716
rect 41509 30685 41521 30688
rect 41555 30685 41567 30719
rect 41509 30679 41567 30685
rect 42150 30676 42156 30728
rect 42208 30676 42214 30728
rect 43272 30725 43300 30756
rect 43257 30719 43315 30725
rect 43257 30685 43269 30719
rect 43303 30685 43315 30719
rect 43257 30679 43315 30685
rect 31570 30648 31576 30660
rect 30147 30620 31064 30648
rect 31128 30620 31576 30648
rect 30147 30617 30159 30620
rect 30101 30611 30159 30617
rect 25464 30552 28764 30580
rect 25464 30540 25470 30552
rect 28810 30540 28816 30592
rect 28868 30540 28874 30592
rect 28902 30540 28908 30592
rect 28960 30580 28966 30592
rect 29733 30583 29791 30589
rect 29733 30580 29745 30583
rect 28960 30552 29745 30580
rect 28960 30540 28966 30552
rect 29733 30549 29745 30552
rect 29779 30549 29791 30583
rect 31036 30580 31064 30620
rect 31570 30608 31576 30620
rect 31628 30608 31634 30660
rect 32798 30620 34284 30648
rect 32398 30580 32404 30592
rect 31036 30552 32404 30580
rect 29733 30543 29791 30549
rect 32398 30540 32404 30552
rect 32456 30540 32462 30592
rect 32582 30540 32588 30592
rect 32640 30580 32646 30592
rect 33045 30583 33103 30589
rect 33045 30580 33057 30583
rect 32640 30552 33057 30580
rect 32640 30540 32646 30552
rect 33045 30549 33057 30552
rect 33091 30549 33103 30583
rect 34256 30580 34284 30620
rect 34606 30608 34612 30660
rect 34664 30648 34670 30660
rect 37829 30651 37887 30657
rect 34664 30620 37412 30648
rect 34664 30608 34670 30620
rect 34790 30580 34796 30592
rect 34256 30552 34796 30580
rect 33045 30543 33103 30549
rect 34790 30540 34796 30552
rect 34848 30540 34854 30592
rect 34977 30583 35035 30589
rect 34977 30549 34989 30583
rect 35023 30580 35035 30583
rect 36538 30580 36544 30592
rect 35023 30552 36544 30580
rect 35023 30549 35035 30552
rect 34977 30543 35035 30549
rect 36538 30540 36544 30552
rect 36596 30540 36602 30592
rect 36725 30583 36783 30589
rect 36725 30549 36737 30583
rect 36771 30580 36783 30583
rect 37090 30580 37096 30592
rect 36771 30552 37096 30580
rect 36771 30549 36783 30552
rect 36725 30543 36783 30549
rect 37090 30540 37096 30552
rect 37148 30540 37154 30592
rect 37384 30589 37412 30620
rect 37829 30617 37841 30651
rect 37875 30648 37887 30651
rect 41230 30648 41236 30660
rect 37875 30620 41236 30648
rect 37875 30617 37887 30620
rect 37829 30611 37887 30617
rect 41230 30608 41236 30620
rect 41288 30608 41294 30660
rect 46106 30648 46112 30660
rect 41340 30620 46112 30648
rect 37369 30583 37427 30589
rect 37369 30549 37381 30583
rect 37415 30549 37427 30583
rect 37369 30543 37427 30549
rect 37734 30540 37740 30592
rect 37792 30540 37798 30592
rect 38657 30583 38715 30589
rect 38657 30549 38669 30583
rect 38703 30580 38715 30583
rect 38746 30580 38752 30592
rect 38703 30552 38752 30580
rect 38703 30549 38715 30552
rect 38657 30543 38715 30549
rect 38746 30540 38752 30552
rect 38804 30540 38810 30592
rect 40034 30540 40040 30592
rect 40092 30540 40098 30592
rect 41340 30589 41368 30620
rect 46106 30608 46112 30620
rect 46164 30608 46170 30660
rect 48682 30608 48688 30660
rect 48740 30608 48746 30660
rect 41325 30583 41383 30589
rect 41325 30549 41337 30583
rect 41371 30549 41383 30583
rect 41325 30543 41383 30549
rect 41966 30540 41972 30592
rect 42024 30540 42030 30592
rect 43073 30583 43131 30589
rect 43073 30549 43085 30583
rect 43119 30580 43131 30583
rect 47026 30580 47032 30592
rect 43119 30552 47032 30580
rect 43119 30549 43131 30552
rect 43073 30543 43131 30549
rect 47026 30540 47032 30552
rect 47084 30540 47090 30592
rect 1104 30490 49864 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 27950 30490
rect 28002 30438 28014 30490
rect 28066 30438 28078 30490
rect 28130 30438 28142 30490
rect 28194 30438 28206 30490
rect 28258 30438 37950 30490
rect 38002 30438 38014 30490
rect 38066 30438 38078 30490
rect 38130 30438 38142 30490
rect 38194 30438 38206 30490
rect 38258 30438 47950 30490
rect 48002 30438 48014 30490
rect 48066 30438 48078 30490
rect 48130 30438 48142 30490
rect 48194 30438 48206 30490
rect 48258 30438 49864 30490
rect 1104 30416 49864 30438
rect 28721 30379 28779 30385
rect 28721 30376 28733 30379
rect 28644 30348 28733 30376
rect 24489 30311 24547 30317
rect 24489 30277 24501 30311
rect 24535 30308 24547 30311
rect 24762 30308 24768 30320
rect 24535 30280 24768 30308
rect 24535 30277 24547 30280
rect 24489 30271 24547 30277
rect 24762 30268 24768 30280
rect 24820 30268 24826 30320
rect 26050 30268 26056 30320
rect 26108 30268 26114 30320
rect 7374 30200 7380 30252
rect 7432 30200 7438 30252
rect 21174 30200 21180 30252
rect 21232 30240 21238 30252
rect 23661 30243 23719 30249
rect 23661 30240 23673 30243
rect 21232 30212 23673 30240
rect 21232 30200 21238 30212
rect 23661 30209 23673 30212
rect 23707 30240 23719 30243
rect 25498 30240 25504 30252
rect 23707 30212 25504 30240
rect 23707 30209 23719 30212
rect 23661 30203 23719 30209
rect 25498 30200 25504 30212
rect 25556 30200 25562 30252
rect 25590 30200 25596 30252
rect 25648 30240 25654 30252
rect 25961 30243 26019 30249
rect 25961 30240 25973 30243
rect 25648 30212 25973 30240
rect 25648 30200 25654 30212
rect 25961 30209 25973 30212
rect 26007 30209 26019 30243
rect 25961 30203 26019 30209
rect 7561 30175 7619 30181
rect 7561 30141 7573 30175
rect 7607 30172 7619 30175
rect 7650 30172 7656 30184
rect 7607 30144 7656 30172
rect 7607 30141 7619 30144
rect 7561 30135 7619 30141
rect 7650 30132 7656 30144
rect 7708 30132 7714 30184
rect 9122 30132 9128 30184
rect 9180 30132 9186 30184
rect 23566 30132 23572 30184
rect 23624 30132 23630 30184
rect 25133 30175 25191 30181
rect 25133 30141 25145 30175
rect 25179 30172 25191 30175
rect 25608 30172 25636 30200
rect 25179 30144 25636 30172
rect 26145 30175 26203 30181
rect 25179 30141 25191 30144
rect 25133 30135 25191 30141
rect 26145 30141 26157 30175
rect 26191 30172 26203 30175
rect 27522 30172 27528 30184
rect 26191 30144 27528 30172
rect 26191 30141 26203 30144
rect 26145 30135 26203 30141
rect 27522 30132 27528 30144
rect 27580 30132 27586 30184
rect 28644 30172 28672 30348
rect 28721 30345 28733 30348
rect 28767 30376 28779 30379
rect 28767 30348 29132 30376
rect 28767 30345 28779 30348
rect 28721 30339 28779 30345
rect 28718 30200 28724 30252
rect 28776 30240 28782 30252
rect 29104 30240 29132 30348
rect 30466 30336 30472 30388
rect 30524 30376 30530 30388
rect 36906 30376 36912 30388
rect 30524 30348 36912 30376
rect 30524 30336 30530 30348
rect 36906 30336 36912 30348
rect 36964 30336 36970 30388
rect 37458 30336 37464 30388
rect 37516 30376 37522 30388
rect 38378 30376 38384 30388
rect 37516 30348 38384 30376
rect 37516 30336 37522 30348
rect 38378 30336 38384 30348
rect 38436 30336 38442 30388
rect 41230 30336 41236 30388
rect 41288 30376 41294 30388
rect 41325 30379 41383 30385
rect 41325 30376 41337 30379
rect 41288 30348 41337 30376
rect 41288 30336 41294 30348
rect 41325 30345 41337 30348
rect 41371 30345 41383 30379
rect 41325 30339 41383 30345
rect 30006 30268 30012 30320
rect 30064 30308 30070 30320
rect 31294 30308 31300 30320
rect 30064 30280 31300 30308
rect 30064 30268 30070 30280
rect 31294 30268 31300 30280
rect 31352 30268 31358 30320
rect 33686 30308 33692 30320
rect 31404 30280 33692 30308
rect 30466 30240 30472 30252
rect 28776 30212 28948 30240
rect 29104 30212 30472 30240
rect 28776 30200 28782 30212
rect 28920 30181 28948 30212
rect 30466 30200 30472 30212
rect 30524 30200 30530 30252
rect 30837 30243 30895 30249
rect 30837 30209 30849 30243
rect 30883 30240 30895 30243
rect 31404 30240 31432 30280
rect 33686 30268 33692 30280
rect 33744 30268 33750 30320
rect 35802 30308 35808 30320
rect 34256 30280 35808 30308
rect 30883 30212 31432 30240
rect 30883 30209 30895 30212
rect 30837 30203 30895 30209
rect 28552 30144 28672 30172
rect 28813 30175 28871 30181
rect 18690 30064 18696 30116
rect 18748 30104 18754 30116
rect 25593 30107 25651 30113
rect 18748 30076 19334 30104
rect 18748 30064 18754 30076
rect 19306 30036 19334 30076
rect 25593 30073 25605 30107
rect 25639 30104 25651 30107
rect 26326 30104 26332 30116
rect 25639 30076 26332 30104
rect 25639 30073 25651 30076
rect 25593 30067 25651 30073
rect 26326 30064 26332 30076
rect 26384 30064 26390 30116
rect 27430 30064 27436 30116
rect 27488 30104 27494 30116
rect 28353 30107 28411 30113
rect 28353 30104 28365 30107
rect 27488 30076 28365 30104
rect 27488 30064 27494 30076
rect 28353 30073 28365 30076
rect 28399 30073 28411 30107
rect 28353 30067 28411 30073
rect 27801 30039 27859 30045
rect 27801 30036 27813 30039
rect 19306 30008 27813 30036
rect 27801 30005 27813 30008
rect 27847 30036 27859 30039
rect 28552 30036 28580 30144
rect 28813 30141 28825 30175
rect 28859 30141 28871 30175
rect 28813 30135 28871 30141
rect 28905 30175 28963 30181
rect 28905 30141 28917 30175
rect 28951 30141 28963 30175
rect 28905 30135 28963 30141
rect 28828 30104 28856 30135
rect 29454 30132 29460 30184
rect 29512 30172 29518 30184
rect 29917 30175 29975 30181
rect 29917 30172 29929 30175
rect 29512 30144 29929 30172
rect 29512 30132 29518 30144
rect 29917 30141 29929 30144
rect 29963 30172 29975 30175
rect 30852 30172 30880 30203
rect 32122 30200 32128 30252
rect 32180 30240 32186 30252
rect 34057 30243 34115 30249
rect 34057 30240 34069 30243
rect 32180 30212 34069 30240
rect 32180 30200 32186 30212
rect 34057 30209 34069 30212
rect 34103 30209 34115 30243
rect 34057 30203 34115 30209
rect 34146 30200 34152 30252
rect 34204 30200 34210 30252
rect 29963 30144 30880 30172
rect 30929 30175 30987 30181
rect 29963 30141 29975 30144
rect 29917 30135 29975 30141
rect 30929 30141 30941 30175
rect 30975 30141 30987 30175
rect 30929 30135 30987 30141
rect 31113 30175 31171 30181
rect 31113 30141 31125 30175
rect 31159 30172 31171 30175
rect 33962 30172 33968 30184
rect 31159 30144 33968 30172
rect 31159 30141 31171 30144
rect 31113 30135 31171 30141
rect 30944 30104 30972 30135
rect 33962 30132 33968 30144
rect 34020 30132 34026 30184
rect 34256 30181 34284 30280
rect 35802 30268 35808 30280
rect 35860 30268 35866 30320
rect 35897 30311 35955 30317
rect 35897 30277 35909 30311
rect 35943 30308 35955 30311
rect 36078 30308 36084 30320
rect 35943 30280 36084 30308
rect 35943 30277 35955 30280
rect 35897 30271 35955 30277
rect 36078 30268 36084 30280
rect 36136 30268 36142 30320
rect 37826 30268 37832 30320
rect 37884 30268 37890 30320
rect 37921 30311 37979 30317
rect 37921 30277 37933 30311
rect 37967 30308 37979 30311
rect 38286 30308 38292 30320
rect 37967 30280 38292 30308
rect 37967 30277 37979 30280
rect 37921 30271 37979 30277
rect 38286 30268 38292 30280
rect 38344 30268 38350 30320
rect 38470 30268 38476 30320
rect 38528 30308 38534 30320
rect 39025 30311 39083 30317
rect 39025 30308 39037 30311
rect 38528 30280 39037 30308
rect 38528 30268 38534 30280
rect 39025 30277 39037 30280
rect 39071 30277 39083 30311
rect 40250 30280 41414 30308
rect 39025 30271 39083 30277
rect 34422 30200 34428 30252
rect 34480 30240 34486 30252
rect 35989 30243 36047 30249
rect 34480 30212 35756 30240
rect 34480 30200 34486 30212
rect 34241 30175 34299 30181
rect 34241 30141 34253 30175
rect 34287 30141 34299 30175
rect 35728 30172 35756 30212
rect 35989 30209 36001 30243
rect 36035 30240 36047 30243
rect 37182 30240 37188 30252
rect 36035 30212 37188 30240
rect 36035 30209 36047 30212
rect 35989 30203 36047 30209
rect 37182 30200 37188 30212
rect 37240 30200 37246 30252
rect 41386 30240 41414 30280
rect 41690 30240 41696 30252
rect 41386 30212 41696 30240
rect 41690 30200 41696 30212
rect 41748 30240 41754 30252
rect 42610 30240 42616 30252
rect 41748 30212 42616 30240
rect 41748 30200 41754 30212
rect 42610 30200 42616 30212
rect 42668 30200 42674 30252
rect 49326 30200 49332 30252
rect 49384 30200 49390 30252
rect 36081 30175 36139 30181
rect 36081 30172 36093 30175
rect 34241 30135 34299 30141
rect 34348 30144 35664 30172
rect 35728 30144 36093 30172
rect 33870 30104 33876 30116
rect 28828 30076 30604 30104
rect 30944 30076 33876 30104
rect 27847 30008 28580 30036
rect 27847 30005 27859 30008
rect 27801 29999 27859 30005
rect 28626 29996 28632 30048
rect 28684 30036 28690 30048
rect 30469 30039 30527 30045
rect 30469 30036 30481 30039
rect 28684 30008 30481 30036
rect 28684 29996 28690 30008
rect 30469 30005 30481 30008
rect 30515 30005 30527 30039
rect 30576 30036 30604 30076
rect 33870 30064 33876 30076
rect 33928 30064 33934 30116
rect 34054 30064 34060 30116
rect 34112 30104 34118 30116
rect 34348 30104 34376 30144
rect 34112 30076 34376 30104
rect 34112 30064 34118 30076
rect 34606 30064 34612 30116
rect 34664 30104 34670 30116
rect 35529 30107 35587 30113
rect 35529 30104 35541 30107
rect 34664 30076 35541 30104
rect 34664 30064 34670 30076
rect 35529 30073 35541 30076
rect 35575 30073 35587 30107
rect 35636 30104 35664 30144
rect 36081 30141 36093 30144
rect 36127 30141 36139 30175
rect 38013 30175 38071 30181
rect 38013 30172 38025 30175
rect 36081 30135 36139 30141
rect 36188 30144 38025 30172
rect 36188 30104 36216 30144
rect 38013 30141 38025 30144
rect 38059 30141 38071 30175
rect 38013 30135 38071 30141
rect 38749 30175 38807 30181
rect 38749 30141 38761 30175
rect 38795 30172 38807 30175
rect 40678 30172 40684 30184
rect 38795 30144 40684 30172
rect 38795 30141 38807 30144
rect 38749 30135 38807 30141
rect 35636 30076 36216 30104
rect 35529 30067 35587 30073
rect 36262 30064 36268 30116
rect 36320 30104 36326 30116
rect 38764 30104 38792 30135
rect 40678 30132 40684 30144
rect 40736 30132 40742 30184
rect 40862 30132 40868 30184
rect 40920 30172 40926 30184
rect 41417 30175 41475 30181
rect 41417 30172 41429 30175
rect 40920 30144 41429 30172
rect 40920 30132 40926 30144
rect 41417 30141 41429 30144
rect 41463 30141 41475 30175
rect 41417 30135 41475 30141
rect 41509 30175 41567 30181
rect 41509 30141 41521 30175
rect 41555 30141 41567 30175
rect 41509 30135 41567 30141
rect 36320 30076 38792 30104
rect 36320 30064 36326 30076
rect 40126 30064 40132 30116
rect 40184 30104 40190 30116
rect 40957 30107 41015 30113
rect 40957 30104 40969 30107
rect 40184 30076 40969 30104
rect 40184 30064 40190 30076
rect 40957 30073 40969 30076
rect 41003 30073 41015 30107
rect 40957 30067 41015 30073
rect 41322 30064 41328 30116
rect 41380 30104 41386 30116
rect 41524 30104 41552 30135
rect 41380 30076 41552 30104
rect 41380 30064 41386 30076
rect 32766 30036 32772 30048
rect 30576 30008 32772 30036
rect 30469 29999 30527 30005
rect 32766 29996 32772 30008
rect 32824 29996 32830 30048
rect 33689 30039 33747 30045
rect 33689 30005 33701 30039
rect 33735 30036 33747 30039
rect 35158 30036 35164 30048
rect 33735 30008 35164 30036
rect 33735 30005 33747 30008
rect 33689 29999 33747 30005
rect 35158 29996 35164 30008
rect 35216 29996 35222 30048
rect 36170 29996 36176 30048
rect 36228 30036 36234 30048
rect 37461 30039 37519 30045
rect 37461 30036 37473 30039
rect 36228 30008 37473 30036
rect 36228 29996 36234 30008
rect 37461 30005 37473 30008
rect 37507 30005 37519 30039
rect 37461 29999 37519 30005
rect 40494 29996 40500 30048
rect 40552 29996 40558 30048
rect 45738 29996 45744 30048
rect 45796 30036 45802 30048
rect 49145 30039 49203 30045
rect 49145 30036 49157 30039
rect 45796 30008 49157 30036
rect 45796 29996 45802 30008
rect 49145 30005 49157 30008
rect 49191 30005 49203 30039
rect 49145 29999 49203 30005
rect 1104 29946 49864 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 32950 29946
rect 33002 29894 33014 29946
rect 33066 29894 33078 29946
rect 33130 29894 33142 29946
rect 33194 29894 33206 29946
rect 33258 29894 42950 29946
rect 43002 29894 43014 29946
rect 43066 29894 43078 29946
rect 43130 29894 43142 29946
rect 43194 29894 43206 29946
rect 43258 29894 49864 29946
rect 1104 29872 49864 29894
rect 10686 29792 10692 29844
rect 10744 29832 10750 29844
rect 25590 29832 25596 29844
rect 10744 29804 25596 29832
rect 10744 29792 10750 29804
rect 25590 29792 25596 29804
rect 25648 29792 25654 29844
rect 28810 29792 28816 29844
rect 28868 29832 28874 29844
rect 28868 29804 30236 29832
rect 28868 29792 28874 29804
rect 25317 29767 25375 29773
rect 25317 29733 25329 29767
rect 25363 29764 25375 29767
rect 25363 29736 30052 29764
rect 25363 29733 25375 29736
rect 25317 29727 25375 29733
rect 1302 29656 1308 29708
rect 1360 29696 1366 29708
rect 2041 29699 2099 29705
rect 2041 29696 2053 29699
rect 1360 29668 2053 29696
rect 1360 29656 1366 29668
rect 2041 29665 2053 29668
rect 2087 29665 2099 29699
rect 2041 29659 2099 29665
rect 21082 29656 21088 29708
rect 21140 29696 21146 29708
rect 21913 29699 21971 29705
rect 21913 29696 21925 29699
rect 21140 29668 21925 29696
rect 21140 29656 21146 29668
rect 21913 29665 21925 29668
rect 21959 29665 21971 29699
rect 21913 29659 21971 29665
rect 25961 29699 26019 29705
rect 25961 29665 25973 29699
rect 26007 29696 26019 29699
rect 27338 29696 27344 29708
rect 26007 29668 27344 29696
rect 26007 29665 26019 29668
rect 25961 29659 26019 29665
rect 27338 29656 27344 29668
rect 27396 29656 27402 29708
rect 27522 29656 27528 29708
rect 27580 29696 27586 29708
rect 29362 29696 29368 29708
rect 27580 29668 29368 29696
rect 27580 29656 27586 29668
rect 29362 29656 29368 29668
rect 29420 29656 29426 29708
rect 30024 29696 30052 29736
rect 30208 29696 30236 29804
rect 30466 29792 30472 29844
rect 30524 29832 30530 29844
rect 30524 29804 31754 29832
rect 30524 29792 30530 29804
rect 31726 29764 31754 29804
rect 32214 29792 32220 29844
rect 32272 29832 32278 29844
rect 34422 29832 34428 29844
rect 32272 29804 34428 29832
rect 32272 29792 32278 29804
rect 34422 29792 34428 29804
rect 34480 29792 34486 29844
rect 34698 29792 34704 29844
rect 34756 29832 34762 29844
rect 34756 29804 36400 29832
rect 34756 29792 34762 29804
rect 35250 29764 35256 29776
rect 31726 29736 35256 29764
rect 35250 29724 35256 29736
rect 35308 29724 35314 29776
rect 36372 29764 36400 29804
rect 36446 29792 36452 29844
rect 36504 29832 36510 29844
rect 38749 29835 38807 29841
rect 38749 29832 38761 29835
rect 36504 29804 38761 29832
rect 36504 29792 36510 29804
rect 38749 29801 38761 29804
rect 38795 29801 38807 29835
rect 38749 29795 38807 29801
rect 42702 29792 42708 29844
rect 42760 29792 42766 29844
rect 36372 29736 36584 29764
rect 30285 29699 30343 29705
rect 30285 29696 30297 29699
rect 30024 29668 30144 29696
rect 30208 29668 30297 29696
rect 1765 29631 1823 29637
rect 1765 29597 1777 29631
rect 1811 29628 1823 29631
rect 4798 29628 4804 29640
rect 1811 29600 4804 29628
rect 1811 29597 1823 29600
rect 1765 29591 1823 29597
rect 4798 29588 4804 29600
rect 4856 29588 4862 29640
rect 25685 29631 25743 29637
rect 25685 29597 25697 29631
rect 25731 29628 25743 29631
rect 26697 29631 26755 29637
rect 26697 29628 26709 29631
rect 25731 29600 26709 29628
rect 25731 29597 25743 29600
rect 25685 29591 25743 29597
rect 26697 29597 26709 29600
rect 26743 29597 26755 29631
rect 26697 29591 26755 29597
rect 27062 29588 27068 29640
rect 27120 29628 27126 29640
rect 30006 29628 30012 29640
rect 27120 29600 30012 29628
rect 27120 29588 27126 29600
rect 30006 29588 30012 29600
rect 30064 29588 30070 29640
rect 30116 29637 30144 29668
rect 30285 29665 30297 29668
rect 30331 29665 30343 29699
rect 30285 29659 30343 29665
rect 30466 29656 30472 29708
rect 30524 29696 30530 29708
rect 32493 29699 32551 29705
rect 32493 29696 32505 29699
rect 30524 29668 32505 29696
rect 30524 29656 30530 29668
rect 32493 29665 32505 29668
rect 32539 29665 32551 29699
rect 32493 29659 32551 29665
rect 33870 29656 33876 29708
rect 33928 29696 33934 29708
rect 34698 29696 34704 29708
rect 33928 29668 34704 29696
rect 33928 29656 33934 29668
rect 34698 29656 34704 29668
rect 34756 29656 34762 29708
rect 36262 29656 36268 29708
rect 36320 29696 36326 29708
rect 36449 29699 36507 29705
rect 36449 29696 36461 29699
rect 36320 29668 36461 29696
rect 36320 29656 36326 29668
rect 36449 29665 36461 29668
rect 36495 29665 36507 29699
rect 36556 29696 36584 29736
rect 38562 29724 38568 29776
rect 38620 29764 38626 29776
rect 38620 29736 41092 29764
rect 38620 29724 38626 29736
rect 36725 29699 36783 29705
rect 36725 29696 36737 29699
rect 36556 29668 36737 29696
rect 36449 29659 36507 29665
rect 36725 29665 36737 29668
rect 36771 29696 36783 29699
rect 37458 29696 37464 29708
rect 36771 29668 37464 29696
rect 36771 29665 36783 29668
rect 36725 29659 36783 29665
rect 37458 29656 37464 29668
rect 37516 29656 37522 29708
rect 39393 29699 39451 29705
rect 39393 29665 39405 29699
rect 39439 29696 39451 29699
rect 39758 29696 39764 29708
rect 39439 29668 39764 29696
rect 39439 29665 39451 29668
rect 39393 29659 39451 29665
rect 39758 29656 39764 29668
rect 39816 29656 39822 29708
rect 40310 29656 40316 29708
rect 40368 29696 40374 29708
rect 40678 29696 40684 29708
rect 40368 29668 40684 29696
rect 40368 29656 40374 29668
rect 40678 29656 40684 29668
rect 40736 29696 40742 29708
rect 40957 29699 41015 29705
rect 40957 29696 40969 29699
rect 40736 29668 40969 29696
rect 40736 29656 40742 29668
rect 40957 29665 40969 29668
rect 41003 29665 41015 29699
rect 41064 29696 41092 29736
rect 48777 29699 48835 29705
rect 48777 29696 48789 29699
rect 41064 29668 48789 29696
rect 40957 29659 41015 29665
rect 48777 29665 48789 29668
rect 48823 29665 48835 29699
rect 48777 29659 48835 29665
rect 30101 29631 30159 29637
rect 30101 29597 30113 29631
rect 30147 29597 30159 29631
rect 30101 29591 30159 29597
rect 32309 29631 32367 29637
rect 32309 29597 32321 29631
rect 32355 29628 32367 29631
rect 34238 29628 34244 29640
rect 32355 29600 34244 29628
rect 32355 29597 32367 29600
rect 32309 29591 32367 29597
rect 34238 29588 34244 29600
rect 34296 29588 34302 29640
rect 39117 29631 39175 29637
rect 39117 29597 39129 29631
rect 39163 29628 39175 29631
rect 40770 29628 40776 29640
rect 39163 29600 40776 29628
rect 39163 29597 39175 29600
rect 39117 29591 39175 29597
rect 40770 29588 40776 29600
rect 40828 29588 40834 29640
rect 48498 29588 48504 29640
rect 48556 29588 48562 29640
rect 21174 29520 21180 29572
rect 21232 29520 21238 29572
rect 28534 29520 28540 29572
rect 28592 29560 28598 29572
rect 28718 29560 28724 29572
rect 28592 29532 28724 29560
rect 28592 29520 28598 29532
rect 28718 29520 28724 29532
rect 28776 29560 28782 29572
rect 29454 29560 29460 29572
rect 28776 29532 29460 29560
rect 28776 29520 28782 29532
rect 29454 29520 29460 29532
rect 29512 29520 29518 29572
rect 36630 29560 36636 29572
rect 29748 29532 36636 29560
rect 22738 29452 22744 29504
rect 22796 29492 22802 29504
rect 23658 29492 23664 29504
rect 22796 29464 23664 29492
rect 22796 29452 22802 29464
rect 23658 29452 23664 29464
rect 23716 29492 23722 29504
rect 29748 29501 29776 29532
rect 36630 29520 36636 29532
rect 36688 29520 36694 29572
rect 37274 29520 37280 29572
rect 37332 29520 37338 29572
rect 40494 29520 40500 29572
rect 40552 29560 40558 29572
rect 41233 29563 41291 29569
rect 41233 29560 41245 29563
rect 40552 29532 41245 29560
rect 40552 29520 40558 29532
rect 41233 29529 41245 29532
rect 41279 29529 41291 29563
rect 41233 29523 41291 29529
rect 41690 29520 41696 29572
rect 41748 29520 41754 29572
rect 25777 29495 25835 29501
rect 25777 29492 25789 29495
rect 23716 29464 25789 29492
rect 23716 29452 23722 29464
rect 25777 29461 25789 29464
rect 25823 29461 25835 29495
rect 25777 29455 25835 29461
rect 29733 29495 29791 29501
rect 29733 29461 29745 29495
rect 29779 29461 29791 29495
rect 29733 29455 29791 29461
rect 29914 29452 29920 29504
rect 29972 29492 29978 29504
rect 30193 29495 30251 29501
rect 30193 29492 30205 29495
rect 29972 29464 30205 29492
rect 29972 29452 29978 29464
rect 30193 29461 30205 29464
rect 30239 29461 30251 29495
rect 30193 29455 30251 29461
rect 31938 29452 31944 29504
rect 31996 29452 32002 29504
rect 32398 29452 32404 29504
rect 32456 29492 32462 29504
rect 35894 29492 35900 29504
rect 32456 29464 35900 29492
rect 32456 29452 32462 29464
rect 35894 29452 35900 29464
rect 35952 29452 35958 29504
rect 36262 29452 36268 29504
rect 36320 29492 36326 29504
rect 38197 29495 38255 29501
rect 38197 29492 38209 29495
rect 36320 29464 38209 29492
rect 36320 29452 36326 29464
rect 38197 29461 38209 29464
rect 38243 29461 38255 29495
rect 38197 29455 38255 29461
rect 39209 29495 39267 29501
rect 39209 29461 39221 29495
rect 39255 29492 39267 29495
rect 41414 29492 41420 29504
rect 39255 29464 41420 29492
rect 39255 29461 39267 29464
rect 39209 29455 39267 29461
rect 41414 29452 41420 29464
rect 41472 29452 41478 29504
rect 1104 29402 49864 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 27950 29402
rect 28002 29350 28014 29402
rect 28066 29350 28078 29402
rect 28130 29350 28142 29402
rect 28194 29350 28206 29402
rect 28258 29350 37950 29402
rect 38002 29350 38014 29402
rect 38066 29350 38078 29402
rect 38130 29350 38142 29402
rect 38194 29350 38206 29402
rect 38258 29350 47950 29402
rect 48002 29350 48014 29402
rect 48066 29350 48078 29402
rect 48130 29350 48142 29402
rect 48194 29350 48206 29402
rect 48258 29350 49864 29402
rect 1104 29328 49864 29350
rect 22005 29291 22063 29297
rect 22005 29257 22017 29291
rect 22051 29288 22063 29291
rect 23290 29288 23296 29300
rect 22051 29260 23296 29288
rect 22051 29257 22063 29260
rect 22005 29251 22063 29257
rect 23290 29248 23296 29260
rect 23348 29248 23354 29300
rect 28810 29288 28816 29300
rect 28000 29260 28816 29288
rect 17218 29180 17224 29232
rect 17276 29220 17282 29232
rect 28000 29229 28028 29260
rect 28810 29248 28816 29260
rect 28868 29248 28874 29300
rect 30098 29248 30104 29300
rect 30156 29288 30162 29300
rect 30466 29288 30472 29300
rect 30156 29260 30472 29288
rect 30156 29248 30162 29260
rect 30466 29248 30472 29260
rect 30524 29248 30530 29300
rect 34146 29248 34152 29300
rect 34204 29288 34210 29300
rect 34422 29288 34428 29300
rect 34204 29260 34428 29288
rect 34204 29248 34210 29260
rect 34422 29248 34428 29260
rect 34480 29248 34486 29300
rect 35526 29248 35532 29300
rect 35584 29288 35590 29300
rect 35713 29291 35771 29297
rect 35713 29288 35725 29291
rect 35584 29260 35725 29288
rect 35584 29248 35590 29260
rect 35713 29257 35725 29260
rect 35759 29257 35771 29291
rect 35713 29251 35771 29257
rect 40034 29248 40040 29300
rect 40092 29288 40098 29300
rect 41233 29291 41291 29297
rect 41233 29288 41245 29291
rect 40092 29260 41245 29288
rect 40092 29248 40098 29260
rect 41233 29257 41245 29260
rect 41279 29257 41291 29291
rect 41233 29251 41291 29257
rect 27985 29223 28043 29229
rect 17276 29192 22508 29220
rect 17276 29180 17282 29192
rect 22370 29112 22376 29164
rect 22428 29112 22434 29164
rect 22480 29161 22508 29192
rect 27985 29189 27997 29223
rect 28031 29189 28043 29223
rect 29730 29220 29736 29232
rect 29210 29192 29736 29220
rect 27985 29183 28043 29189
rect 29730 29180 29736 29192
rect 29788 29180 29794 29232
rect 30285 29223 30343 29229
rect 30285 29189 30297 29223
rect 30331 29220 30343 29223
rect 33502 29220 33508 29232
rect 30331 29192 33508 29220
rect 30331 29189 30343 29192
rect 30285 29183 30343 29189
rect 33502 29180 33508 29192
rect 33560 29220 33566 29232
rect 33778 29220 33784 29232
rect 33560 29192 33784 29220
rect 33560 29180 33566 29192
rect 33778 29180 33784 29192
rect 33836 29180 33842 29232
rect 34790 29180 34796 29232
rect 34848 29180 34854 29232
rect 37642 29180 37648 29232
rect 37700 29220 37706 29232
rect 41322 29220 41328 29232
rect 37700 29192 41328 29220
rect 37700 29180 37706 29192
rect 41322 29180 41328 29192
rect 41380 29180 41386 29232
rect 22465 29155 22523 29161
rect 22465 29121 22477 29155
rect 22511 29152 22523 29155
rect 23290 29152 23296 29164
rect 22511 29124 23296 29152
rect 22511 29121 22523 29124
rect 22465 29115 22523 29121
rect 23290 29112 23296 29124
rect 23348 29112 23354 29164
rect 27062 29112 27068 29164
rect 27120 29152 27126 29164
rect 27709 29155 27767 29161
rect 27709 29152 27721 29155
rect 27120 29124 27721 29152
rect 27120 29112 27126 29124
rect 27709 29121 27721 29124
rect 27755 29121 27767 29155
rect 27709 29115 27767 29121
rect 29270 29112 29276 29164
rect 29328 29152 29334 29164
rect 29546 29152 29552 29164
rect 29328 29124 29552 29152
rect 29328 29112 29334 29124
rect 29546 29112 29552 29124
rect 29604 29152 29610 29164
rect 32398 29152 32404 29164
rect 29604 29124 32404 29152
rect 29604 29112 29610 29124
rect 32398 29112 32404 29124
rect 32456 29112 32462 29164
rect 41138 29112 41144 29164
rect 41196 29112 41202 29164
rect 41248 29124 45554 29152
rect 22649 29087 22707 29093
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 25130 29084 25136 29096
rect 22695 29056 25136 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 25130 29044 25136 29056
rect 25188 29044 25194 29096
rect 30377 29087 30435 29093
rect 30377 29084 30389 29087
rect 26160 29056 30389 29084
rect 26160 29028 26188 29056
rect 7742 28976 7748 29028
rect 7800 29016 7806 29028
rect 21177 29019 21235 29025
rect 21177 29016 21189 29019
rect 7800 28988 21189 29016
rect 7800 28976 7806 28988
rect 21177 28985 21189 28988
rect 21223 29016 21235 29019
rect 22370 29016 22376 29028
rect 21223 28988 22376 29016
rect 21223 28985 21235 28988
rect 21177 28979 21235 28985
rect 22370 28976 22376 28988
rect 22428 28976 22434 29028
rect 25682 28976 25688 29028
rect 25740 29016 25746 29028
rect 26142 29016 26148 29028
rect 25740 28988 26148 29016
rect 25740 28976 25746 28988
rect 26142 28976 26148 28988
rect 26200 28976 26206 29028
rect 28994 28976 29000 29028
rect 29052 29016 29058 29028
rect 29917 29019 29975 29025
rect 29917 29016 29929 29019
rect 29052 28988 29929 29016
rect 29052 28976 29058 28988
rect 29917 28985 29929 28988
rect 29963 28985 29975 29019
rect 29917 28979 29975 28985
rect 30208 28994 30236 29056
rect 30377 29053 30389 29056
rect 30423 29053 30435 29087
rect 30377 29047 30435 29053
rect 30466 29044 30472 29096
rect 30524 29044 30530 29096
rect 33962 29044 33968 29096
rect 34020 29044 34026 29096
rect 37274 29044 37280 29096
rect 37332 29084 37338 29096
rect 37826 29084 37832 29096
rect 37332 29056 37832 29084
rect 37332 29044 37338 29056
rect 37826 29044 37832 29056
rect 37884 29044 37890 29096
rect 38654 29044 38660 29096
rect 38712 29084 38718 29096
rect 39022 29084 39028 29096
rect 38712 29056 39028 29084
rect 38712 29044 38718 29056
rect 39022 29044 39028 29056
rect 39080 29084 39086 29096
rect 41248 29084 41276 29124
rect 39080 29056 41276 29084
rect 41417 29087 41475 29093
rect 39080 29044 39086 29056
rect 41417 29053 41429 29087
rect 41463 29084 41475 29087
rect 42702 29084 42708 29096
rect 41463 29056 42708 29084
rect 41463 29053 41475 29056
rect 41417 29047 41475 29053
rect 42702 29044 42708 29056
rect 42760 29044 42766 29096
rect 32122 29016 32128 29028
rect 30208 28966 30328 28994
rect 28534 28908 28540 28960
rect 28592 28948 28598 28960
rect 29454 28948 29460 28960
rect 28592 28920 29460 28948
rect 28592 28908 28598 28920
rect 29454 28908 29460 28920
rect 29512 28908 29518 28960
rect 30300 28948 30328 28966
rect 30576 28988 32128 29016
rect 30576 28948 30604 28988
rect 32122 28976 32128 28988
rect 32180 28976 32186 29028
rect 35802 28976 35808 29028
rect 35860 29016 35866 29028
rect 39390 29016 39396 29028
rect 35860 28988 39396 29016
rect 35860 28976 35866 28988
rect 39390 28976 39396 28988
rect 39448 28976 39454 29028
rect 40773 29019 40831 29025
rect 40773 28985 40785 29019
rect 40819 29016 40831 29019
rect 44174 29016 44180 29028
rect 40819 28988 44180 29016
rect 40819 28985 40831 28988
rect 40773 28979 40831 28985
rect 44174 28976 44180 28988
rect 44232 28976 44238 29028
rect 45526 29016 45554 29124
rect 49326 29112 49332 29164
rect 49384 29112 49390 29164
rect 49145 29019 49203 29025
rect 49145 29016 49157 29019
rect 45526 28988 49157 29016
rect 49145 28985 49157 28988
rect 49191 28985 49203 29019
rect 49145 28979 49203 28985
rect 30300 28920 30604 28948
rect 32030 28908 32036 28960
rect 32088 28948 32094 28960
rect 32582 28948 32588 28960
rect 32088 28920 32588 28948
rect 32088 28908 32094 28920
rect 32582 28908 32588 28920
rect 32640 28908 32646 28960
rect 34228 28951 34286 28957
rect 34228 28917 34240 28951
rect 34274 28948 34286 28951
rect 36262 28948 36268 28960
rect 34274 28920 36268 28948
rect 34274 28917 34286 28920
rect 34228 28911 34286 28917
rect 36262 28908 36268 28920
rect 36320 28908 36326 28960
rect 36354 28908 36360 28960
rect 36412 28908 36418 28960
rect 1104 28858 49864 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 32950 28858
rect 33002 28806 33014 28858
rect 33066 28806 33078 28858
rect 33130 28806 33142 28858
rect 33194 28806 33206 28858
rect 33258 28806 42950 28858
rect 43002 28806 43014 28858
rect 43066 28806 43078 28858
rect 43130 28806 43142 28858
rect 43194 28806 43206 28858
rect 43258 28806 49864 28858
rect 1104 28784 49864 28806
rect 22186 28704 22192 28756
rect 22244 28704 22250 28756
rect 35434 28704 35440 28756
rect 35492 28744 35498 28756
rect 39114 28744 39120 28756
rect 35492 28716 39120 28744
rect 35492 28704 35498 28716
rect 39114 28704 39120 28716
rect 39172 28704 39178 28756
rect 27614 28636 27620 28688
rect 27672 28676 27678 28688
rect 28810 28676 28816 28688
rect 27672 28648 28816 28676
rect 27672 28636 27678 28648
rect 28810 28636 28816 28648
rect 28868 28636 28874 28688
rect 36814 28676 36820 28688
rect 35360 28648 36820 28676
rect 22554 28568 22560 28620
rect 22612 28608 22618 28620
rect 22649 28611 22707 28617
rect 22649 28608 22661 28611
rect 22612 28580 22661 28608
rect 22612 28568 22618 28580
rect 22649 28577 22661 28580
rect 22695 28577 22707 28611
rect 22649 28571 22707 28577
rect 22833 28611 22891 28617
rect 22833 28577 22845 28611
rect 22879 28608 22891 28611
rect 23382 28608 23388 28620
rect 22879 28580 23388 28608
rect 22879 28577 22891 28580
rect 22833 28571 22891 28577
rect 23382 28568 23388 28580
rect 23440 28568 23446 28620
rect 29454 28568 29460 28620
rect 29512 28608 29518 28620
rect 31297 28611 31355 28617
rect 31297 28608 31309 28611
rect 29512 28580 31309 28608
rect 29512 28568 29518 28580
rect 31297 28577 31309 28580
rect 31343 28577 31355 28611
rect 31297 28571 31355 28577
rect 32858 28568 32864 28620
rect 32916 28608 32922 28620
rect 34057 28611 34115 28617
rect 34057 28608 34069 28611
rect 32916 28580 34069 28608
rect 32916 28568 32922 28580
rect 34057 28577 34069 28580
rect 34103 28577 34115 28611
rect 34057 28571 34115 28577
rect 34146 28568 34152 28620
rect 34204 28568 34210 28620
rect 24946 28500 24952 28552
rect 25004 28540 25010 28552
rect 26329 28543 26387 28549
rect 26329 28540 26341 28543
rect 25004 28512 26341 28540
rect 25004 28500 25010 28512
rect 26329 28509 26341 28512
rect 26375 28540 26387 28543
rect 27614 28540 27620 28552
rect 26375 28512 27620 28540
rect 26375 28509 26387 28512
rect 26329 28503 26387 28509
rect 27614 28500 27620 28512
rect 27672 28500 27678 28552
rect 29914 28500 29920 28552
rect 29972 28500 29978 28552
rect 31113 28543 31171 28549
rect 31113 28509 31125 28543
rect 31159 28540 31171 28543
rect 33318 28540 33324 28552
rect 31159 28512 33324 28540
rect 31159 28509 31171 28512
rect 31113 28503 31171 28509
rect 33318 28500 33324 28512
rect 33376 28540 33382 28552
rect 33778 28540 33784 28552
rect 33376 28512 33784 28540
rect 33376 28500 33382 28512
rect 33778 28500 33784 28512
rect 33836 28500 33842 28552
rect 33965 28543 34023 28549
rect 33965 28509 33977 28543
rect 34011 28540 34023 28543
rect 35360 28540 35388 28648
rect 36814 28636 36820 28648
rect 36872 28636 36878 28688
rect 39206 28636 39212 28688
rect 39264 28676 39270 28688
rect 39482 28676 39488 28688
rect 39264 28648 39488 28676
rect 39264 28636 39270 28648
rect 39482 28636 39488 28648
rect 39540 28676 39546 28688
rect 49145 28679 49203 28685
rect 49145 28676 49157 28679
rect 39540 28648 49157 28676
rect 39540 28636 39546 28648
rect 49145 28645 49157 28648
rect 49191 28645 49203 28679
rect 49145 28639 49203 28645
rect 35529 28611 35587 28617
rect 35529 28577 35541 28611
rect 35575 28608 35587 28611
rect 35802 28608 35808 28620
rect 35575 28580 35808 28608
rect 35575 28577 35587 28580
rect 35529 28571 35587 28577
rect 35802 28568 35808 28580
rect 35860 28568 35866 28620
rect 36262 28568 36268 28620
rect 36320 28608 36326 28620
rect 36633 28611 36691 28617
rect 36633 28608 36645 28611
rect 36320 28580 36645 28608
rect 36320 28568 36326 28580
rect 36633 28577 36645 28580
rect 36679 28577 36691 28611
rect 36633 28571 36691 28577
rect 37921 28611 37979 28617
rect 37921 28577 37933 28611
rect 37967 28608 37979 28611
rect 38286 28608 38292 28620
rect 37967 28580 38292 28608
rect 37967 28577 37979 28580
rect 37921 28571 37979 28577
rect 38286 28568 38292 28580
rect 38344 28568 38350 28620
rect 40218 28608 40224 28620
rect 38580 28580 40224 28608
rect 34011 28512 35388 28540
rect 34011 28509 34023 28512
rect 33965 28503 34023 28509
rect 36354 28500 36360 28552
rect 36412 28540 36418 28552
rect 36449 28543 36507 28549
rect 36449 28540 36461 28543
rect 36412 28512 36461 28540
rect 36412 28500 36418 28512
rect 36449 28509 36461 28512
rect 36495 28509 36507 28543
rect 36449 28503 36507 28509
rect 37645 28543 37703 28549
rect 37645 28509 37657 28543
rect 37691 28540 37703 28543
rect 38580 28540 38608 28580
rect 40218 28568 40224 28580
rect 40276 28568 40282 28620
rect 40678 28568 40684 28620
rect 40736 28568 40742 28620
rect 37691 28512 38608 28540
rect 38657 28543 38715 28549
rect 37691 28509 37703 28512
rect 37645 28503 37703 28509
rect 38657 28509 38669 28543
rect 38703 28540 38715 28543
rect 39022 28540 39028 28552
rect 38703 28512 39028 28540
rect 38703 28509 38715 28512
rect 38657 28503 38715 28509
rect 39022 28500 39028 28512
rect 39080 28500 39086 28552
rect 40405 28543 40463 28549
rect 40405 28509 40417 28543
rect 40451 28540 40463 28543
rect 41046 28540 41052 28552
rect 40451 28512 41052 28540
rect 40451 28509 40463 28512
rect 40405 28503 40463 28509
rect 41046 28500 41052 28512
rect 41104 28500 41110 28552
rect 49326 28500 49332 28552
rect 49384 28500 49390 28552
rect 22066 28444 22600 28472
rect 7098 28364 7104 28416
rect 7156 28404 7162 28416
rect 19334 28404 19340 28416
rect 7156 28376 19340 28404
rect 7156 28364 7162 28376
rect 19334 28364 19340 28376
rect 19392 28404 19398 28416
rect 21637 28407 21695 28413
rect 21637 28404 21649 28407
rect 19392 28376 21649 28404
rect 19392 28364 19398 28376
rect 21637 28373 21649 28376
rect 21683 28404 21695 28407
rect 22066 28404 22094 28444
rect 22572 28416 22600 28444
rect 25498 28432 25504 28484
rect 25556 28432 25562 28484
rect 27062 28432 27068 28484
rect 27120 28432 27126 28484
rect 30190 28432 30196 28484
rect 30248 28472 30254 28484
rect 30248 28444 31248 28472
rect 30248 28432 30254 28444
rect 21683 28376 22094 28404
rect 21683 28373 21695 28376
rect 21637 28367 21695 28373
rect 22554 28364 22560 28416
rect 22612 28364 22618 28416
rect 25516 28404 25544 28432
rect 28350 28404 28356 28416
rect 25516 28376 28356 28404
rect 28350 28364 28356 28376
rect 28408 28364 28414 28416
rect 30745 28407 30803 28413
rect 30745 28373 30757 28407
rect 30791 28404 30803 28407
rect 31110 28404 31116 28416
rect 30791 28376 31116 28404
rect 30791 28373 30803 28376
rect 30745 28367 30803 28373
rect 31110 28364 31116 28376
rect 31168 28364 31174 28416
rect 31220 28413 31248 28444
rect 35158 28432 35164 28484
rect 35216 28472 35222 28484
rect 37737 28475 37795 28481
rect 37737 28472 37749 28475
rect 35216 28444 37749 28472
rect 35216 28432 35222 28444
rect 37737 28441 37749 28444
rect 37783 28441 37795 28475
rect 37737 28435 37795 28441
rect 38930 28432 38936 28484
rect 38988 28472 38994 28484
rect 40497 28475 40555 28481
rect 40497 28472 40509 28475
rect 38988 28444 40509 28472
rect 38988 28432 38994 28444
rect 40497 28441 40509 28444
rect 40543 28441 40555 28475
rect 40497 28435 40555 28441
rect 31205 28407 31263 28413
rect 31205 28373 31217 28407
rect 31251 28404 31263 28407
rect 31294 28404 31300 28416
rect 31251 28376 31300 28404
rect 31251 28373 31263 28376
rect 31205 28367 31263 28373
rect 31294 28364 31300 28376
rect 31352 28364 31358 28416
rect 32858 28364 32864 28416
rect 32916 28404 32922 28416
rect 33597 28407 33655 28413
rect 33597 28404 33609 28407
rect 32916 28376 33609 28404
rect 32916 28364 32922 28376
rect 33597 28373 33609 28376
rect 33643 28373 33655 28407
rect 33597 28367 33655 28373
rect 34885 28407 34943 28413
rect 34885 28373 34897 28407
rect 34931 28404 34943 28407
rect 35066 28404 35072 28416
rect 34931 28376 35072 28404
rect 34931 28373 34943 28376
rect 34885 28367 34943 28373
rect 35066 28364 35072 28376
rect 35124 28364 35130 28416
rect 35250 28364 35256 28416
rect 35308 28364 35314 28416
rect 35345 28407 35403 28413
rect 35345 28373 35357 28407
rect 35391 28404 35403 28407
rect 35434 28404 35440 28416
rect 35391 28376 35440 28404
rect 35391 28373 35403 28376
rect 35345 28367 35403 28373
rect 35434 28364 35440 28376
rect 35492 28364 35498 28416
rect 36078 28364 36084 28416
rect 36136 28364 36142 28416
rect 36538 28364 36544 28416
rect 36596 28364 36602 28416
rect 37274 28364 37280 28416
rect 37332 28364 37338 28416
rect 40037 28407 40095 28413
rect 40037 28373 40049 28407
rect 40083 28404 40095 28407
rect 40218 28404 40224 28416
rect 40083 28376 40224 28404
rect 40083 28373 40095 28376
rect 40037 28367 40095 28373
rect 40218 28364 40224 28376
rect 40276 28364 40282 28416
rect 1104 28314 49864 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 27950 28314
rect 28002 28262 28014 28314
rect 28066 28262 28078 28314
rect 28130 28262 28142 28314
rect 28194 28262 28206 28314
rect 28258 28262 37950 28314
rect 38002 28262 38014 28314
rect 38066 28262 38078 28314
rect 38130 28262 38142 28314
rect 38194 28262 38206 28314
rect 38258 28262 47950 28314
rect 48002 28262 48014 28314
rect 48066 28262 48078 28314
rect 48130 28262 48142 28314
rect 48194 28262 48206 28314
rect 48258 28262 49864 28314
rect 1104 28240 49864 28262
rect 4798 28160 4804 28212
rect 4856 28160 4862 28212
rect 26421 28203 26479 28209
rect 22480 28172 24716 28200
rect 20533 28135 20591 28141
rect 20533 28101 20545 28135
rect 20579 28132 20591 28135
rect 21174 28132 21180 28144
rect 20579 28104 21180 28132
rect 20579 28101 20591 28104
rect 20533 28095 20591 28101
rect 21174 28092 21180 28104
rect 21232 28092 21238 28144
rect 4985 28067 5043 28073
rect 4985 28033 4997 28067
rect 5031 28064 5043 28067
rect 5031 28036 6914 28064
rect 5031 28033 5043 28036
rect 4985 28027 5043 28033
rect 6886 27928 6914 28036
rect 7558 28024 7564 28076
rect 7616 28024 7622 28076
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22480 28073 22508 28172
rect 24688 28132 24716 28172
rect 26421 28169 26433 28203
rect 26467 28200 26479 28203
rect 30282 28200 30288 28212
rect 26467 28172 30288 28200
rect 26467 28169 26479 28172
rect 26421 28163 26479 28169
rect 24946 28132 24952 28144
rect 24688 28104 24952 28132
rect 22465 28067 22523 28073
rect 22465 28064 22477 28067
rect 22152 28036 22477 28064
rect 22152 28024 22158 28036
rect 22465 28033 22477 28036
rect 22511 28033 22523 28067
rect 22465 28027 22523 28033
rect 23842 28024 23848 28076
rect 23900 28024 23906 28076
rect 24688 28073 24716 28104
rect 24946 28092 24952 28104
rect 25004 28092 25010 28144
rect 26234 28132 26240 28144
rect 26174 28104 26240 28132
rect 26234 28092 26240 28104
rect 26292 28092 26298 28144
rect 24673 28067 24731 28073
rect 24673 28033 24685 28067
rect 24719 28033 24731 28067
rect 24673 28027 24731 28033
rect 7742 27956 7748 28008
rect 7800 27956 7806 28008
rect 9401 27999 9459 28005
rect 9401 27965 9413 27999
rect 9447 27996 9459 27999
rect 9490 27996 9496 28008
rect 9447 27968 9496 27996
rect 9447 27965 9459 27968
rect 9401 27959 9459 27965
rect 9490 27956 9496 27968
rect 9548 27956 9554 28008
rect 21361 27999 21419 28005
rect 21361 27965 21373 27999
rect 21407 27996 21419 27999
rect 21450 27996 21456 28008
rect 21407 27968 21456 27996
rect 21407 27965 21419 27968
rect 21361 27959 21419 27965
rect 21450 27956 21456 27968
rect 21508 27956 21514 28008
rect 22741 27999 22799 28005
rect 22741 27965 22753 27999
rect 22787 27996 22799 27999
rect 23382 27996 23388 28008
rect 22787 27968 23388 27996
rect 22787 27965 22799 27968
rect 22741 27959 22799 27965
rect 23382 27956 23388 27968
rect 23440 27996 23446 28008
rect 24949 27999 25007 28005
rect 23440 27968 24808 27996
rect 23440 27956 23446 27968
rect 9674 27928 9680 27940
rect 6886 27900 9680 27928
rect 9674 27888 9680 27900
rect 9732 27888 9738 27940
rect 24210 27820 24216 27872
rect 24268 27820 24274 27872
rect 24780 27860 24808 27968
rect 24949 27965 24961 27999
rect 24995 27996 25007 27999
rect 26694 27996 26700 28008
rect 24995 27968 26700 27996
rect 24995 27965 25007 27968
rect 24949 27959 25007 27965
rect 26694 27956 26700 27968
rect 26752 27956 26758 28008
rect 26804 27860 26832 28172
rect 30282 28160 30288 28172
rect 30340 28160 30346 28212
rect 32122 28160 32128 28212
rect 32180 28200 32186 28212
rect 33410 28200 33416 28212
rect 32180 28172 33416 28200
rect 32180 28160 32186 28172
rect 27798 28092 27804 28144
rect 27856 28132 27862 28144
rect 28261 28135 28319 28141
rect 28261 28132 28273 28135
rect 27856 28104 28273 28132
rect 27856 28092 27862 28104
rect 28261 28101 28273 28104
rect 28307 28132 28319 28135
rect 28534 28132 28540 28144
rect 28307 28104 28540 28132
rect 28307 28101 28319 28104
rect 28261 28095 28319 28101
rect 28534 28092 28540 28104
rect 28592 28092 28598 28144
rect 29730 28132 29736 28144
rect 29486 28104 29736 28132
rect 29730 28092 29736 28104
rect 29788 28132 29794 28144
rect 30190 28132 30196 28144
rect 29788 28104 30196 28132
rect 29788 28092 29794 28104
rect 30190 28092 30196 28104
rect 30248 28092 30254 28144
rect 32030 28132 32036 28144
rect 31726 28104 32036 28132
rect 29546 28024 29552 28076
rect 29604 28064 29610 28076
rect 31205 28067 31263 28073
rect 31205 28064 31217 28067
rect 29604 28036 31217 28064
rect 29604 28024 29610 28036
rect 31205 28033 31217 28036
rect 31251 28033 31263 28067
rect 31205 28027 31263 28033
rect 27614 27956 27620 28008
rect 27672 27996 27678 28008
rect 27985 27999 28043 28005
rect 27985 27996 27997 27999
rect 27672 27968 27997 27996
rect 27672 27956 27678 27968
rect 27985 27965 27997 27968
rect 28031 27965 28043 27999
rect 27985 27959 28043 27965
rect 24780 27832 26832 27860
rect 28000 27860 28028 27959
rect 29730 27956 29736 28008
rect 29788 27996 29794 28008
rect 30742 27996 30748 28008
rect 29788 27968 30748 27996
rect 29788 27956 29794 27968
rect 30742 27956 30748 27968
rect 30800 27956 30806 28008
rect 31297 27999 31355 28005
rect 31297 27965 31309 27999
rect 31343 27965 31355 27999
rect 31297 27959 31355 27965
rect 31481 27999 31539 28005
rect 31481 27965 31493 27999
rect 31527 27996 31539 27999
rect 31726 27996 31754 28104
rect 32030 28092 32036 28104
rect 32088 28092 32094 28144
rect 32600 28141 32628 28172
rect 33410 28160 33416 28172
rect 33468 28160 33474 28212
rect 35894 28160 35900 28212
rect 35952 28200 35958 28212
rect 36357 28203 36415 28209
rect 36357 28200 36369 28203
rect 35952 28172 36369 28200
rect 35952 28160 35958 28172
rect 36357 28169 36369 28172
rect 36403 28169 36415 28203
rect 36357 28163 36415 28169
rect 36538 28160 36544 28212
rect 36596 28200 36602 28212
rect 37461 28203 37519 28209
rect 37461 28200 37473 28203
rect 36596 28172 37473 28200
rect 36596 28160 36602 28172
rect 37461 28169 37473 28172
rect 37507 28169 37519 28203
rect 37461 28163 37519 28169
rect 37921 28203 37979 28209
rect 37921 28169 37933 28203
rect 37967 28200 37979 28203
rect 38654 28200 38660 28212
rect 37967 28172 38660 28200
rect 37967 28169 37979 28172
rect 37921 28163 37979 28169
rect 38654 28160 38660 28172
rect 38712 28160 38718 28212
rect 39022 28160 39028 28212
rect 39080 28160 39086 28212
rect 32585 28135 32643 28141
rect 32585 28101 32597 28135
rect 32631 28101 32643 28135
rect 33870 28132 33876 28144
rect 33810 28104 33876 28132
rect 32585 28095 32643 28101
rect 33870 28092 33876 28104
rect 33928 28132 33934 28144
rect 34790 28132 34796 28144
rect 33928 28104 34796 28132
rect 33928 28092 33934 28104
rect 34790 28092 34796 28104
rect 34848 28092 34854 28144
rect 36449 28135 36507 28141
rect 36449 28101 36461 28135
rect 36495 28132 36507 28135
rect 36814 28132 36820 28144
rect 36495 28104 36820 28132
rect 36495 28101 36507 28104
rect 36449 28095 36507 28101
rect 36814 28092 36820 28104
rect 36872 28092 36878 28144
rect 38580 28104 41414 28132
rect 37458 28024 37464 28076
rect 37516 28064 37522 28076
rect 37829 28067 37887 28073
rect 37516 28036 37780 28064
rect 37516 28024 37522 28036
rect 31527 27968 31754 27996
rect 31527 27965 31539 27968
rect 31481 27959 31539 27965
rect 30837 27931 30895 27937
rect 30837 27928 30849 27931
rect 29288 27900 30849 27928
rect 28442 27860 28448 27872
rect 28000 27832 28448 27860
rect 28442 27820 28448 27832
rect 28500 27820 28506 27872
rect 28626 27820 28632 27872
rect 28684 27860 28690 27872
rect 29288 27860 29316 27900
rect 30837 27897 30849 27900
rect 30883 27897 30895 27931
rect 30837 27891 30895 27897
rect 28684 27832 29316 27860
rect 29733 27863 29791 27869
rect 28684 27820 28690 27832
rect 29733 27829 29745 27863
rect 29779 27860 29791 27863
rect 29822 27860 29828 27872
rect 29779 27832 29828 27860
rect 29779 27829 29791 27832
rect 29733 27823 29791 27829
rect 29822 27820 29828 27832
rect 29880 27820 29886 27872
rect 31312 27860 31340 27959
rect 32306 27956 32312 28008
rect 32364 27956 32370 28008
rect 34514 27996 34520 28008
rect 32416 27968 34520 27996
rect 32416 27860 32444 27968
rect 34514 27956 34520 27968
rect 34572 27956 34578 28008
rect 36633 27999 36691 28005
rect 36633 27965 36645 27999
rect 36679 27996 36691 27999
rect 37642 27996 37648 28008
rect 36679 27968 37648 27996
rect 36679 27965 36691 27968
rect 36633 27959 36691 27965
rect 37642 27956 37648 27968
rect 37700 27956 37706 28008
rect 37752 27996 37780 28036
rect 37829 28033 37841 28067
rect 37875 28064 37887 28067
rect 38470 28064 38476 28076
rect 37875 28036 38476 28064
rect 37875 28033 37887 28036
rect 37829 28027 37887 28033
rect 38470 28024 38476 28036
rect 38528 28024 38534 28076
rect 38013 27999 38071 28005
rect 38013 27996 38025 27999
rect 37752 27968 38025 27996
rect 38013 27965 38025 27968
rect 38059 27996 38071 27999
rect 38580 27996 38608 28104
rect 38654 28024 38660 28076
rect 38712 28064 38718 28076
rect 39482 28064 39488 28076
rect 38712 28036 39488 28064
rect 38712 28024 38718 28036
rect 39482 28024 39488 28036
rect 39540 28024 39546 28076
rect 41386 28064 41414 28104
rect 46934 28092 46940 28144
rect 46992 28132 46998 28144
rect 48041 28135 48099 28141
rect 48041 28132 48053 28135
rect 46992 28104 48053 28132
rect 46992 28092 46998 28104
rect 48041 28101 48053 28104
rect 48087 28101 48099 28135
rect 48041 28095 48099 28101
rect 41598 28064 41604 28076
rect 41386 28036 41604 28064
rect 41598 28024 41604 28036
rect 41656 28024 41662 28076
rect 38059 27968 38608 27996
rect 38059 27965 38071 27968
rect 38013 27959 38071 27965
rect 39114 27956 39120 28008
rect 39172 27956 39178 28008
rect 39301 27999 39359 28005
rect 39301 27965 39313 27999
rect 39347 27996 39359 27999
rect 40494 27996 40500 28008
rect 39347 27968 40500 27996
rect 39347 27965 39359 27968
rect 39301 27959 39359 27965
rect 40494 27956 40500 27968
rect 40552 27956 40558 28008
rect 33778 27888 33784 27940
rect 33836 27928 33842 27940
rect 38378 27928 38384 27940
rect 33836 27900 38384 27928
rect 33836 27888 33842 27900
rect 38378 27888 38384 27900
rect 38436 27888 38442 27940
rect 38657 27931 38715 27937
rect 38657 27897 38669 27931
rect 38703 27928 38715 27931
rect 41138 27928 41144 27940
rect 38703 27900 41144 27928
rect 38703 27897 38715 27900
rect 38657 27891 38715 27897
rect 41138 27888 41144 27900
rect 41196 27888 41202 27940
rect 31312 27832 32444 27860
rect 32582 27820 32588 27872
rect 32640 27860 32646 27872
rect 34057 27863 34115 27869
rect 34057 27860 34069 27863
rect 32640 27832 34069 27860
rect 32640 27820 32646 27832
rect 34057 27829 34069 27832
rect 34103 27860 34115 27863
rect 34146 27860 34152 27872
rect 34103 27832 34152 27860
rect 34103 27829 34115 27832
rect 34057 27823 34115 27829
rect 34146 27820 34152 27832
rect 34204 27820 34210 27872
rect 35158 27820 35164 27872
rect 35216 27860 35222 27872
rect 35434 27860 35440 27872
rect 35216 27832 35440 27860
rect 35216 27820 35222 27832
rect 35434 27820 35440 27832
rect 35492 27820 35498 27872
rect 35986 27820 35992 27872
rect 36044 27820 36050 27872
rect 37182 27820 37188 27872
rect 37240 27860 37246 27872
rect 41230 27860 41236 27872
rect 37240 27832 41236 27860
rect 37240 27820 37246 27832
rect 41230 27820 41236 27832
rect 41288 27820 41294 27872
rect 47762 27820 47768 27872
rect 47820 27860 47826 27872
rect 48133 27863 48191 27869
rect 48133 27860 48145 27863
rect 47820 27832 48145 27860
rect 47820 27820 47826 27832
rect 48133 27829 48145 27832
rect 48179 27829 48191 27863
rect 48133 27823 48191 27829
rect 1104 27770 49864 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 32950 27770
rect 33002 27718 33014 27770
rect 33066 27718 33078 27770
rect 33130 27718 33142 27770
rect 33194 27718 33206 27770
rect 33258 27718 42950 27770
rect 43002 27718 43014 27770
rect 43066 27718 43078 27770
rect 43130 27718 43142 27770
rect 43194 27718 43206 27770
rect 43258 27718 49864 27770
rect 1104 27696 49864 27718
rect 28350 27616 28356 27668
rect 28408 27656 28414 27668
rect 30650 27656 30656 27668
rect 28408 27628 30656 27656
rect 28408 27616 28414 27628
rect 30650 27616 30656 27628
rect 30708 27616 30714 27668
rect 30742 27616 30748 27668
rect 30800 27656 30806 27668
rect 39114 27656 39120 27668
rect 30800 27628 39120 27656
rect 30800 27616 30806 27628
rect 39114 27616 39120 27628
rect 39172 27616 39178 27668
rect 40300 27659 40358 27665
rect 40300 27625 40312 27659
rect 40346 27656 40358 27659
rect 40770 27656 40776 27668
rect 40346 27628 40776 27656
rect 40346 27625 40358 27628
rect 40300 27619 40358 27625
rect 40770 27616 40776 27628
rect 40828 27616 40834 27668
rect 7650 27548 7656 27600
rect 7708 27588 7714 27600
rect 7791 27591 7849 27597
rect 7791 27588 7803 27591
rect 7708 27560 7803 27588
rect 7708 27548 7714 27560
rect 7791 27557 7803 27560
rect 7837 27557 7849 27591
rect 7791 27551 7849 27557
rect 27617 27591 27675 27597
rect 27617 27557 27629 27591
rect 27663 27588 27675 27591
rect 29546 27588 29552 27600
rect 27663 27560 29552 27588
rect 27663 27557 27675 27560
rect 27617 27551 27675 27557
rect 29546 27548 29552 27560
rect 29604 27548 29610 27600
rect 30668 27588 30696 27616
rect 30668 27560 31754 27588
rect 1302 27480 1308 27532
rect 1360 27520 1366 27532
rect 2041 27523 2099 27529
rect 2041 27520 2053 27523
rect 1360 27492 2053 27520
rect 1360 27480 1366 27492
rect 2041 27489 2053 27492
rect 2087 27489 2099 27523
rect 2041 27483 2099 27489
rect 24946 27480 24952 27532
rect 25004 27480 25010 27532
rect 28261 27523 28319 27529
rect 28261 27489 28273 27523
rect 28307 27520 28319 27523
rect 30282 27520 30288 27532
rect 28307 27492 30288 27520
rect 28307 27489 28319 27492
rect 28261 27483 28319 27489
rect 30282 27480 30288 27492
rect 30340 27480 30346 27532
rect 30745 27523 30803 27529
rect 30745 27520 30757 27523
rect 30484 27492 30757 27520
rect 1765 27455 1823 27461
rect 1765 27421 1777 27455
rect 1811 27452 1823 27455
rect 4982 27452 4988 27464
rect 1811 27424 4988 27452
rect 1811 27421 1823 27424
rect 1765 27415 1823 27421
rect 4982 27412 4988 27424
rect 5040 27412 5046 27464
rect 7720 27455 7778 27461
rect 7720 27452 7732 27455
rect 6886 27424 7732 27452
rect 4890 27344 4896 27396
rect 4948 27384 4954 27396
rect 6886 27384 6914 27424
rect 7720 27421 7732 27424
rect 7766 27452 7778 27455
rect 9766 27452 9772 27464
rect 7766 27424 9772 27452
rect 7766 27421 7778 27424
rect 7720 27415 7778 27421
rect 9766 27412 9772 27424
rect 9824 27412 9830 27464
rect 23106 27412 23112 27464
rect 23164 27452 23170 27464
rect 23385 27455 23443 27461
rect 23385 27452 23397 27455
rect 23164 27424 23397 27452
rect 23164 27412 23170 27424
rect 23385 27421 23397 27424
rect 23431 27421 23443 27455
rect 23385 27415 23443 27421
rect 27985 27455 28043 27461
rect 27985 27421 27997 27455
rect 28031 27452 28043 27455
rect 29914 27452 29920 27464
rect 28031 27424 29920 27452
rect 28031 27421 28043 27424
rect 27985 27415 28043 27421
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 4948 27356 6914 27384
rect 4948 27344 4954 27356
rect 25222 27344 25228 27396
rect 25280 27344 25286 27396
rect 26234 27344 26240 27396
rect 26292 27344 26298 27396
rect 27614 27344 27620 27396
rect 27672 27384 27678 27396
rect 30484 27384 30512 27492
rect 30745 27489 30757 27492
rect 30791 27489 30803 27523
rect 30745 27483 30803 27489
rect 31726 27452 31754 27560
rect 32766 27548 32772 27600
rect 32824 27588 32830 27600
rect 32824 27560 35664 27588
rect 32824 27548 32830 27560
rect 32030 27480 32036 27532
rect 32088 27520 32094 27532
rect 32214 27520 32220 27532
rect 32088 27492 32220 27520
rect 32088 27480 32094 27492
rect 32214 27480 32220 27492
rect 32272 27520 32278 27532
rect 32309 27523 32367 27529
rect 32309 27520 32321 27523
rect 32272 27492 32321 27520
rect 32272 27480 32278 27492
rect 32309 27489 32321 27492
rect 32355 27489 32367 27523
rect 32309 27483 32367 27489
rect 35342 27480 35348 27532
rect 35400 27480 35406 27532
rect 35526 27480 35532 27532
rect 35584 27480 35590 27532
rect 35636 27520 35664 27560
rect 41598 27548 41604 27600
rect 41656 27588 41662 27600
rect 41785 27591 41843 27597
rect 41785 27588 41797 27591
rect 41656 27560 41797 27588
rect 41656 27548 41662 27560
rect 41785 27557 41797 27560
rect 41831 27557 41843 27591
rect 41785 27551 41843 27557
rect 40037 27523 40095 27529
rect 35636 27492 38516 27520
rect 32953 27455 33011 27461
rect 32953 27452 32965 27455
rect 31726 27424 32965 27452
rect 32953 27421 32965 27424
rect 32999 27452 33011 27455
rect 34882 27452 34888 27464
rect 32999 27424 34888 27452
rect 32999 27421 33011 27424
rect 32953 27415 33011 27421
rect 34882 27412 34888 27424
rect 34940 27412 34946 27464
rect 35253 27455 35311 27461
rect 35253 27421 35265 27455
rect 35299 27452 35311 27455
rect 36078 27452 36084 27464
rect 35299 27424 36084 27452
rect 35299 27421 35311 27424
rect 35253 27415 35311 27421
rect 36078 27412 36084 27424
rect 36136 27412 36142 27464
rect 37001 27455 37059 27461
rect 37001 27421 37013 27455
rect 37047 27421 37059 27455
rect 38488 27452 38516 27492
rect 40037 27489 40049 27523
rect 40083 27520 40095 27523
rect 40310 27520 40316 27532
rect 40083 27492 40316 27520
rect 40083 27489 40095 27492
rect 40037 27483 40095 27489
rect 40310 27480 40316 27492
rect 40368 27480 40374 27532
rect 47118 27520 47124 27532
rect 41616 27492 47124 27520
rect 38488 27424 38608 27452
rect 37001 27415 37059 27421
rect 27672 27356 30512 27384
rect 30561 27387 30619 27393
rect 27672 27344 27678 27356
rect 30561 27353 30573 27387
rect 30607 27384 30619 27387
rect 31478 27384 31484 27396
rect 30607 27356 31484 27384
rect 30607 27353 30619 27356
rect 30561 27347 30619 27353
rect 31478 27344 31484 27356
rect 31536 27344 31542 27396
rect 32125 27387 32183 27393
rect 32125 27384 32137 27387
rect 31588 27356 32137 27384
rect 26694 27276 26700 27328
rect 26752 27316 26758 27328
rect 27246 27316 27252 27328
rect 26752 27288 27252 27316
rect 26752 27276 26758 27288
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 28077 27319 28135 27325
rect 28077 27285 28089 27319
rect 28123 27316 28135 27319
rect 28534 27316 28540 27328
rect 28123 27288 28540 27316
rect 28123 27285 28135 27288
rect 28077 27279 28135 27285
rect 28534 27276 28540 27288
rect 28592 27276 28598 27328
rect 30190 27276 30196 27328
rect 30248 27276 30254 27328
rect 30650 27276 30656 27328
rect 30708 27276 30714 27328
rect 30742 27276 30748 27328
rect 30800 27316 30806 27328
rect 31588 27316 31616 27356
rect 32125 27353 32137 27356
rect 32171 27353 32183 27387
rect 32125 27347 32183 27353
rect 32306 27344 32312 27396
rect 32364 27384 32370 27396
rect 33781 27387 33839 27393
rect 33781 27384 33793 27387
rect 32364 27356 33793 27384
rect 32364 27344 32370 27356
rect 33781 27353 33793 27356
rect 33827 27384 33839 27387
rect 33962 27384 33968 27396
rect 33827 27356 33968 27384
rect 33827 27353 33839 27356
rect 33781 27347 33839 27353
rect 33962 27344 33968 27356
rect 34020 27384 34026 27396
rect 37016 27384 37044 27415
rect 34020 27356 37044 27384
rect 34020 27344 34026 27356
rect 37182 27344 37188 27396
rect 37240 27384 37246 27396
rect 37277 27387 37335 27393
rect 37277 27384 37289 27387
rect 37240 27356 37289 27384
rect 37240 27344 37246 27356
rect 37277 27353 37289 27356
rect 37323 27353 37335 27387
rect 37277 27347 37335 27353
rect 37918 27344 37924 27396
rect 37976 27344 37982 27396
rect 38580 27384 38608 27424
rect 41414 27412 41420 27464
rect 41472 27412 41478 27464
rect 38580 27356 40632 27384
rect 30800 27288 31616 27316
rect 30800 27276 30806 27288
rect 31754 27276 31760 27328
rect 31812 27276 31818 27328
rect 32217 27319 32275 27325
rect 32217 27285 32229 27319
rect 32263 27316 32275 27319
rect 32582 27316 32588 27328
rect 32263 27288 32588 27316
rect 32263 27285 32275 27288
rect 32217 27279 32275 27285
rect 32582 27276 32588 27288
rect 32640 27276 32646 27328
rect 34790 27276 34796 27328
rect 34848 27316 34854 27328
rect 34885 27319 34943 27325
rect 34885 27316 34897 27319
rect 34848 27288 34897 27316
rect 34848 27276 34854 27288
rect 34885 27285 34897 27288
rect 34931 27285 34943 27319
rect 34885 27279 34943 27285
rect 35894 27276 35900 27328
rect 35952 27316 35958 27328
rect 36078 27316 36084 27328
rect 35952 27288 36084 27316
rect 35952 27276 35958 27288
rect 36078 27276 36084 27288
rect 36136 27316 36142 27328
rect 37200 27316 37228 27344
rect 36136 27288 37228 27316
rect 36136 27276 36142 27288
rect 38286 27276 38292 27328
rect 38344 27316 38350 27328
rect 38749 27319 38807 27325
rect 38749 27316 38761 27319
rect 38344 27288 38761 27316
rect 38344 27276 38350 27288
rect 38749 27285 38761 27288
rect 38795 27285 38807 27319
rect 40604 27316 40632 27356
rect 41616 27316 41644 27492
rect 47118 27480 47124 27492
rect 47176 27480 47182 27532
rect 44174 27412 44180 27464
rect 44232 27412 44238 27464
rect 47210 27412 47216 27464
rect 47268 27412 47274 27464
rect 48498 27412 48504 27464
rect 48556 27412 48562 27464
rect 48777 27455 48835 27461
rect 48777 27421 48789 27455
rect 48823 27421 48835 27455
rect 48777 27415 48835 27421
rect 47397 27387 47455 27393
rect 47397 27353 47409 27387
rect 47443 27384 47455 27387
rect 47578 27384 47584 27396
rect 47443 27356 47584 27384
rect 47443 27353 47455 27356
rect 47397 27347 47455 27353
rect 47578 27344 47584 27356
rect 47636 27344 47642 27396
rect 47670 27344 47676 27396
rect 47728 27384 47734 27396
rect 48792 27384 48820 27415
rect 47728 27356 48820 27384
rect 47728 27344 47734 27356
rect 40604 27288 41644 27316
rect 38749 27279 38807 27285
rect 43990 27276 43996 27328
rect 44048 27276 44054 27328
rect 1104 27226 49864 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 27950 27226
rect 28002 27174 28014 27226
rect 28066 27174 28078 27226
rect 28130 27174 28142 27226
rect 28194 27174 28206 27226
rect 28258 27174 37950 27226
rect 38002 27174 38014 27226
rect 38066 27174 38078 27226
rect 38130 27174 38142 27226
rect 38194 27174 38206 27226
rect 38258 27174 47950 27226
rect 48002 27174 48014 27226
rect 48066 27174 48078 27226
rect 48130 27174 48142 27226
rect 48194 27174 48206 27226
rect 48258 27174 49864 27226
rect 1104 27152 49864 27174
rect 23106 27072 23112 27124
rect 23164 27072 23170 27124
rect 26694 27072 26700 27124
rect 26752 27112 26758 27124
rect 27154 27112 27160 27124
rect 26752 27084 27160 27112
rect 26752 27072 26758 27084
rect 27154 27072 27160 27084
rect 27212 27112 27218 27124
rect 30650 27112 30656 27124
rect 27212 27084 30656 27112
rect 27212 27072 27218 27084
rect 30650 27072 30656 27084
rect 30708 27072 30714 27124
rect 30834 27072 30840 27124
rect 30892 27112 30898 27124
rect 31113 27115 31171 27121
rect 31113 27112 31125 27115
rect 30892 27084 31125 27112
rect 30892 27072 30898 27084
rect 31113 27081 31125 27084
rect 31159 27112 31171 27115
rect 31202 27112 31208 27124
rect 31159 27084 31208 27112
rect 31159 27081 31171 27084
rect 31113 27075 31171 27081
rect 31202 27072 31208 27084
rect 31260 27072 31266 27124
rect 31846 27072 31852 27124
rect 31904 27112 31910 27124
rect 31904 27084 36952 27112
rect 31904 27072 31910 27084
rect 22554 27004 22560 27056
rect 22612 27044 22618 27056
rect 23201 27047 23259 27053
rect 23201 27044 23213 27047
rect 22612 27016 23213 27044
rect 22612 27004 22618 27016
rect 23201 27013 23213 27016
rect 23247 27013 23259 27047
rect 23201 27007 23259 27013
rect 24121 27047 24179 27053
rect 24121 27013 24133 27047
rect 24167 27044 24179 27047
rect 25866 27044 25872 27056
rect 24167 27016 25872 27044
rect 24167 27013 24179 27016
rect 24121 27007 24179 27013
rect 25866 27004 25872 27016
rect 25924 27004 25930 27056
rect 33870 27004 33876 27056
rect 33928 27044 33934 27056
rect 34517 27047 34575 27053
rect 34517 27044 34529 27047
rect 33928 27016 34529 27044
rect 33928 27004 33934 27016
rect 34517 27013 34529 27016
rect 34563 27013 34575 27047
rect 34517 27007 34575 27013
rect 34974 27004 34980 27056
rect 35032 27004 35038 27056
rect 7834 26936 7840 26988
rect 7892 26936 7898 26988
rect 30282 26976 30288 26988
rect 29946 26948 30288 26976
rect 30282 26936 30288 26948
rect 30340 26936 30346 26988
rect 31294 26936 31300 26988
rect 31352 26976 31358 26988
rect 36924 26985 36952 27084
rect 37090 27072 37096 27124
rect 37148 27112 37154 27124
rect 40586 27112 40592 27124
rect 37148 27084 40592 27112
rect 37148 27072 37154 27084
rect 40586 27072 40592 27084
rect 40644 27072 40650 27124
rect 40678 27072 40684 27124
rect 40736 27112 40742 27124
rect 42061 27115 42119 27121
rect 42061 27112 42073 27115
rect 40736 27084 42073 27112
rect 40736 27072 40742 27084
rect 42061 27081 42073 27084
rect 42107 27081 42119 27115
rect 42061 27075 42119 27081
rect 42150 27072 42156 27124
rect 42208 27112 42214 27124
rect 48774 27112 48780 27124
rect 42208 27084 48780 27112
rect 42208 27072 42214 27084
rect 48774 27072 48780 27084
rect 48832 27072 48838 27124
rect 38565 27047 38623 27053
rect 38565 27013 38577 27047
rect 38611 27044 38623 27047
rect 38611 27016 39896 27044
rect 38611 27013 38623 27016
rect 38565 27007 38623 27013
rect 39868 26988 39896 27016
rect 41598 27004 41604 27056
rect 41656 27004 41662 27056
rect 44818 27004 44824 27056
rect 44876 27044 44882 27056
rect 47857 27047 47915 27053
rect 47857 27044 47869 27047
rect 44876 27016 47869 27044
rect 44876 27004 44882 27016
rect 47857 27013 47869 27016
rect 47903 27013 47915 27047
rect 47857 27007 47915 27013
rect 33413 26979 33471 26985
rect 33413 26976 33425 26979
rect 31352 26948 33425 26976
rect 31352 26936 31358 26948
rect 33413 26945 33425 26948
rect 33459 26945 33471 26979
rect 33413 26939 33471 26945
rect 36909 26979 36967 26985
rect 36909 26945 36921 26979
rect 36955 26945 36967 26979
rect 36909 26939 36967 26945
rect 37734 26936 37740 26988
rect 37792 26936 37798 26988
rect 39850 26936 39856 26988
rect 39908 26976 39914 26988
rect 40310 26976 40316 26988
rect 40368 26985 40374 26988
rect 39908 26948 40316 26976
rect 39908 26936 39914 26948
rect 40310 26936 40316 26948
rect 40368 26939 40378 26985
rect 40368 26936 40374 26939
rect 47026 26936 47032 26988
rect 47084 26936 47090 26988
rect 47118 26936 47124 26988
rect 47176 26976 47182 26988
rect 48777 26979 48835 26985
rect 48777 26976 48789 26979
rect 47176 26948 48789 26976
rect 47176 26936 47182 26948
rect 48777 26945 48789 26948
rect 48823 26945 48835 26979
rect 48777 26939 48835 26945
rect 8021 26911 8079 26917
rect 8021 26877 8033 26911
rect 8067 26908 8079 26911
rect 8294 26908 8300 26920
rect 8067 26880 8300 26908
rect 8067 26877 8079 26880
rect 8021 26871 8079 26877
rect 8294 26868 8300 26880
rect 8352 26868 8358 26920
rect 9582 26868 9588 26920
rect 9640 26868 9646 26920
rect 23382 26868 23388 26920
rect 23440 26868 23446 26920
rect 28442 26868 28448 26920
rect 28500 26908 28506 26920
rect 28537 26911 28595 26917
rect 28537 26908 28549 26911
rect 28500 26880 28549 26908
rect 28500 26868 28506 26880
rect 28537 26877 28549 26880
rect 28583 26877 28595 26911
rect 28537 26871 28595 26877
rect 28813 26911 28871 26917
rect 28813 26877 28825 26911
rect 28859 26908 28871 26911
rect 29822 26908 29828 26920
rect 28859 26880 29828 26908
rect 28859 26877 28871 26880
rect 28813 26871 28871 26877
rect 29822 26868 29828 26880
rect 29880 26908 29886 26920
rect 29880 26880 29960 26908
rect 29880 26868 29886 26880
rect 22741 26843 22799 26849
rect 22741 26809 22753 26843
rect 22787 26840 22799 26843
rect 28166 26840 28172 26852
rect 22787 26812 28172 26840
rect 22787 26809 22799 26812
rect 22741 26803 22799 26809
rect 28166 26800 28172 26812
rect 28224 26800 28230 26852
rect 29932 26840 29960 26880
rect 31018 26868 31024 26920
rect 31076 26908 31082 26920
rect 31205 26911 31263 26917
rect 31205 26908 31217 26911
rect 31076 26880 31217 26908
rect 31076 26868 31082 26880
rect 31205 26877 31217 26880
rect 31251 26877 31263 26911
rect 31205 26871 31263 26877
rect 31386 26868 31392 26920
rect 31444 26868 31450 26920
rect 33226 26868 33232 26920
rect 33284 26908 33290 26920
rect 33505 26911 33563 26917
rect 33505 26908 33517 26911
rect 33284 26880 33517 26908
rect 33284 26868 33290 26880
rect 33505 26877 33517 26880
rect 33551 26877 33563 26911
rect 33505 26871 33563 26877
rect 33689 26911 33747 26917
rect 33689 26877 33701 26911
rect 33735 26908 33747 26911
rect 34054 26908 34060 26920
rect 33735 26880 34060 26908
rect 33735 26877 33747 26880
rect 33689 26871 33747 26877
rect 34054 26868 34060 26880
rect 34112 26868 34118 26920
rect 34248 26911 34306 26917
rect 34248 26877 34260 26911
rect 34294 26877 34306 26911
rect 34248 26871 34306 26877
rect 29932 26812 31340 26840
rect 31312 26784 31340 26812
rect 31478 26800 31484 26852
rect 31536 26840 31542 26852
rect 34146 26840 34152 26852
rect 31536 26812 34152 26840
rect 31536 26800 31542 26812
rect 34146 26800 34152 26812
rect 34204 26800 34210 26852
rect 24026 26732 24032 26784
rect 24084 26772 24090 26784
rect 24213 26775 24271 26781
rect 24213 26772 24225 26775
rect 24084 26744 24225 26772
rect 24084 26732 24090 26744
rect 24213 26741 24225 26744
rect 24259 26741 24271 26775
rect 24213 26735 24271 26741
rect 26970 26732 26976 26784
rect 27028 26772 27034 26784
rect 27341 26775 27399 26781
rect 27341 26772 27353 26775
rect 27028 26744 27353 26772
rect 27028 26732 27034 26744
rect 27341 26741 27353 26744
rect 27387 26741 27399 26775
rect 27341 26735 27399 26741
rect 30098 26732 30104 26784
rect 30156 26772 30162 26784
rect 30285 26775 30343 26781
rect 30285 26772 30297 26775
rect 30156 26744 30297 26772
rect 30156 26732 30162 26744
rect 30285 26741 30297 26744
rect 30331 26741 30343 26775
rect 30285 26735 30343 26741
rect 30374 26732 30380 26784
rect 30432 26772 30438 26784
rect 30745 26775 30803 26781
rect 30745 26772 30757 26775
rect 30432 26744 30757 26772
rect 30432 26732 30438 26744
rect 30745 26741 30757 26744
rect 30791 26741 30803 26775
rect 30745 26735 30803 26741
rect 31294 26732 31300 26784
rect 31352 26732 31358 26784
rect 33045 26775 33103 26781
rect 33045 26741 33057 26775
rect 33091 26772 33103 26775
rect 33962 26772 33968 26784
rect 33091 26744 33968 26772
rect 33091 26741 33103 26744
rect 33045 26735 33103 26741
rect 33962 26732 33968 26744
rect 34020 26732 34026 26784
rect 34256 26772 34284 26871
rect 40126 26868 40132 26920
rect 40184 26908 40190 26920
rect 40589 26911 40647 26917
rect 40589 26908 40601 26911
rect 40184 26880 40601 26908
rect 40184 26868 40190 26880
rect 40589 26877 40601 26880
rect 40635 26877 40647 26911
rect 47670 26908 47676 26920
rect 40589 26871 40647 26877
rect 41616 26880 47676 26908
rect 35802 26800 35808 26852
rect 35860 26840 35866 26852
rect 35860 26812 40448 26840
rect 35860 26800 35866 26812
rect 34974 26772 34980 26784
rect 34256 26744 34980 26772
rect 34974 26732 34980 26744
rect 35032 26732 35038 26784
rect 35989 26775 36047 26781
rect 35989 26741 36001 26775
rect 36035 26772 36047 26775
rect 36078 26772 36084 26784
rect 36035 26744 36084 26772
rect 36035 26741 36047 26744
rect 35989 26735 36047 26741
rect 36078 26732 36084 26744
rect 36136 26732 36142 26784
rect 36725 26775 36783 26781
rect 36725 26741 36737 26775
rect 36771 26772 36783 26775
rect 39022 26772 39028 26784
rect 36771 26744 39028 26772
rect 36771 26741 36783 26744
rect 36725 26735 36783 26741
rect 39022 26732 39028 26744
rect 39080 26732 39086 26784
rect 40420 26772 40448 26812
rect 41616 26772 41644 26880
rect 47670 26868 47676 26880
rect 47728 26868 47734 26920
rect 48498 26868 48504 26920
rect 48556 26868 48562 26920
rect 40420 26744 41644 26772
rect 46750 26732 46756 26784
rect 46808 26772 46814 26784
rect 46845 26775 46903 26781
rect 46845 26772 46857 26775
rect 46808 26744 46857 26772
rect 46808 26732 46814 26744
rect 46845 26741 46857 26744
rect 46891 26741 46903 26775
rect 46845 26735 46903 26741
rect 47670 26732 47676 26784
rect 47728 26772 47734 26784
rect 47949 26775 48007 26781
rect 47949 26772 47961 26775
rect 47728 26744 47961 26772
rect 47728 26732 47734 26744
rect 47949 26741 47961 26744
rect 47995 26741 48007 26775
rect 47949 26735 48007 26741
rect 1104 26682 49864 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 32950 26682
rect 33002 26630 33014 26682
rect 33066 26630 33078 26682
rect 33130 26630 33142 26682
rect 33194 26630 33206 26682
rect 33258 26630 42950 26682
rect 43002 26630 43014 26682
rect 43066 26630 43078 26682
rect 43130 26630 43142 26682
rect 43194 26630 43206 26682
rect 43258 26630 49864 26682
rect 1104 26608 49864 26630
rect 7742 26528 7748 26580
rect 7800 26568 7806 26580
rect 7883 26571 7941 26577
rect 7883 26568 7895 26571
rect 7800 26540 7895 26568
rect 7800 26528 7806 26540
rect 7883 26537 7895 26540
rect 7929 26537 7941 26571
rect 7883 26531 7941 26537
rect 9674 26528 9680 26580
rect 9732 26528 9738 26580
rect 25038 26528 25044 26580
rect 25096 26568 25102 26580
rect 25314 26568 25320 26580
rect 25096 26540 25320 26568
rect 25096 26528 25102 26540
rect 25314 26528 25320 26540
rect 25372 26568 25378 26580
rect 25774 26568 25780 26580
rect 25372 26540 25780 26568
rect 25372 26528 25378 26540
rect 25774 26528 25780 26540
rect 25832 26528 25838 26580
rect 27154 26528 27160 26580
rect 27212 26568 27218 26580
rect 27798 26568 27804 26580
rect 27212 26540 27804 26568
rect 27212 26528 27218 26540
rect 27798 26528 27804 26540
rect 27856 26528 27862 26580
rect 30745 26571 30803 26577
rect 30745 26537 30757 26571
rect 30791 26568 30803 26571
rect 35526 26568 35532 26580
rect 30791 26540 35532 26568
rect 30791 26537 30803 26540
rect 30745 26531 30803 26537
rect 35526 26528 35532 26540
rect 35584 26528 35590 26580
rect 40126 26528 40132 26580
rect 40184 26568 40190 26580
rect 41782 26568 41788 26580
rect 40184 26540 41788 26568
rect 40184 26528 40190 26540
rect 41782 26528 41788 26540
rect 41840 26528 41846 26580
rect 23750 26460 23756 26512
rect 23808 26500 23814 26512
rect 23845 26503 23903 26509
rect 23845 26500 23857 26503
rect 23808 26472 23857 26500
rect 23808 26460 23814 26472
rect 23845 26469 23857 26472
rect 23891 26469 23903 26503
rect 23845 26463 23903 26469
rect 24210 26460 24216 26512
rect 24268 26500 24274 26512
rect 26605 26503 26663 26509
rect 24268 26472 25268 26500
rect 24268 26460 24274 26472
rect 9125 26435 9183 26441
rect 9125 26401 9137 26435
rect 9171 26432 9183 26435
rect 10870 26432 10876 26444
rect 9171 26404 10876 26432
rect 9171 26401 9183 26404
rect 9125 26395 9183 26401
rect 10870 26392 10876 26404
rect 10928 26392 10934 26444
rect 22094 26392 22100 26444
rect 22152 26392 22158 26444
rect 22373 26435 22431 26441
rect 22373 26401 22385 26435
rect 22419 26432 22431 26435
rect 24228 26432 24256 26460
rect 22419 26404 24256 26432
rect 22419 26401 22431 26404
rect 22373 26395 22431 26401
rect 25038 26392 25044 26444
rect 25096 26392 25102 26444
rect 25133 26435 25191 26441
rect 25133 26401 25145 26435
rect 25179 26401 25191 26435
rect 25240 26432 25268 26472
rect 26605 26469 26617 26503
rect 26651 26500 26663 26503
rect 26651 26472 31156 26500
rect 26651 26469 26663 26472
rect 26605 26463 26663 26469
rect 25240 26404 27108 26432
rect 25133 26395 25191 26401
rect 7742 26324 7748 26376
rect 7800 26373 7806 26376
rect 7800 26367 7838 26373
rect 7826 26333 7838 26367
rect 7800 26327 7838 26333
rect 9309 26367 9367 26373
rect 9309 26333 9321 26367
rect 9355 26364 9367 26367
rect 9766 26364 9772 26376
rect 9355 26336 9772 26364
rect 9355 26333 9367 26336
rect 9309 26327 9367 26333
rect 7800 26324 7806 26327
rect 9766 26324 9772 26336
rect 9824 26364 9830 26376
rect 10962 26364 10968 26376
rect 9824 26336 10968 26364
rect 9824 26324 9830 26336
rect 10962 26324 10968 26336
rect 11020 26324 11026 26376
rect 23750 26324 23756 26376
rect 23808 26364 23814 26376
rect 25148 26364 25176 26395
rect 23808 26336 25176 26364
rect 23808 26324 23814 26336
rect 26970 26324 26976 26376
rect 27028 26324 27034 26376
rect 27080 26364 27108 26404
rect 27154 26392 27160 26444
rect 27212 26392 27218 26444
rect 28353 26435 28411 26441
rect 28353 26432 28365 26435
rect 27264 26404 28365 26432
rect 27264 26364 27292 26404
rect 28353 26401 28365 26404
rect 28399 26401 28411 26435
rect 28353 26395 28411 26401
rect 29362 26392 29368 26444
rect 29420 26432 29426 26444
rect 30742 26432 30748 26444
rect 29420 26404 30748 26432
rect 29420 26392 29426 26404
rect 30742 26392 30748 26404
rect 30800 26392 30806 26444
rect 27080 26336 27292 26364
rect 28166 26324 28172 26376
rect 28224 26324 28230 26376
rect 28261 26367 28319 26373
rect 28261 26333 28273 26367
rect 28307 26364 28319 26367
rect 28902 26364 28908 26376
rect 28307 26336 28908 26364
rect 28307 26333 28319 26336
rect 28261 26327 28319 26333
rect 28902 26324 28908 26336
rect 28960 26324 28966 26376
rect 29086 26324 29092 26376
rect 29144 26364 29150 26376
rect 31018 26364 31024 26376
rect 29144 26336 31024 26364
rect 29144 26324 29150 26336
rect 31018 26324 31024 26336
rect 31076 26324 31082 26376
rect 31128 26373 31156 26472
rect 38378 26460 38384 26512
rect 38436 26500 38442 26512
rect 38749 26503 38807 26509
rect 38749 26500 38761 26503
rect 38436 26472 38761 26500
rect 38436 26460 38442 26472
rect 38749 26469 38761 26472
rect 38795 26469 38807 26503
rect 38749 26463 38807 26469
rect 39022 26460 39028 26512
rect 39080 26500 39086 26512
rect 39080 26472 40172 26500
rect 39080 26460 39086 26472
rect 31202 26392 31208 26444
rect 31260 26392 31266 26444
rect 31294 26392 31300 26444
rect 31352 26392 31358 26444
rect 31846 26392 31852 26444
rect 31904 26432 31910 26444
rect 32030 26432 32036 26444
rect 31904 26404 32036 26432
rect 31904 26392 31910 26404
rect 32030 26392 32036 26404
rect 32088 26392 32094 26444
rect 32214 26392 32220 26444
rect 32272 26392 32278 26444
rect 33870 26392 33876 26444
rect 33928 26432 33934 26444
rect 33965 26435 34023 26441
rect 33965 26432 33977 26435
rect 33928 26404 33977 26432
rect 33928 26392 33934 26404
rect 33965 26401 33977 26404
rect 34011 26401 34023 26435
rect 33965 26395 34023 26401
rect 35986 26392 35992 26444
rect 36044 26432 36050 26444
rect 39209 26435 39267 26441
rect 39209 26432 39221 26435
rect 36044 26404 39221 26432
rect 36044 26392 36050 26404
rect 39209 26401 39221 26404
rect 39255 26401 39267 26435
rect 39209 26395 39267 26401
rect 39390 26392 39396 26444
rect 39448 26392 39454 26444
rect 39850 26392 39856 26444
rect 39908 26432 39914 26444
rect 40037 26435 40095 26441
rect 40037 26432 40049 26435
rect 39908 26404 40049 26432
rect 39908 26392 39914 26404
rect 40037 26401 40049 26404
rect 40083 26401 40095 26435
rect 40144 26432 40172 26472
rect 40144 26404 41736 26432
rect 40037 26395 40095 26401
rect 31113 26367 31171 26373
rect 31113 26333 31125 26367
rect 31159 26333 31171 26367
rect 31113 26327 31171 26333
rect 34882 26324 34888 26376
rect 34940 26364 34946 26376
rect 36909 26367 36967 26373
rect 36909 26364 36921 26367
rect 34940 26336 36921 26364
rect 34940 26324 34946 26336
rect 36909 26333 36921 26336
rect 36955 26364 36967 26367
rect 37734 26364 37740 26376
rect 36955 26336 37740 26364
rect 36955 26333 36967 26336
rect 36909 26327 36967 26333
rect 37734 26324 37740 26336
rect 37792 26324 37798 26376
rect 39117 26367 39175 26373
rect 39117 26333 39129 26367
rect 39163 26364 39175 26367
rect 39942 26364 39948 26376
rect 39163 26336 39948 26364
rect 39163 26333 39175 26336
rect 39117 26327 39175 26333
rect 39942 26324 39948 26336
rect 40000 26324 40006 26376
rect 41414 26324 41420 26376
rect 41472 26324 41478 26376
rect 41708 26364 41736 26404
rect 48774 26392 48780 26444
rect 48832 26392 48838 26444
rect 42794 26364 42800 26376
rect 41708 26336 42800 26364
rect 42794 26324 42800 26336
rect 42852 26324 42858 26376
rect 43990 26324 43996 26376
rect 44048 26364 44054 26376
rect 47397 26367 47455 26373
rect 47397 26364 47409 26367
rect 44048 26336 47409 26364
rect 44048 26324 44054 26336
rect 47397 26333 47409 26336
rect 47443 26333 47455 26367
rect 47397 26327 47455 26333
rect 48041 26367 48099 26373
rect 48041 26333 48053 26367
rect 48087 26364 48099 26367
rect 48222 26364 48228 26376
rect 48087 26336 48228 26364
rect 48087 26333 48099 26336
rect 48041 26327 48099 26333
rect 48222 26324 48228 26336
rect 48280 26364 48286 26376
rect 48501 26367 48559 26373
rect 48501 26364 48513 26367
rect 48280 26336 48513 26364
rect 48280 26324 48286 26336
rect 48501 26333 48513 26336
rect 48547 26333 48559 26367
rect 48501 26327 48559 26333
rect 23658 26296 23664 26308
rect 23598 26268 23664 26296
rect 23658 26256 23664 26268
rect 23716 26296 23722 26308
rect 23842 26296 23848 26308
rect 23716 26268 23848 26296
rect 23716 26256 23722 26268
rect 23842 26256 23848 26268
rect 23900 26256 23906 26308
rect 24949 26299 25007 26305
rect 24949 26265 24961 26299
rect 24995 26296 25007 26299
rect 32030 26296 32036 26308
rect 24995 26268 32036 26296
rect 24995 26265 25007 26268
rect 24949 26259 25007 26265
rect 32030 26256 32036 26268
rect 32088 26296 32094 26308
rect 32398 26296 32404 26308
rect 32088 26268 32404 26296
rect 32088 26256 32094 26268
rect 32398 26256 32404 26268
rect 32456 26256 32462 26308
rect 32490 26256 32496 26308
rect 32548 26256 32554 26308
rect 32582 26256 32588 26308
rect 32640 26256 32646 26308
rect 33778 26296 33784 26308
rect 33718 26268 33784 26296
rect 33778 26256 33784 26268
rect 33836 26296 33842 26308
rect 33836 26268 34928 26296
rect 33836 26256 33842 26268
rect 24578 26188 24584 26240
rect 24636 26188 24642 26240
rect 26878 26188 26884 26240
rect 26936 26228 26942 26240
rect 27065 26231 27123 26237
rect 27065 26228 27077 26231
rect 26936 26200 27077 26228
rect 26936 26188 26942 26200
rect 27065 26197 27077 26200
rect 27111 26197 27123 26231
rect 27065 26191 27123 26197
rect 27798 26188 27804 26240
rect 27856 26188 27862 26240
rect 32122 26188 32128 26240
rect 32180 26228 32186 26240
rect 32600 26228 32628 26256
rect 34900 26240 34928 26268
rect 34974 26256 34980 26308
rect 35032 26296 35038 26308
rect 35621 26299 35679 26305
rect 35621 26296 35633 26299
rect 35032 26268 35633 26296
rect 35032 26256 35038 26268
rect 35621 26265 35633 26268
rect 35667 26265 35679 26299
rect 35621 26259 35679 26265
rect 37645 26299 37703 26305
rect 37645 26265 37657 26299
rect 37691 26296 37703 26299
rect 38562 26296 38568 26308
rect 37691 26268 38568 26296
rect 37691 26265 37703 26268
rect 37645 26259 37703 26265
rect 38562 26256 38568 26268
rect 38620 26256 38626 26308
rect 39482 26256 39488 26308
rect 39540 26296 39546 26308
rect 40313 26299 40371 26305
rect 40313 26296 40325 26299
rect 39540 26268 40325 26296
rect 39540 26256 39546 26268
rect 40313 26265 40325 26268
rect 40359 26265 40371 26299
rect 40313 26259 40371 26265
rect 32180 26200 32628 26228
rect 32180 26188 32186 26200
rect 34882 26188 34888 26240
rect 34940 26188 34946 26240
rect 47210 26188 47216 26240
rect 47268 26188 47274 26240
rect 1104 26138 49864 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 27950 26138
rect 28002 26086 28014 26138
rect 28066 26086 28078 26138
rect 28130 26086 28142 26138
rect 28194 26086 28206 26138
rect 28258 26086 37950 26138
rect 38002 26086 38014 26138
rect 38066 26086 38078 26138
rect 38130 26086 38142 26138
rect 38194 26086 38206 26138
rect 38258 26086 47950 26138
rect 48002 26086 48014 26138
rect 48066 26086 48078 26138
rect 48130 26086 48142 26138
rect 48194 26086 48206 26138
rect 48258 26086 49864 26138
rect 1104 26064 49864 26086
rect 26970 25984 26976 26036
rect 27028 26024 27034 26036
rect 29086 26024 29092 26036
rect 27028 25996 29092 26024
rect 27028 25984 27034 25996
rect 29086 25984 29092 25996
rect 29144 25984 29150 26036
rect 31481 26027 31539 26033
rect 31481 25993 31493 26027
rect 31527 26024 31539 26027
rect 32309 26027 32367 26033
rect 32309 26024 32321 26027
rect 31527 25996 32321 26024
rect 31527 25993 31539 25996
rect 31481 25987 31539 25993
rect 32309 25993 32321 25996
rect 32355 25993 32367 26027
rect 32309 25987 32367 25993
rect 32674 25984 32680 26036
rect 32732 26024 32738 26036
rect 37829 26027 37887 26033
rect 37829 26024 37841 26027
rect 32732 25996 37841 26024
rect 32732 25984 32738 25996
rect 37829 25993 37841 25996
rect 37875 25993 37887 26027
rect 37829 25987 37887 25993
rect 37921 26027 37979 26033
rect 37921 25993 37933 26027
rect 37967 26024 37979 26027
rect 38654 26024 38660 26036
rect 37967 25996 38660 26024
rect 37967 25993 37979 25996
rect 37921 25987 37979 25993
rect 38654 25984 38660 25996
rect 38712 25984 38718 26036
rect 38838 25984 38844 26036
rect 38896 26024 38902 26036
rect 39025 26027 39083 26033
rect 39025 26024 39037 26027
rect 38896 25996 39037 26024
rect 38896 25984 38902 25996
rect 39025 25993 39037 25996
rect 39071 25993 39083 26027
rect 39025 25987 39083 25993
rect 39117 26027 39175 26033
rect 39117 25993 39129 26027
rect 39163 26024 39175 26027
rect 39298 26024 39304 26036
rect 39163 25996 39304 26024
rect 39163 25993 39175 25996
rect 39117 25987 39175 25993
rect 39298 25984 39304 25996
rect 39356 25984 39362 26036
rect 40770 25984 40776 26036
rect 40828 26024 40834 26036
rect 42061 26027 42119 26033
rect 42061 26024 42073 26027
rect 40828 25996 42073 26024
rect 40828 25984 40834 25996
rect 42061 25993 42073 25996
rect 42107 25993 42119 26027
rect 42061 25987 42119 25993
rect 30282 25956 30288 25968
rect 29946 25928 30288 25956
rect 30282 25916 30288 25928
rect 30340 25916 30346 25968
rect 32766 25916 32772 25968
rect 32824 25916 32830 25968
rect 34698 25916 34704 25968
rect 34756 25956 34762 25968
rect 35345 25959 35403 25965
rect 35345 25956 35357 25959
rect 34756 25928 35357 25956
rect 34756 25916 34762 25928
rect 35345 25925 35357 25928
rect 35391 25956 35403 25959
rect 35802 25956 35808 25968
rect 35391 25928 35808 25956
rect 35391 25925 35403 25928
rect 35345 25919 35403 25925
rect 35802 25916 35808 25928
rect 35860 25916 35866 25968
rect 38562 25916 38568 25968
rect 38620 25956 38626 25968
rect 40589 25959 40647 25965
rect 38620 25928 40356 25956
rect 38620 25916 38626 25928
rect 7466 25848 7472 25900
rect 7524 25888 7530 25900
rect 7561 25891 7619 25897
rect 7561 25888 7573 25891
rect 7524 25860 7573 25888
rect 7524 25848 7530 25860
rect 7561 25857 7573 25860
rect 7607 25857 7619 25891
rect 7561 25851 7619 25857
rect 24121 25891 24179 25897
rect 24121 25857 24133 25891
rect 24167 25888 24179 25891
rect 25133 25891 25191 25897
rect 25133 25888 25145 25891
rect 24167 25860 25145 25888
rect 24167 25857 24179 25860
rect 24121 25851 24179 25857
rect 25133 25857 25145 25860
rect 25179 25857 25191 25891
rect 25133 25851 25191 25857
rect 30558 25848 30564 25900
rect 30616 25888 30622 25900
rect 31389 25891 31447 25897
rect 31389 25888 31401 25891
rect 30616 25860 31401 25888
rect 30616 25848 30622 25860
rect 31389 25857 31401 25860
rect 31435 25857 31447 25891
rect 31389 25851 31447 25857
rect 34514 25848 34520 25900
rect 34572 25888 34578 25900
rect 35253 25891 35311 25897
rect 35253 25888 35265 25891
rect 34572 25860 35265 25888
rect 34572 25848 34578 25860
rect 35253 25857 35265 25860
rect 35299 25857 35311 25891
rect 40126 25888 40132 25900
rect 35253 25851 35311 25857
rect 38120 25860 40132 25888
rect 7745 25823 7803 25829
rect 7745 25789 7757 25823
rect 7791 25820 7803 25823
rect 9030 25820 9036 25832
rect 7791 25792 9036 25820
rect 7791 25789 7803 25792
rect 7745 25783 7803 25789
rect 9030 25780 9036 25792
rect 9088 25780 9094 25832
rect 9398 25780 9404 25832
rect 9456 25780 9462 25832
rect 22370 25780 22376 25832
rect 22428 25820 22434 25832
rect 24213 25823 24271 25829
rect 24213 25820 24225 25823
rect 22428 25792 24225 25820
rect 22428 25780 22434 25792
rect 24213 25789 24225 25792
rect 24259 25789 24271 25823
rect 24213 25783 24271 25789
rect 24397 25823 24455 25829
rect 24397 25789 24409 25823
rect 24443 25820 24455 25823
rect 25222 25820 25228 25832
rect 24443 25792 25228 25820
rect 24443 25789 24455 25792
rect 24397 25783 24455 25789
rect 25222 25780 25228 25792
rect 25280 25780 25286 25832
rect 28442 25780 28448 25832
rect 28500 25780 28506 25832
rect 28721 25823 28779 25829
rect 28721 25820 28733 25823
rect 28552 25792 28733 25820
rect 26234 25712 26240 25764
rect 26292 25752 26298 25764
rect 28552 25752 28580 25792
rect 28721 25789 28733 25792
rect 28767 25820 28779 25823
rect 30098 25820 30104 25832
rect 28767 25792 30104 25820
rect 28767 25789 28779 25792
rect 28721 25783 28779 25789
rect 30098 25780 30104 25792
rect 30156 25780 30162 25832
rect 31665 25823 31723 25829
rect 31665 25789 31677 25823
rect 31711 25820 31723 25823
rect 32490 25820 32496 25832
rect 31711 25792 32496 25820
rect 31711 25789 31723 25792
rect 31665 25783 31723 25789
rect 32490 25780 32496 25792
rect 32548 25780 32554 25832
rect 32953 25823 33011 25829
rect 32953 25789 32965 25823
rect 32999 25820 33011 25823
rect 34698 25820 34704 25832
rect 32999 25792 34704 25820
rect 32999 25789 33011 25792
rect 32953 25783 33011 25789
rect 26292 25724 28580 25752
rect 26292 25712 26298 25724
rect 32214 25712 32220 25764
rect 32272 25752 32278 25764
rect 32968 25752 32996 25783
rect 34698 25780 34704 25792
rect 34756 25780 34762 25832
rect 35529 25823 35587 25829
rect 35529 25789 35541 25823
rect 35575 25820 35587 25823
rect 36078 25820 36084 25832
rect 35575 25792 36084 25820
rect 35575 25789 35587 25792
rect 35529 25783 35587 25789
rect 36078 25780 36084 25792
rect 36136 25780 36142 25832
rect 37458 25780 37464 25832
rect 37516 25820 37522 25832
rect 37642 25820 37648 25832
rect 37516 25792 37648 25820
rect 37516 25780 37522 25792
rect 37642 25780 37648 25792
rect 37700 25780 37706 25832
rect 38120 25829 38148 25860
rect 40126 25848 40132 25860
rect 40184 25848 40190 25900
rect 40328 25897 40356 25928
rect 40589 25925 40601 25959
rect 40635 25956 40647 25959
rect 40678 25956 40684 25968
rect 40635 25928 40684 25956
rect 40635 25925 40647 25928
rect 40589 25919 40647 25925
rect 40678 25916 40684 25928
rect 40736 25916 40742 25968
rect 46106 25916 46112 25968
rect 46164 25916 46170 25968
rect 40313 25891 40371 25897
rect 40313 25857 40325 25891
rect 40359 25857 40371 25891
rect 40313 25851 40371 25857
rect 41598 25848 41604 25900
rect 41656 25888 41662 25900
rect 41656 25874 41722 25888
rect 41656 25860 41736 25874
rect 41656 25848 41662 25860
rect 38105 25823 38163 25829
rect 38105 25789 38117 25823
rect 38151 25789 38163 25823
rect 38105 25783 38163 25789
rect 39206 25780 39212 25832
rect 39264 25780 39270 25832
rect 32272 25724 32996 25752
rect 32272 25712 32278 25724
rect 37826 25712 37832 25764
rect 37884 25752 37890 25764
rect 39666 25752 39672 25764
rect 37884 25724 39672 25752
rect 37884 25712 37890 25724
rect 39666 25712 39672 25724
rect 39724 25712 39730 25764
rect 23753 25687 23811 25693
rect 23753 25653 23765 25687
rect 23799 25684 23811 25687
rect 25774 25684 25780 25696
rect 23799 25656 25780 25684
rect 23799 25653 23811 25656
rect 23753 25647 23811 25653
rect 25774 25644 25780 25656
rect 25832 25644 25838 25696
rect 25866 25644 25872 25696
rect 25924 25684 25930 25696
rect 26053 25687 26111 25693
rect 26053 25684 26065 25687
rect 25924 25656 26065 25684
rect 25924 25644 25930 25656
rect 26053 25653 26065 25656
rect 26099 25653 26111 25687
rect 26053 25647 26111 25653
rect 27430 25644 27436 25696
rect 27488 25684 27494 25696
rect 28534 25684 28540 25696
rect 27488 25656 28540 25684
rect 27488 25644 27494 25656
rect 28534 25644 28540 25656
rect 28592 25644 28598 25696
rect 29914 25644 29920 25696
rect 29972 25684 29978 25696
rect 30193 25687 30251 25693
rect 30193 25684 30205 25687
rect 29972 25656 30205 25684
rect 29972 25644 29978 25656
rect 30193 25653 30205 25656
rect 30239 25653 30251 25687
rect 30193 25647 30251 25653
rect 31018 25644 31024 25696
rect 31076 25644 31082 25696
rect 34885 25687 34943 25693
rect 34885 25653 34897 25687
rect 34931 25684 34943 25687
rect 36814 25684 36820 25696
rect 34931 25656 36820 25684
rect 34931 25653 34943 25656
rect 34885 25647 34943 25653
rect 36814 25644 36820 25656
rect 36872 25644 36878 25696
rect 36906 25644 36912 25696
rect 36964 25644 36970 25696
rect 37458 25644 37464 25696
rect 37516 25644 37522 25696
rect 38654 25644 38660 25696
rect 38712 25644 38718 25696
rect 39574 25644 39580 25696
rect 39632 25684 39638 25696
rect 41708 25684 41736 25860
rect 41966 25848 41972 25900
rect 42024 25888 42030 25900
rect 46845 25891 46903 25897
rect 46845 25888 46857 25891
rect 42024 25860 46857 25888
rect 42024 25848 42030 25860
rect 46845 25857 46857 25860
rect 46891 25857 46903 25891
rect 46845 25851 46903 25857
rect 49326 25848 49332 25900
rect 49384 25848 49390 25900
rect 46290 25712 46296 25764
rect 46348 25712 46354 25764
rect 47026 25712 47032 25764
rect 47084 25712 47090 25764
rect 39632 25656 41736 25684
rect 39632 25644 39638 25656
rect 49142 25644 49148 25696
rect 49200 25644 49206 25696
rect 1104 25594 49864 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 32950 25594
rect 33002 25542 33014 25594
rect 33066 25542 33078 25594
rect 33130 25542 33142 25594
rect 33194 25542 33206 25594
rect 33258 25542 42950 25594
rect 43002 25542 43014 25594
rect 43066 25542 43078 25594
rect 43130 25542 43142 25594
rect 43194 25542 43206 25594
rect 43258 25542 49864 25594
rect 1104 25520 49864 25542
rect 4982 25440 4988 25492
rect 5040 25440 5046 25492
rect 10781 25483 10839 25489
rect 10781 25449 10793 25483
rect 10827 25449 10839 25483
rect 10781 25443 10839 25449
rect 1302 25304 1308 25356
rect 1360 25344 1366 25356
rect 2041 25347 2099 25353
rect 2041 25344 2053 25347
rect 1360 25316 2053 25344
rect 1360 25304 1366 25316
rect 2041 25313 2053 25316
rect 2087 25313 2099 25347
rect 10796 25344 10824 25443
rect 10962 25440 10968 25492
rect 11020 25480 11026 25492
rect 11057 25483 11115 25489
rect 11057 25480 11069 25483
rect 11020 25452 11069 25480
rect 11020 25440 11026 25452
rect 11057 25449 11069 25452
rect 11103 25449 11115 25483
rect 11057 25443 11115 25449
rect 25222 25440 25228 25492
rect 25280 25480 25286 25492
rect 27709 25483 27767 25489
rect 27709 25480 27721 25483
rect 25280 25452 27721 25480
rect 25280 25440 25286 25452
rect 27709 25449 27721 25452
rect 27755 25480 27767 25483
rect 30006 25480 30012 25492
rect 27755 25452 30012 25480
rect 27755 25449 27767 25452
rect 27709 25443 27767 25449
rect 30006 25440 30012 25452
rect 30064 25440 30070 25492
rect 37550 25440 37556 25492
rect 37608 25480 37614 25492
rect 37608 25452 39436 25480
rect 37608 25440 37614 25452
rect 10870 25372 10876 25424
rect 10928 25412 10934 25424
rect 14277 25415 14335 25421
rect 14277 25412 14289 25415
rect 10928 25384 14289 25412
rect 10928 25372 10934 25384
rect 14277 25381 14289 25384
rect 14323 25381 14335 25415
rect 14277 25375 14335 25381
rect 27246 25372 27252 25424
rect 27304 25412 27310 25424
rect 36170 25412 36176 25424
rect 27304 25384 28948 25412
rect 27304 25372 27310 25384
rect 11054 25344 11060 25356
rect 10796 25316 11060 25344
rect 2041 25307 2099 25313
rect 11054 25304 11060 25316
rect 11112 25304 11118 25356
rect 22925 25347 22983 25353
rect 22925 25313 22937 25347
rect 22971 25344 22983 25347
rect 24210 25344 24216 25356
rect 22971 25316 24216 25344
rect 22971 25313 22983 25316
rect 22925 25307 22983 25313
rect 24210 25304 24216 25316
rect 24268 25304 24274 25356
rect 25130 25304 25136 25356
rect 25188 25304 25194 25356
rect 25774 25304 25780 25356
rect 25832 25344 25838 25356
rect 28920 25353 28948 25384
rect 34900 25384 36176 25412
rect 28905 25347 28963 25353
rect 25832 25316 28764 25344
rect 25832 25304 25838 25316
rect 1765 25279 1823 25285
rect 1765 25245 1777 25279
rect 1811 25276 1823 25279
rect 4154 25276 4160 25288
rect 1811 25248 4160 25276
rect 1811 25245 1823 25248
rect 1765 25239 1823 25245
rect 4154 25236 4160 25248
rect 4212 25236 4218 25288
rect 5169 25279 5227 25285
rect 5169 25245 5181 25279
rect 5215 25276 5227 25279
rect 5994 25276 6000 25288
rect 5215 25248 6000 25276
rect 5215 25245 5227 25248
rect 5169 25239 5227 25245
rect 5994 25236 6000 25248
rect 6052 25236 6058 25288
rect 10594 25236 10600 25288
rect 10652 25236 10658 25288
rect 14461 25279 14519 25285
rect 14461 25245 14473 25279
rect 14507 25276 14519 25279
rect 16482 25276 16488 25288
rect 14507 25248 16488 25276
rect 14507 25245 14519 25248
rect 14461 25239 14519 25245
rect 16482 25236 16488 25248
rect 16540 25236 16546 25288
rect 24029 25279 24087 25285
rect 24029 25245 24041 25279
rect 24075 25276 24087 25279
rect 24949 25279 25007 25285
rect 24949 25276 24961 25279
rect 24075 25248 24961 25276
rect 24075 25245 24087 25248
rect 24029 25239 24087 25245
rect 24949 25245 24961 25248
rect 24995 25245 25007 25279
rect 24949 25239 25007 25245
rect 25958 25236 25964 25288
rect 26016 25236 26022 25288
rect 28736 25285 28764 25316
rect 28905 25313 28917 25347
rect 28951 25313 28963 25347
rect 28905 25307 28963 25313
rect 30006 25304 30012 25356
rect 30064 25344 30070 25356
rect 31389 25347 31447 25353
rect 31389 25344 31401 25347
rect 30064 25316 31401 25344
rect 30064 25304 30070 25316
rect 31389 25313 31401 25316
rect 31435 25313 31447 25347
rect 31389 25307 31447 25313
rect 31754 25304 31760 25356
rect 31812 25344 31818 25356
rect 32493 25347 32551 25353
rect 32493 25344 32505 25347
rect 31812 25316 32505 25344
rect 31812 25304 31818 25316
rect 32493 25313 32505 25316
rect 32539 25313 32551 25347
rect 32493 25307 32551 25313
rect 32582 25304 32588 25356
rect 32640 25304 32646 25356
rect 33962 25304 33968 25356
rect 34020 25304 34026 25356
rect 34054 25304 34060 25356
rect 34112 25304 34118 25356
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25245 28779 25279
rect 28721 25239 28779 25245
rect 28813 25279 28871 25285
rect 28813 25245 28825 25279
rect 28859 25276 28871 25279
rect 28994 25276 29000 25288
rect 28859 25248 29000 25276
rect 28859 25245 28871 25248
rect 28813 25239 28871 25245
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 29086 25236 29092 25288
rect 29144 25276 29150 25288
rect 29917 25279 29975 25285
rect 29917 25276 29929 25279
rect 29144 25248 29929 25276
rect 29144 25236 29150 25248
rect 29917 25245 29929 25248
rect 29963 25245 29975 25279
rect 29917 25239 29975 25245
rect 31297 25279 31355 25285
rect 31297 25245 31309 25279
rect 31343 25276 31355 25279
rect 31938 25276 31944 25288
rect 31343 25248 31944 25276
rect 31343 25245 31355 25248
rect 31297 25239 31355 25245
rect 31938 25236 31944 25248
rect 31996 25236 32002 25288
rect 32401 25279 32459 25285
rect 32401 25245 32413 25279
rect 32447 25276 32459 25279
rect 34606 25276 34612 25288
rect 32447 25248 34612 25276
rect 32447 25245 32459 25248
rect 32401 25239 32459 25245
rect 34606 25236 34612 25248
rect 34664 25236 34670 25288
rect 22741 25211 22799 25217
rect 22741 25177 22753 25211
rect 22787 25208 22799 25211
rect 25498 25208 25504 25220
rect 22787 25180 25504 25208
rect 22787 25177 22799 25180
rect 22741 25171 22799 25177
rect 25498 25168 25504 25180
rect 25556 25208 25562 25220
rect 25682 25208 25688 25220
rect 25556 25180 25688 25208
rect 25556 25168 25562 25180
rect 25682 25168 25688 25180
rect 25740 25168 25746 25220
rect 26237 25211 26295 25217
rect 26237 25177 26249 25211
rect 26283 25177 26295 25211
rect 26237 25171 26295 25177
rect 22278 25100 22284 25152
rect 22336 25100 22342 25152
rect 22646 25100 22652 25152
rect 22704 25100 22710 25152
rect 23290 25100 23296 25152
rect 23348 25140 23354 25152
rect 24581 25143 24639 25149
rect 24581 25140 24593 25143
rect 23348 25112 24593 25140
rect 23348 25100 23354 25112
rect 24581 25109 24593 25112
rect 24627 25109 24639 25143
rect 24581 25103 24639 25109
rect 25041 25143 25099 25149
rect 25041 25109 25053 25143
rect 25087 25140 25099 25143
rect 26142 25140 26148 25152
rect 25087 25112 26148 25140
rect 25087 25109 25099 25112
rect 25041 25103 25099 25109
rect 26142 25100 26148 25112
rect 26200 25100 26206 25152
rect 26252 25140 26280 25171
rect 26326 25168 26332 25220
rect 26384 25208 26390 25220
rect 26384 25180 26726 25208
rect 26384 25168 26390 25180
rect 29178 25168 29184 25220
rect 29236 25208 29242 25220
rect 31205 25211 31263 25217
rect 31205 25208 31217 25211
rect 29236 25180 31217 25208
rect 29236 25168 29242 25180
rect 31205 25177 31217 25180
rect 31251 25177 31263 25211
rect 31205 25171 31263 25177
rect 33873 25211 33931 25217
rect 33873 25177 33885 25211
rect 33919 25208 33931 25211
rect 34900 25208 34928 25384
rect 36170 25372 36176 25384
rect 36228 25372 36234 25424
rect 39408 25412 39436 25452
rect 39482 25440 39488 25492
rect 39540 25440 39546 25492
rect 39666 25440 39672 25492
rect 39724 25480 39730 25492
rect 49142 25480 49148 25492
rect 39724 25452 49148 25480
rect 39724 25440 39730 25452
rect 49142 25440 49148 25452
rect 49200 25440 49206 25492
rect 39408 25384 41414 25412
rect 35618 25304 35624 25356
rect 35676 25344 35682 25356
rect 35713 25347 35771 25353
rect 35713 25344 35725 25347
rect 35676 25316 35725 25344
rect 35676 25304 35682 25316
rect 35713 25313 35725 25316
rect 35759 25313 35771 25347
rect 35713 25307 35771 25313
rect 36814 25304 36820 25356
rect 36872 25344 36878 25356
rect 37001 25347 37059 25353
rect 37001 25344 37013 25347
rect 36872 25316 37013 25344
rect 36872 25304 36878 25316
rect 37001 25313 37013 25316
rect 37047 25313 37059 25347
rect 37001 25307 37059 25313
rect 37185 25347 37243 25353
rect 37185 25313 37197 25347
rect 37231 25344 37243 25347
rect 37366 25344 37372 25356
rect 37231 25316 37372 25344
rect 37231 25313 37243 25316
rect 37185 25307 37243 25313
rect 37366 25304 37372 25316
rect 37424 25304 37430 25356
rect 37458 25304 37464 25356
rect 37516 25344 37522 25356
rect 40497 25347 40555 25353
rect 40497 25344 40509 25347
rect 37516 25316 40509 25344
rect 37516 25304 37522 25316
rect 40497 25313 40509 25316
rect 40543 25313 40555 25347
rect 40497 25307 40555 25313
rect 40678 25304 40684 25356
rect 40736 25304 40742 25356
rect 34974 25236 34980 25288
rect 35032 25276 35038 25288
rect 37737 25279 37795 25285
rect 37737 25276 37749 25279
rect 35032 25248 37749 25276
rect 35032 25236 35038 25248
rect 37737 25245 37749 25248
rect 37783 25245 37795 25279
rect 37737 25239 37795 25245
rect 33919 25180 34928 25208
rect 33919 25177 33931 25180
rect 33873 25171 33931 25177
rect 35066 25168 35072 25220
rect 35124 25208 35130 25220
rect 35621 25211 35679 25217
rect 35621 25208 35633 25211
rect 35124 25180 35633 25208
rect 35124 25168 35130 25180
rect 35621 25177 35633 25180
rect 35667 25177 35679 25211
rect 35621 25171 35679 25177
rect 36464 25180 36860 25208
rect 27614 25140 27620 25152
rect 26252 25112 27620 25140
rect 27614 25100 27620 25112
rect 27672 25100 27678 25152
rect 28353 25143 28411 25149
rect 28353 25109 28365 25143
rect 28399 25140 28411 25143
rect 30650 25140 30656 25152
rect 28399 25112 30656 25140
rect 28399 25109 28411 25112
rect 28353 25103 28411 25109
rect 30650 25100 30656 25112
rect 30708 25100 30714 25152
rect 30837 25143 30895 25149
rect 30837 25109 30849 25143
rect 30883 25140 30895 25143
rect 31110 25140 31116 25152
rect 30883 25112 31116 25140
rect 30883 25109 30895 25112
rect 30837 25103 30895 25109
rect 31110 25100 31116 25112
rect 31168 25100 31174 25152
rect 31386 25100 31392 25152
rect 31444 25140 31450 25152
rect 32033 25143 32091 25149
rect 32033 25140 32045 25143
rect 31444 25112 32045 25140
rect 31444 25100 31450 25112
rect 32033 25109 32045 25112
rect 32079 25109 32091 25143
rect 32033 25103 32091 25109
rect 32766 25100 32772 25152
rect 32824 25140 32830 25152
rect 33505 25143 33563 25149
rect 33505 25140 33517 25143
rect 32824 25112 33517 25140
rect 32824 25100 32830 25112
rect 33505 25109 33517 25112
rect 33551 25109 33563 25143
rect 33505 25103 33563 25109
rect 34146 25100 34152 25152
rect 34204 25140 34210 25152
rect 35161 25143 35219 25149
rect 35161 25140 35173 25143
rect 34204 25112 35173 25140
rect 34204 25100 34210 25112
rect 35161 25109 35173 25112
rect 35207 25109 35219 25143
rect 35161 25103 35219 25109
rect 35529 25143 35587 25149
rect 35529 25109 35541 25143
rect 35575 25140 35587 25143
rect 36464 25140 36492 25180
rect 35575 25112 36492 25140
rect 35575 25109 35587 25112
rect 35529 25103 35587 25109
rect 36538 25100 36544 25152
rect 36596 25100 36602 25152
rect 36832 25140 36860 25180
rect 36906 25168 36912 25220
rect 36964 25168 36970 25220
rect 37366 25168 37372 25220
rect 37424 25208 37430 25220
rect 38013 25211 38071 25217
rect 38013 25208 38025 25211
rect 37424 25180 38025 25208
rect 37424 25168 37430 25180
rect 38013 25177 38025 25180
rect 38059 25208 38071 25211
rect 38286 25208 38292 25220
rect 38059 25180 38292 25208
rect 38059 25177 38071 25180
rect 38013 25171 38071 25177
rect 38286 25168 38292 25180
rect 38344 25168 38350 25220
rect 39574 25208 39580 25220
rect 39238 25180 39580 25208
rect 39574 25168 39580 25180
rect 39632 25168 39638 25220
rect 41386 25208 41414 25384
rect 45278 25236 45284 25288
rect 45336 25236 45342 25288
rect 46014 25236 46020 25288
rect 46072 25236 46078 25288
rect 44453 25211 44511 25217
rect 44453 25208 44465 25211
rect 41386 25180 44465 25208
rect 44453 25177 44465 25180
rect 44499 25177 44511 25211
rect 44453 25171 44511 25177
rect 44634 25168 44640 25220
rect 44692 25168 44698 25220
rect 45462 25168 45468 25220
rect 45520 25168 45526 25220
rect 46201 25211 46259 25217
rect 46201 25177 46213 25211
rect 46247 25208 46259 25211
rect 47854 25208 47860 25220
rect 46247 25180 47860 25208
rect 46247 25177 46259 25180
rect 46201 25171 46259 25177
rect 47854 25168 47860 25180
rect 47912 25168 47918 25220
rect 38746 25140 38752 25152
rect 36832 25112 38752 25140
rect 38746 25100 38752 25112
rect 38804 25100 38810 25152
rect 40034 25100 40040 25152
rect 40092 25100 40098 25152
rect 40402 25100 40408 25152
rect 40460 25100 40466 25152
rect 1104 25050 49864 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 27950 25050
rect 28002 24998 28014 25050
rect 28066 24998 28078 25050
rect 28130 24998 28142 25050
rect 28194 24998 28206 25050
rect 28258 24998 37950 25050
rect 38002 24998 38014 25050
rect 38066 24998 38078 25050
rect 38130 24998 38142 25050
rect 38194 24998 38206 25050
rect 38258 24998 47950 25050
rect 48002 24998 48014 25050
rect 48066 24998 48078 25050
rect 48130 24998 48142 25050
rect 48194 24998 48206 25050
rect 48258 24998 49864 25050
rect 1104 24976 49864 24998
rect 9398 24896 9404 24948
rect 9456 24936 9462 24948
rect 27430 24936 27436 24948
rect 9456 24908 27436 24936
rect 9456 24896 9462 24908
rect 27430 24896 27436 24908
rect 27488 24896 27494 24948
rect 28442 24936 28448 24948
rect 27724 24908 28448 24936
rect 21358 24868 21364 24880
rect 21206 24840 21364 24868
rect 21358 24828 21364 24840
rect 21416 24868 21422 24880
rect 23658 24868 23664 24880
rect 21416 24840 23664 24868
rect 21416 24828 21422 24840
rect 23658 24828 23664 24840
rect 23716 24828 23722 24880
rect 25866 24828 25872 24880
rect 25924 24828 25930 24880
rect 25958 24828 25964 24880
rect 26016 24828 26022 24880
rect 26142 24828 26148 24880
rect 26200 24868 26206 24880
rect 26970 24868 26976 24880
rect 26200 24840 26976 24868
rect 26200 24828 26206 24840
rect 26970 24828 26976 24840
rect 27028 24828 27034 24880
rect 27724 24868 27752 24908
rect 28442 24896 28448 24908
rect 28500 24936 28506 24948
rect 28500 24908 28764 24936
rect 28500 24896 28506 24908
rect 27172 24840 27752 24868
rect 8440 24803 8498 24809
rect 8440 24769 8452 24803
rect 8486 24800 8498 24803
rect 9306 24800 9312 24812
rect 8486 24772 9312 24800
rect 8486 24769 8498 24772
rect 8440 24763 8498 24769
rect 9306 24760 9312 24772
rect 9364 24760 9370 24812
rect 22646 24760 22652 24812
rect 22704 24800 22710 24812
rect 22925 24803 22983 24809
rect 22925 24800 22937 24803
rect 22704 24772 22937 24800
rect 22704 24760 22710 24772
rect 22925 24769 22937 24772
rect 22971 24769 22983 24803
rect 25976 24800 26004 24828
rect 27172 24809 27200 24840
rect 27890 24828 27896 24880
rect 27948 24828 27954 24880
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 25976 24772 27169 24800
rect 22925 24763 22983 24769
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 28736 24800 28764 24908
rect 30282 24896 30288 24948
rect 30340 24936 30346 24948
rect 30340 24908 30972 24936
rect 30340 24896 30346 24908
rect 29641 24871 29699 24877
rect 29641 24837 29653 24871
rect 29687 24868 29699 24871
rect 29914 24868 29920 24880
rect 29687 24840 29920 24868
rect 29687 24837 29699 24840
rect 29641 24831 29699 24837
rect 29914 24828 29920 24840
rect 29972 24828 29978 24880
rect 30944 24868 30972 24908
rect 31018 24896 31024 24948
rect 31076 24936 31082 24948
rect 32861 24939 32919 24945
rect 32861 24936 32873 24939
rect 31076 24908 32873 24936
rect 31076 24896 31082 24908
rect 32861 24905 32873 24908
rect 32907 24905 32919 24939
rect 32861 24899 32919 24905
rect 36538 24896 36544 24948
rect 36596 24936 36602 24948
rect 37829 24939 37887 24945
rect 37829 24936 37841 24939
rect 36596 24908 37841 24936
rect 36596 24896 36602 24908
rect 37829 24905 37841 24908
rect 37875 24905 37887 24939
rect 37829 24899 37887 24905
rect 31662 24868 31668 24880
rect 30866 24840 31668 24868
rect 31662 24828 31668 24840
rect 31720 24828 31726 24880
rect 34882 24828 34888 24880
rect 34940 24828 34946 24880
rect 36170 24828 36176 24880
rect 36228 24868 36234 24880
rect 36722 24868 36728 24880
rect 36228 24840 36728 24868
rect 36228 24828 36234 24840
rect 36722 24828 36728 24840
rect 36780 24828 36786 24880
rect 29365 24803 29423 24809
rect 29365 24800 29377 24803
rect 28736 24772 29377 24800
rect 27157 24763 27215 24769
rect 29365 24769 29377 24772
rect 29411 24769 29423 24803
rect 29365 24763 29423 24769
rect 32858 24760 32864 24812
rect 32916 24800 32922 24812
rect 32953 24803 33011 24809
rect 32953 24800 32965 24803
rect 32916 24772 32965 24800
rect 32916 24760 32922 24772
rect 32953 24769 32965 24772
rect 32999 24769 33011 24803
rect 33686 24800 33692 24812
rect 32953 24763 33011 24769
rect 33060 24772 33692 24800
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 8527 24735 8585 24741
rect 8527 24732 8539 24735
rect 8352 24704 8539 24732
rect 8352 24692 8358 24704
rect 8527 24701 8539 24704
rect 8573 24701 8585 24735
rect 8527 24695 8585 24701
rect 19702 24692 19708 24744
rect 19760 24692 19766 24744
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 21266 24732 21272 24744
rect 20027 24704 21272 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 21266 24692 21272 24704
rect 21324 24692 21330 24744
rect 25590 24692 25596 24744
rect 25648 24732 25654 24744
rect 25958 24732 25964 24744
rect 25648 24704 25964 24732
rect 25648 24692 25654 24704
rect 25958 24692 25964 24704
rect 26016 24692 26022 24744
rect 26145 24735 26203 24741
rect 26145 24701 26157 24735
rect 26191 24732 26203 24735
rect 26234 24732 26240 24744
rect 26191 24704 26240 24732
rect 26191 24701 26203 24704
rect 26145 24695 26203 24701
rect 26234 24692 26240 24704
rect 26292 24692 26298 24744
rect 29178 24732 29184 24744
rect 27264 24704 29184 24732
rect 21082 24624 21088 24676
rect 21140 24664 21146 24676
rect 25130 24664 25136 24676
rect 21140 24636 25136 24664
rect 21140 24624 21146 24636
rect 25130 24624 25136 24636
rect 25188 24624 25194 24676
rect 25501 24667 25559 24673
rect 25501 24633 25513 24667
rect 25547 24664 25559 24667
rect 27264 24664 27292 24704
rect 29178 24692 29184 24704
rect 29236 24692 29242 24744
rect 31113 24735 31171 24741
rect 31113 24701 31125 24735
rect 31159 24732 31171 24735
rect 31294 24732 31300 24744
rect 31159 24704 31300 24732
rect 31159 24701 31171 24704
rect 31113 24695 31171 24701
rect 31294 24692 31300 24704
rect 31352 24692 31358 24744
rect 32674 24692 32680 24744
rect 32732 24732 32738 24744
rect 33060 24732 33088 24772
rect 33686 24760 33692 24772
rect 33744 24760 33750 24812
rect 36630 24760 36636 24812
rect 36688 24800 36694 24812
rect 36909 24803 36967 24809
rect 36909 24800 36921 24803
rect 36688 24772 36921 24800
rect 36688 24760 36694 24772
rect 36909 24769 36921 24772
rect 36955 24769 36967 24803
rect 36909 24763 36967 24769
rect 37274 24760 37280 24812
rect 37332 24800 37338 24812
rect 37921 24803 37979 24809
rect 37921 24800 37933 24803
rect 37332 24772 37933 24800
rect 37332 24760 37338 24772
rect 37921 24769 37933 24772
rect 37967 24769 37979 24803
rect 37921 24763 37979 24769
rect 40221 24803 40279 24809
rect 40221 24769 40233 24803
rect 40267 24800 40279 24803
rect 40402 24800 40408 24812
rect 40267 24772 40408 24800
rect 40267 24769 40279 24772
rect 40221 24763 40279 24769
rect 40402 24760 40408 24772
rect 40460 24760 40466 24812
rect 47210 24760 47216 24812
rect 47268 24800 47274 24812
rect 47949 24803 48007 24809
rect 47949 24800 47961 24803
rect 47268 24772 47961 24800
rect 47268 24760 47274 24772
rect 47949 24769 47961 24772
rect 47995 24769 48007 24803
rect 47949 24763 48007 24769
rect 32732 24704 33088 24732
rect 33137 24735 33195 24741
rect 32732 24692 32738 24704
rect 33137 24701 33149 24735
rect 33183 24732 33195 24735
rect 33870 24732 33876 24744
rect 33183 24704 33876 24732
rect 33183 24701 33195 24704
rect 33137 24695 33195 24701
rect 33870 24692 33876 24704
rect 33928 24692 33934 24744
rect 33965 24735 34023 24741
rect 33965 24701 33977 24735
rect 34011 24701 34023 24735
rect 33965 24695 34023 24701
rect 25547 24636 27292 24664
rect 25547 24633 25559 24636
rect 25501 24627 25559 24633
rect 32306 24624 32312 24676
rect 32364 24664 32370 24676
rect 33980 24664 34008 24695
rect 34238 24692 34244 24744
rect 34296 24692 34302 24744
rect 34698 24692 34704 24744
rect 34756 24732 34762 24744
rect 35989 24735 36047 24741
rect 35989 24732 36001 24735
rect 34756 24704 36001 24732
rect 34756 24692 34762 24704
rect 35989 24701 36001 24704
rect 36035 24701 36047 24735
rect 35989 24695 36047 24701
rect 38105 24735 38163 24741
rect 38105 24701 38117 24735
rect 38151 24732 38163 24735
rect 39482 24732 39488 24744
rect 38151 24704 39488 24732
rect 38151 24701 38163 24704
rect 38105 24695 38163 24701
rect 39482 24692 39488 24704
rect 39540 24692 39546 24744
rect 49142 24692 49148 24744
rect 49200 24692 49206 24744
rect 32364 24636 34008 24664
rect 32364 24624 32370 24636
rect 21453 24599 21511 24605
rect 21453 24565 21465 24599
rect 21499 24596 21511 24599
rect 21542 24596 21548 24608
rect 21499 24568 21548 24596
rect 21499 24565 21511 24568
rect 21453 24559 21511 24565
rect 21542 24556 21548 24568
rect 21600 24556 21606 24608
rect 27420 24599 27478 24605
rect 27420 24565 27432 24599
rect 27466 24596 27478 24599
rect 27522 24596 27528 24608
rect 27466 24568 27528 24596
rect 27466 24565 27478 24568
rect 27420 24559 27478 24565
rect 27522 24556 27528 24568
rect 27580 24556 27586 24608
rect 27614 24556 27620 24608
rect 27672 24596 27678 24608
rect 28905 24599 28963 24605
rect 28905 24596 28917 24599
rect 27672 24568 28917 24596
rect 27672 24556 27678 24568
rect 28905 24565 28917 24568
rect 28951 24596 28963 24599
rect 30282 24596 30288 24608
rect 28951 24568 30288 24596
rect 28951 24565 28963 24568
rect 28905 24559 28963 24565
rect 30282 24556 30288 24568
rect 30340 24556 30346 24608
rect 31202 24556 31208 24608
rect 31260 24596 31266 24608
rect 32214 24596 32220 24608
rect 31260 24568 32220 24596
rect 31260 24556 31266 24568
rect 32214 24556 32220 24568
rect 32272 24556 32278 24608
rect 32398 24556 32404 24608
rect 32456 24596 32462 24608
rect 32493 24599 32551 24605
rect 32493 24596 32505 24599
rect 32456 24568 32505 24596
rect 32456 24556 32462 24568
rect 32493 24565 32505 24568
rect 32539 24565 32551 24599
rect 33980 24596 34008 24636
rect 36725 24667 36783 24673
rect 36725 24633 36737 24667
rect 36771 24664 36783 24667
rect 36771 24636 41414 24664
rect 36771 24633 36783 24636
rect 36725 24627 36783 24633
rect 34974 24596 34980 24608
rect 33980 24568 34980 24596
rect 32493 24559 32551 24565
rect 34974 24556 34980 24568
rect 35032 24556 35038 24608
rect 35434 24556 35440 24608
rect 35492 24596 35498 24608
rect 37461 24599 37519 24605
rect 37461 24596 37473 24599
rect 35492 24568 37473 24596
rect 35492 24556 35498 24568
rect 37461 24565 37473 24568
rect 37507 24565 37519 24599
rect 41386 24596 41414 24636
rect 43806 24596 43812 24608
rect 41386 24568 43812 24596
rect 37461 24559 37519 24565
rect 43806 24556 43812 24568
rect 43864 24556 43870 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 10965 24395 11023 24401
rect 10965 24361 10977 24395
rect 11011 24392 11023 24395
rect 14090 24392 14096 24404
rect 11011 24364 14096 24392
rect 11011 24361 11023 24364
rect 10965 24355 11023 24361
rect 14090 24352 14096 24364
rect 14148 24352 14154 24404
rect 21818 24352 21824 24404
rect 21876 24392 21882 24404
rect 21876 24364 26740 24392
rect 21876 24352 21882 24364
rect 19702 24216 19708 24268
rect 19760 24256 19766 24268
rect 20809 24259 20867 24265
rect 20809 24256 20821 24259
rect 19760 24228 20821 24256
rect 19760 24216 19766 24228
rect 20809 24225 20821 24228
rect 20855 24256 20867 24259
rect 21450 24256 21456 24268
rect 20855 24228 21456 24256
rect 20855 24225 20867 24228
rect 20809 24219 20867 24225
rect 21450 24216 21456 24228
rect 21508 24216 21514 24268
rect 25498 24216 25504 24268
rect 25556 24216 25562 24268
rect 26712 24265 26740 24364
rect 26786 24352 26792 24404
rect 26844 24392 26850 24404
rect 34422 24392 34428 24404
rect 26844 24364 34428 24392
rect 26844 24352 26850 24364
rect 34422 24352 34428 24364
rect 34480 24392 34486 24404
rect 34606 24392 34612 24404
rect 34480 24364 34612 24392
rect 34480 24352 34486 24364
rect 34606 24352 34612 24364
rect 34664 24352 34670 24404
rect 27430 24284 27436 24336
rect 27488 24324 27494 24336
rect 31202 24324 31208 24336
rect 27488 24296 28120 24324
rect 27488 24284 27494 24296
rect 28092 24268 28120 24296
rect 28276 24296 31208 24324
rect 25593 24259 25651 24265
rect 25593 24225 25605 24259
rect 25639 24225 25651 24259
rect 25593 24219 25651 24225
rect 26697 24259 26755 24265
rect 26697 24225 26709 24259
rect 26743 24225 26755 24259
rect 26697 24219 26755 24225
rect 26881 24259 26939 24265
rect 26881 24225 26893 24259
rect 26927 24256 26939 24259
rect 27522 24256 27528 24268
rect 26927 24228 27528 24256
rect 26927 24225 26939 24228
rect 26881 24219 26939 24225
rect 10594 24148 10600 24200
rect 10652 24188 10658 24200
rect 10689 24191 10747 24197
rect 10689 24188 10701 24191
rect 10652 24160 10701 24188
rect 10652 24148 10658 24160
rect 10689 24157 10701 24160
rect 10735 24188 10747 24191
rect 12618 24188 12624 24200
rect 10735 24160 12624 24188
rect 10735 24157 10747 24160
rect 10689 24151 10747 24157
rect 12618 24148 12624 24160
rect 12676 24148 12682 24200
rect 22830 24148 22836 24200
rect 22888 24188 22894 24200
rect 25608 24188 25636 24219
rect 27522 24216 27528 24228
rect 27580 24216 27586 24268
rect 28074 24216 28080 24268
rect 28132 24216 28138 24268
rect 28276 24265 28304 24296
rect 31202 24284 31208 24296
rect 31260 24284 31266 24336
rect 39482 24324 39488 24336
rect 34900 24296 35112 24324
rect 28261 24259 28319 24265
rect 28261 24225 28273 24259
rect 28307 24225 28319 24259
rect 28261 24219 28319 24225
rect 30190 24216 30196 24268
rect 30248 24216 30254 24268
rect 30282 24216 30288 24268
rect 30340 24216 30346 24268
rect 32858 24216 32864 24268
rect 32916 24256 32922 24268
rect 34241 24259 34299 24265
rect 34241 24256 34253 24259
rect 32916 24228 34253 24256
rect 32916 24216 32922 24228
rect 34241 24225 34253 24228
rect 34287 24256 34299 24259
rect 34900 24256 34928 24296
rect 34287 24228 34928 24256
rect 34287 24225 34299 24228
rect 34241 24219 34299 24225
rect 34974 24216 34980 24268
rect 35032 24216 35038 24268
rect 35084 24256 35112 24296
rect 37660 24296 39488 24324
rect 35253 24259 35311 24265
rect 35253 24256 35265 24259
rect 35084 24228 35265 24256
rect 35253 24225 35265 24228
rect 35299 24256 35311 24259
rect 35710 24256 35716 24268
rect 35299 24228 35716 24256
rect 35299 24225 35311 24228
rect 35253 24219 35311 24225
rect 35710 24216 35716 24228
rect 35768 24256 35774 24268
rect 37660 24256 37688 24296
rect 39482 24284 39488 24296
rect 39540 24284 39546 24336
rect 35768 24228 37688 24256
rect 35768 24216 35774 24228
rect 37734 24216 37740 24268
rect 37792 24216 37798 24268
rect 40218 24216 40224 24268
rect 40276 24256 40282 24268
rect 40497 24259 40555 24265
rect 40497 24256 40509 24259
rect 40276 24228 40509 24256
rect 40276 24216 40282 24228
rect 40497 24225 40509 24228
rect 40543 24225 40555 24259
rect 40497 24219 40555 24225
rect 40681 24259 40739 24265
rect 40681 24225 40693 24259
rect 40727 24256 40739 24259
rect 40770 24256 40776 24268
rect 40727 24228 40776 24256
rect 40727 24225 40739 24228
rect 40681 24219 40739 24225
rect 40770 24216 40776 24228
rect 40828 24216 40834 24268
rect 30101 24191 30159 24197
rect 30101 24188 30113 24191
rect 22888 24160 25636 24188
rect 26252 24160 30113 24188
rect 22888 24148 22894 24160
rect 21082 24080 21088 24132
rect 21140 24080 21146 24132
rect 23658 24120 23664 24132
rect 22310 24092 23664 24120
rect 23658 24080 23664 24092
rect 23716 24080 23722 24132
rect 11146 24012 11152 24064
rect 11204 24012 11210 24064
rect 21266 24012 21272 24064
rect 21324 24052 21330 24064
rect 22554 24052 22560 24064
rect 21324 24024 22560 24052
rect 21324 24012 21330 24024
rect 22554 24012 22560 24024
rect 22612 24012 22618 24064
rect 23842 24012 23848 24064
rect 23900 24052 23906 24064
rect 25041 24055 25099 24061
rect 25041 24052 25053 24055
rect 23900 24024 25053 24052
rect 23900 24012 23906 24024
rect 25041 24021 25053 24024
rect 25087 24021 25099 24055
rect 25041 24015 25099 24021
rect 25409 24055 25467 24061
rect 25409 24021 25421 24055
rect 25455 24052 25467 24055
rect 26142 24052 26148 24064
rect 25455 24024 26148 24052
rect 25455 24021 25467 24024
rect 25409 24015 25467 24021
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 26252 24061 26280 24160
rect 30101 24157 30113 24160
rect 30147 24157 30159 24191
rect 30101 24151 30159 24157
rect 30466 24148 30472 24200
rect 30524 24188 30530 24200
rect 32674 24188 32680 24200
rect 30524 24160 32680 24188
rect 30524 24148 30530 24160
rect 32674 24148 32680 24160
rect 32732 24148 32738 24200
rect 33410 24148 33416 24200
rect 33468 24188 33474 24200
rect 33965 24191 34023 24197
rect 33965 24188 33977 24191
rect 33468 24160 33977 24188
rect 33468 24148 33474 24160
rect 33965 24157 33977 24160
rect 34011 24188 34023 24191
rect 34422 24188 34428 24200
rect 34011 24160 34428 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 34422 24148 34428 24160
rect 34480 24148 34486 24200
rect 37645 24191 37703 24197
rect 37645 24157 37657 24191
rect 37691 24188 37703 24191
rect 37826 24188 37832 24200
rect 37691 24160 37832 24188
rect 37691 24157 37703 24160
rect 37645 24151 37703 24157
rect 37826 24148 37832 24160
rect 37884 24148 37890 24200
rect 40034 24148 40040 24200
rect 40092 24188 40098 24200
rect 40405 24191 40463 24197
rect 40405 24188 40417 24191
rect 40092 24160 40417 24188
rect 40092 24148 40098 24160
rect 40405 24157 40417 24160
rect 40451 24157 40463 24191
rect 40405 24151 40463 24157
rect 47762 24148 47768 24200
rect 47820 24188 47826 24200
rect 47949 24191 48007 24197
rect 47949 24188 47961 24191
rect 47820 24160 47961 24188
rect 47820 24148 47826 24160
rect 47949 24157 47961 24160
rect 47995 24157 48007 24191
rect 47949 24151 48007 24157
rect 27985 24123 28043 24129
rect 27985 24089 27997 24123
rect 28031 24120 28043 24123
rect 29086 24120 29092 24132
rect 28031 24092 29092 24120
rect 28031 24089 28043 24092
rect 27985 24083 28043 24089
rect 29086 24080 29092 24092
rect 29144 24080 29150 24132
rect 34698 24120 34704 24132
rect 29748 24092 34704 24120
rect 26237 24055 26295 24061
rect 26237 24021 26249 24055
rect 26283 24021 26295 24055
rect 26237 24015 26295 24021
rect 26602 24012 26608 24064
rect 26660 24012 26666 24064
rect 27614 24012 27620 24064
rect 27672 24012 27678 24064
rect 28074 24012 28080 24064
rect 28132 24052 28138 24064
rect 28442 24052 28448 24064
rect 28132 24024 28448 24052
rect 28132 24012 28138 24024
rect 28442 24012 28448 24024
rect 28500 24012 28506 24064
rect 29748 24061 29776 24092
rect 34698 24080 34704 24092
rect 34756 24080 34762 24132
rect 35710 24120 35716 24132
rect 35084 24092 35716 24120
rect 29733 24055 29791 24061
rect 29733 24021 29745 24055
rect 29779 24021 29791 24055
rect 29733 24015 29791 24021
rect 30190 24012 30196 24064
rect 30248 24052 30254 24064
rect 33410 24052 33416 24064
rect 30248 24024 33416 24052
rect 30248 24012 30254 24024
rect 33410 24012 33416 24024
rect 33468 24012 33474 24064
rect 33597 24055 33655 24061
rect 33597 24021 33609 24055
rect 33643 24052 33655 24055
rect 33870 24052 33876 24064
rect 33643 24024 33876 24052
rect 33643 24021 33655 24024
rect 33597 24015 33655 24021
rect 33870 24012 33876 24024
rect 33928 24012 33934 24064
rect 34057 24055 34115 24061
rect 34057 24021 34069 24055
rect 34103 24052 34115 24055
rect 34422 24052 34428 24064
rect 34103 24024 34428 24052
rect 34103 24021 34115 24024
rect 34057 24015 34115 24021
rect 34422 24012 34428 24024
rect 34480 24012 34486 24064
rect 34514 24012 34520 24064
rect 34572 24052 34578 24064
rect 35084 24052 35112 24092
rect 35710 24080 35716 24092
rect 35768 24080 35774 24132
rect 37366 24080 37372 24132
rect 37424 24120 37430 24132
rect 37553 24123 37611 24129
rect 37553 24120 37565 24123
rect 37424 24092 37565 24120
rect 37424 24080 37430 24092
rect 37553 24089 37565 24092
rect 37599 24120 37611 24123
rect 38470 24120 38476 24132
rect 37599 24092 38476 24120
rect 37599 24089 37611 24092
rect 37553 24083 37611 24089
rect 38470 24080 38476 24092
rect 38528 24080 38534 24132
rect 49142 24080 49148 24132
rect 49200 24080 49206 24132
rect 34572 24024 35112 24052
rect 34572 24012 34578 24024
rect 35158 24012 35164 24064
rect 35216 24052 35222 24064
rect 35618 24052 35624 24064
rect 35216 24024 35624 24052
rect 35216 24012 35222 24024
rect 35618 24012 35624 24024
rect 35676 24052 35682 24064
rect 36725 24055 36783 24061
rect 36725 24052 36737 24055
rect 35676 24024 36737 24052
rect 35676 24012 35682 24024
rect 36725 24021 36737 24024
rect 36771 24021 36783 24055
rect 36725 24015 36783 24021
rect 37185 24055 37243 24061
rect 37185 24021 37197 24055
rect 37231 24052 37243 24055
rect 37458 24052 37464 24064
rect 37231 24024 37464 24052
rect 37231 24021 37243 24024
rect 37185 24015 37243 24021
rect 37458 24012 37464 24024
rect 37516 24012 37522 24064
rect 37642 24012 37648 24064
rect 37700 24052 37706 24064
rect 37826 24052 37832 24064
rect 37700 24024 37832 24052
rect 37700 24012 37706 24024
rect 37826 24012 37832 24024
rect 37884 24012 37890 24064
rect 40034 24012 40040 24064
rect 40092 24012 40098 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 5994 23808 6000 23860
rect 6052 23848 6058 23860
rect 9493 23851 9551 23857
rect 9493 23848 9505 23851
rect 6052 23820 9505 23848
rect 6052 23808 6058 23820
rect 9493 23817 9505 23820
rect 9539 23817 9551 23851
rect 9493 23811 9551 23817
rect 11054 23808 11060 23860
rect 11112 23848 11118 23860
rect 16301 23851 16359 23857
rect 16301 23848 16313 23851
rect 11112 23820 16313 23848
rect 11112 23808 11118 23820
rect 12636 23789 12664 23820
rect 16301 23817 16313 23820
rect 16347 23817 16359 23851
rect 16301 23811 16359 23817
rect 16482 23808 16488 23860
rect 16540 23848 16546 23860
rect 19337 23851 19395 23857
rect 19337 23848 19349 23851
rect 16540 23820 19349 23848
rect 16540 23808 16546 23820
rect 19337 23817 19349 23820
rect 19383 23817 19395 23851
rect 19337 23811 19395 23817
rect 19705 23851 19763 23857
rect 19705 23817 19717 23851
rect 19751 23848 19763 23851
rect 20717 23851 20775 23857
rect 20717 23848 20729 23851
rect 19751 23820 20729 23848
rect 19751 23817 19763 23820
rect 19705 23811 19763 23817
rect 20717 23817 20729 23820
rect 20763 23817 20775 23851
rect 20717 23811 20775 23817
rect 21085 23851 21143 23857
rect 21085 23817 21097 23851
rect 21131 23848 21143 23851
rect 23290 23848 23296 23860
rect 21131 23820 23296 23848
rect 21131 23817 21143 23820
rect 21085 23811 21143 23817
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 26237 23851 26295 23857
rect 26237 23817 26249 23851
rect 26283 23848 26295 23851
rect 26786 23848 26792 23860
rect 26283 23820 26792 23848
rect 26283 23817 26295 23820
rect 26237 23811 26295 23817
rect 26786 23808 26792 23820
rect 26844 23808 26850 23860
rect 27801 23851 27859 23857
rect 27801 23817 27813 23851
rect 27847 23848 27859 23851
rect 28629 23851 28687 23857
rect 28629 23848 28641 23851
rect 27847 23820 28641 23848
rect 27847 23817 27859 23820
rect 27801 23811 27859 23817
rect 28629 23817 28641 23820
rect 28675 23848 28687 23851
rect 30466 23848 30472 23860
rect 28675 23820 30472 23848
rect 28675 23817 28687 23820
rect 28629 23811 28687 23817
rect 30466 23808 30472 23820
rect 30524 23808 30530 23860
rect 34054 23808 34060 23860
rect 34112 23808 34118 23860
rect 34422 23808 34428 23860
rect 34480 23848 34486 23860
rect 37090 23848 37096 23860
rect 34480 23820 37096 23848
rect 34480 23808 34486 23820
rect 37090 23808 37096 23820
rect 37148 23808 37154 23860
rect 39390 23808 39396 23860
rect 39448 23848 39454 23860
rect 40497 23851 40555 23857
rect 40497 23848 40509 23851
rect 39448 23820 40509 23848
rect 39448 23808 39454 23820
rect 40497 23817 40509 23820
rect 40543 23817 40555 23851
rect 40497 23811 40555 23817
rect 12621 23783 12679 23789
rect 12621 23749 12633 23783
rect 12667 23749 12679 23783
rect 15286 23780 15292 23792
rect 13846 23752 15292 23780
rect 12621 23743 12679 23749
rect 15286 23740 15292 23752
rect 15344 23740 15350 23792
rect 20990 23740 20996 23792
rect 21048 23780 21054 23792
rect 21818 23780 21824 23792
rect 21048 23752 21824 23780
rect 21048 23740 21054 23752
rect 21818 23740 21824 23752
rect 21876 23740 21882 23792
rect 23658 23780 23664 23792
rect 23506 23752 23664 23780
rect 23658 23740 23664 23752
rect 23716 23740 23722 23792
rect 26602 23780 26608 23792
rect 25424 23752 26608 23780
rect 8849 23715 8907 23721
rect 8849 23681 8861 23715
rect 8895 23712 8907 23715
rect 12158 23712 12164 23724
rect 8895 23684 12164 23712
rect 8895 23681 8907 23684
rect 8849 23675 8907 23681
rect 12158 23672 12164 23684
rect 12216 23672 12222 23724
rect 12345 23715 12403 23721
rect 12345 23681 12357 23715
rect 12391 23681 12403 23715
rect 12345 23675 12403 23681
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 9033 23647 9091 23653
rect 9033 23644 9045 23647
rect 7892 23616 9045 23644
rect 7892 23604 7898 23616
rect 9033 23613 9045 23616
rect 9079 23644 9091 23647
rect 11146 23644 11152 23656
rect 9079 23616 11152 23644
rect 9079 23613 9091 23616
rect 9033 23607 9091 23613
rect 11146 23604 11152 23616
rect 11204 23604 11210 23656
rect 12360 23644 12388 23675
rect 21450 23672 21456 23724
rect 21508 23712 21514 23724
rect 25424 23721 25452 23752
rect 26602 23740 26608 23752
rect 26660 23740 26666 23792
rect 27614 23740 27620 23792
rect 27672 23780 27678 23792
rect 30558 23780 30564 23792
rect 27672 23752 30564 23780
rect 27672 23740 27678 23752
rect 30558 23740 30564 23752
rect 30616 23740 30622 23792
rect 32490 23780 32496 23792
rect 31726 23752 32496 23780
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21508 23684 22017 23712
rect 21508 23672 21514 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 25409 23715 25467 23721
rect 22005 23675 22063 23681
rect 23492 23684 24164 23712
rect 14553 23647 14611 23653
rect 14553 23644 14565 23647
rect 12360 23616 14565 23644
rect 14553 23613 14565 23616
rect 14599 23613 14611 23647
rect 14553 23607 14611 23613
rect 14829 23647 14887 23653
rect 14829 23613 14841 23647
rect 14875 23644 14887 23647
rect 16482 23644 16488 23656
rect 14875 23616 16488 23644
rect 14875 23613 14887 23616
rect 14829 23607 14887 23613
rect 14090 23536 14096 23588
rect 14148 23536 14154 23588
rect 14568 23508 14596 23607
rect 16482 23604 16488 23616
rect 16540 23604 16546 23656
rect 19797 23647 19855 23653
rect 19797 23613 19809 23647
rect 19843 23613 19855 23647
rect 19797 23607 19855 23613
rect 19981 23647 20039 23653
rect 19981 23613 19993 23647
rect 20027 23613 20039 23647
rect 19981 23607 20039 23613
rect 16206 23508 16212 23520
rect 14568 23480 16212 23508
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 19812 23508 19840 23607
rect 19996 23576 20024 23607
rect 20898 23604 20904 23656
rect 20956 23644 20962 23656
rect 21177 23647 21235 23653
rect 21177 23644 21189 23647
rect 20956 23616 21189 23644
rect 20956 23604 20962 23616
rect 21177 23613 21189 23616
rect 21223 23613 21235 23647
rect 21177 23607 21235 23613
rect 21266 23604 21272 23656
rect 21324 23604 21330 23656
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 22066 23616 22293 23644
rect 21542 23576 21548 23588
rect 19996 23548 21548 23576
rect 21542 23536 21548 23548
rect 21600 23576 21606 23588
rect 22066 23576 22094 23616
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 22281 23607 22339 23613
rect 21600 23548 22094 23576
rect 21600 23536 21606 23548
rect 22094 23508 22100 23520
rect 19812 23480 22100 23508
rect 22094 23468 22100 23480
rect 22152 23468 22158 23520
rect 22462 23468 22468 23520
rect 22520 23508 22526 23520
rect 23492 23508 23520 23684
rect 24029 23647 24087 23653
rect 24029 23613 24041 23647
rect 24075 23613 24087 23647
rect 24136 23644 24164 23684
rect 25409 23681 25421 23715
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 26142 23672 26148 23724
rect 26200 23712 26206 23724
rect 31570 23712 31576 23724
rect 26200 23684 31576 23712
rect 26200 23672 26206 23684
rect 31570 23672 31576 23684
rect 31628 23712 31634 23724
rect 31726 23712 31754 23752
rect 32490 23740 32496 23752
rect 32548 23740 32554 23792
rect 33870 23740 33876 23792
rect 33928 23780 33934 23792
rect 34977 23783 35035 23789
rect 34977 23780 34989 23783
rect 33928 23752 34989 23780
rect 33928 23740 33934 23752
rect 34977 23749 34989 23752
rect 35023 23749 35035 23783
rect 34977 23743 35035 23749
rect 37734 23740 37740 23792
rect 37792 23780 37798 23792
rect 39025 23783 39083 23789
rect 39025 23780 39037 23783
rect 37792 23752 39037 23780
rect 37792 23740 37798 23752
rect 39025 23749 39037 23752
rect 39071 23749 39083 23783
rect 39025 23743 39083 23749
rect 39574 23740 39580 23792
rect 39632 23740 39638 23792
rect 31628 23684 31754 23712
rect 31628 23672 31634 23684
rect 32306 23672 32312 23724
rect 32364 23672 32370 23724
rect 33686 23672 33692 23724
rect 33744 23712 33750 23724
rect 34514 23712 34520 23724
rect 33744 23684 34520 23712
rect 33744 23672 33750 23684
rect 34514 23672 34520 23684
rect 34572 23672 34578 23724
rect 34885 23715 34943 23721
rect 34885 23681 34897 23715
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 26329 23647 26387 23653
rect 26329 23644 26341 23647
rect 24136 23616 26341 23644
rect 24029 23607 24087 23613
rect 26329 23613 26341 23616
rect 26375 23613 26387 23647
rect 26329 23607 26387 23613
rect 23658 23536 23664 23588
rect 23716 23576 23722 23588
rect 24044 23576 24072 23607
rect 26418 23604 26424 23656
rect 26476 23604 26482 23656
rect 26510 23604 26516 23656
rect 26568 23644 26574 23656
rect 28721 23647 28779 23653
rect 28721 23644 28733 23647
rect 26568 23616 28733 23644
rect 26568 23604 26574 23616
rect 28721 23613 28733 23616
rect 28767 23613 28779 23647
rect 28721 23607 28779 23613
rect 28813 23647 28871 23653
rect 28813 23613 28825 23647
rect 28859 23613 28871 23647
rect 28813 23607 28871 23613
rect 24670 23576 24676 23588
rect 23716 23548 24676 23576
rect 23716 23536 23722 23548
rect 24670 23536 24676 23548
rect 24728 23576 24734 23588
rect 28828 23576 28856 23607
rect 32674 23604 32680 23656
rect 32732 23644 32738 23656
rect 34900 23644 34928 23675
rect 38562 23672 38568 23724
rect 38620 23712 38626 23724
rect 38749 23715 38807 23721
rect 38749 23712 38761 23715
rect 38620 23684 38761 23712
rect 38620 23672 38626 23684
rect 38749 23681 38761 23684
rect 38795 23681 38807 23715
rect 38749 23675 38807 23681
rect 46750 23672 46756 23724
rect 46808 23712 46814 23724
rect 47949 23715 48007 23721
rect 47949 23712 47961 23715
rect 46808 23684 47961 23712
rect 46808 23672 46814 23684
rect 47949 23681 47961 23684
rect 47995 23681 48007 23715
rect 47949 23675 48007 23681
rect 32732 23616 34928 23644
rect 32732 23604 32738 23616
rect 35158 23604 35164 23656
rect 35216 23604 35222 23656
rect 49142 23604 49148 23656
rect 49200 23604 49206 23656
rect 24728 23548 28856 23576
rect 24728 23536 24734 23548
rect 22520 23480 23520 23508
rect 24765 23511 24823 23517
rect 22520 23468 22526 23480
rect 24765 23477 24777 23511
rect 24811 23508 24823 23511
rect 24946 23508 24952 23520
rect 24811 23480 24952 23508
rect 24811 23477 24823 23480
rect 24765 23471 24823 23477
rect 24946 23468 24952 23480
rect 25004 23468 25010 23520
rect 25866 23468 25872 23520
rect 25924 23468 25930 23520
rect 26142 23468 26148 23520
rect 26200 23508 26206 23520
rect 28261 23511 28319 23517
rect 28261 23508 28273 23511
rect 26200 23480 28273 23508
rect 26200 23468 26206 23480
rect 28261 23477 28273 23480
rect 28307 23477 28319 23511
rect 28261 23471 28319 23477
rect 32572 23511 32630 23517
rect 32572 23477 32584 23511
rect 32618 23508 32630 23511
rect 34330 23508 34336 23520
rect 32618 23480 34336 23508
rect 32618 23477 32630 23480
rect 32572 23471 32630 23477
rect 34330 23468 34336 23480
rect 34388 23468 34394 23520
rect 34514 23468 34520 23520
rect 34572 23468 34578 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 4154 23264 4160 23316
rect 4212 23304 4218 23316
rect 5169 23307 5227 23313
rect 5169 23304 5181 23307
rect 4212 23276 5181 23304
rect 4212 23264 4218 23276
rect 5169 23273 5181 23276
rect 5215 23273 5227 23307
rect 5169 23267 5227 23273
rect 26970 23264 26976 23316
rect 27028 23304 27034 23316
rect 27522 23304 27528 23316
rect 27028 23276 27528 23304
rect 27028 23264 27034 23276
rect 27522 23264 27528 23276
rect 27580 23264 27586 23316
rect 27614 23264 27620 23316
rect 27672 23304 27678 23316
rect 28905 23307 28963 23313
rect 28905 23304 28917 23307
rect 27672 23276 28917 23304
rect 27672 23264 27678 23276
rect 28905 23273 28917 23276
rect 28951 23273 28963 23307
rect 28905 23267 28963 23273
rect 31846 23264 31852 23316
rect 31904 23304 31910 23316
rect 32582 23304 32588 23316
rect 31904 23276 32588 23304
rect 31904 23264 31910 23276
rect 32582 23264 32588 23276
rect 32640 23264 32646 23316
rect 34238 23264 34244 23316
rect 34296 23304 34302 23316
rect 36633 23307 36691 23313
rect 36633 23304 36645 23307
rect 34296 23276 36645 23304
rect 34296 23264 34302 23276
rect 36633 23273 36645 23276
rect 36679 23273 36691 23307
rect 36633 23267 36691 23273
rect 34057 23239 34115 23245
rect 34057 23205 34069 23239
rect 34103 23236 34115 23239
rect 34330 23236 34336 23248
rect 34103 23208 34336 23236
rect 34103 23205 34115 23208
rect 34057 23199 34115 23205
rect 34330 23196 34336 23208
rect 34388 23196 34394 23248
rect 37461 23239 37519 23245
rect 37461 23205 37473 23239
rect 37507 23236 37519 23239
rect 44082 23236 44088 23248
rect 37507 23208 44088 23236
rect 37507 23205 37519 23208
rect 37461 23199 37519 23205
rect 44082 23196 44088 23208
rect 44140 23196 44146 23248
rect 1302 23128 1308 23180
rect 1360 23168 1366 23180
rect 2041 23171 2099 23177
rect 2041 23168 2053 23171
rect 1360 23140 2053 23168
rect 1360 23128 1366 23140
rect 2041 23137 2053 23140
rect 2087 23137 2099 23171
rect 5534 23168 5540 23180
rect 2041 23131 2099 23137
rect 3528 23140 5540 23168
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 3528 23100 3556 23140
rect 5534 23128 5540 23140
rect 5592 23128 5598 23180
rect 9030 23128 9036 23180
rect 9088 23168 9094 23180
rect 9263 23171 9321 23177
rect 9263 23168 9275 23171
rect 9088 23140 9275 23168
rect 9088 23128 9094 23140
rect 9263 23137 9275 23140
rect 9309 23137 9321 23171
rect 9263 23131 9321 23137
rect 16206 23128 16212 23180
rect 16264 23168 16270 23180
rect 17129 23171 17187 23177
rect 17129 23168 17141 23171
rect 16264 23140 17141 23168
rect 16264 23128 16270 23140
rect 17129 23137 17141 23140
rect 17175 23168 17187 23171
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 17175 23140 19441 23168
rect 17175 23137 17187 23140
rect 17129 23131 17187 23137
rect 19429 23137 19441 23140
rect 19475 23168 19487 23171
rect 19702 23168 19708 23180
rect 19475 23140 19708 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 19702 23128 19708 23140
rect 19760 23128 19766 23180
rect 21358 23168 21364 23180
rect 20824 23140 21364 23168
rect 20824 23112 20852 23140
rect 21358 23128 21364 23140
rect 21416 23128 21422 23180
rect 23658 23128 23664 23180
rect 23716 23128 23722 23180
rect 25222 23128 25228 23180
rect 25280 23128 25286 23180
rect 27154 23128 27160 23180
rect 27212 23168 27218 23180
rect 29822 23168 29828 23180
rect 27212 23140 29828 23168
rect 27212 23128 27218 23140
rect 29822 23128 29828 23140
rect 29880 23168 29886 23180
rect 30101 23171 30159 23177
rect 30101 23168 30113 23171
rect 29880 23140 30113 23168
rect 29880 23128 29886 23140
rect 30101 23137 30113 23140
rect 30147 23168 30159 23171
rect 34885 23171 34943 23177
rect 30147 23140 31754 23168
rect 30147 23137 30159 23140
rect 30101 23131 30159 23137
rect 1811 23072 3556 23100
rect 4157 23103 4215 23109
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 4157 23069 4169 23103
rect 4203 23100 4215 23103
rect 4890 23100 4896 23112
rect 4203 23072 4896 23100
rect 4203 23069 4215 23072
rect 4157 23063 4215 23069
rect 4890 23060 4896 23072
rect 4948 23060 4954 23112
rect 9176 23103 9234 23109
rect 9176 23069 9188 23103
rect 9222 23100 9234 23103
rect 9766 23100 9772 23112
rect 9222 23072 9772 23100
rect 9222 23069 9234 23072
rect 9176 23063 9234 23069
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 20806 23060 20812 23112
rect 20864 23060 20870 23112
rect 23385 23103 23443 23109
rect 23385 23069 23397 23103
rect 23431 23100 23443 23103
rect 24854 23100 24860 23112
rect 23431 23072 24860 23100
rect 23431 23069 23443 23072
rect 23385 23063 23443 23069
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 24946 23060 24952 23112
rect 25004 23060 25010 23112
rect 28534 23060 28540 23112
rect 28592 23100 28598 23112
rect 28810 23100 28816 23112
rect 28592 23072 28816 23100
rect 28592 23060 28598 23072
rect 28810 23060 28816 23072
rect 28868 23060 28874 23112
rect 31726 23100 31754 23140
rect 34885 23137 34897 23171
rect 34931 23168 34943 23171
rect 37550 23168 37556 23180
rect 34931 23140 37556 23168
rect 34931 23137 34943 23140
rect 34885 23131 34943 23137
rect 37550 23128 37556 23140
rect 37608 23128 37614 23180
rect 38746 23128 38752 23180
rect 38804 23168 38810 23180
rect 38841 23171 38899 23177
rect 38841 23168 38853 23171
rect 38804 23140 38853 23168
rect 38804 23128 38810 23140
rect 38841 23137 38853 23140
rect 38887 23168 38899 23171
rect 39390 23168 39396 23180
rect 38887 23140 39396 23168
rect 38887 23137 38899 23140
rect 38841 23131 38899 23137
rect 39390 23128 39396 23140
rect 39448 23128 39454 23180
rect 32309 23103 32367 23109
rect 32309 23100 32321 23103
rect 31726 23072 32321 23100
rect 32309 23069 32321 23072
rect 32355 23069 32367 23103
rect 32309 23063 32367 23069
rect 5077 23035 5135 23041
rect 5077 23001 5089 23035
rect 5123 23032 5135 23035
rect 9674 23032 9680 23044
rect 5123 23004 9680 23032
rect 5123 23001 5135 23004
rect 5077 22995 5135 23001
rect 9674 22992 9680 23004
rect 9732 22992 9738 23044
rect 15286 22992 15292 23044
rect 15344 23032 15350 23044
rect 16206 23032 16212 23044
rect 15344 23004 16212 23032
rect 15344 22992 15350 23004
rect 16206 22992 16212 23004
rect 16264 22992 16270 23044
rect 17402 22992 17408 23044
rect 17460 22992 17466 23044
rect 17788 23004 17894 23032
rect 18800 23004 19334 23032
rect 2774 22924 2780 22976
rect 2832 22964 2838 22976
rect 4249 22967 4307 22973
rect 4249 22964 4261 22967
rect 2832 22936 4261 22964
rect 2832 22924 2838 22936
rect 4249 22933 4261 22936
rect 4295 22933 4307 22967
rect 16224 22964 16252 22992
rect 17788 22964 17816 23004
rect 18800 22964 18828 23004
rect 16224 22936 18828 22964
rect 4249 22927 4307 22933
rect 18874 22924 18880 22976
rect 18932 22924 18938 22976
rect 19306 22964 19334 23004
rect 19702 22992 19708 23044
rect 19760 22992 19766 23044
rect 20824 22964 20852 23060
rect 22186 22992 22192 23044
rect 22244 23032 22250 23044
rect 22738 23032 22744 23044
rect 22244 23004 22744 23032
rect 22244 22992 22250 23004
rect 22738 22992 22744 23004
rect 22796 23032 22802 23044
rect 23477 23035 23535 23041
rect 23477 23032 23489 23035
rect 22796 23004 23489 23032
rect 22796 22992 22802 23004
rect 23477 23001 23489 23004
rect 23523 23001 23535 23035
rect 23477 22995 23535 23001
rect 24762 22992 24768 23044
rect 24820 23032 24826 23044
rect 27433 23035 27491 23041
rect 24820 23004 27384 23032
rect 24820 22992 24826 23004
rect 19306 22936 20852 22964
rect 21174 22924 21180 22976
rect 21232 22924 21238 22976
rect 22646 22924 22652 22976
rect 22704 22964 22710 22976
rect 23017 22967 23075 22973
rect 23017 22964 23029 22967
rect 22704 22936 23029 22964
rect 22704 22924 22710 22936
rect 23017 22933 23029 22936
rect 23063 22933 23075 22967
rect 23017 22927 23075 22933
rect 24581 22967 24639 22973
rect 24581 22933 24593 22967
rect 24627 22964 24639 22967
rect 24946 22964 24952 22976
rect 24627 22936 24952 22964
rect 24627 22933 24639 22936
rect 24581 22927 24639 22933
rect 24946 22924 24952 22936
rect 25004 22924 25010 22976
rect 25038 22924 25044 22976
rect 25096 22924 25102 22976
rect 27356 22964 27384 23004
rect 27433 23001 27445 23035
rect 27479 23032 27491 23035
rect 27522 23032 27528 23044
rect 27479 23004 27528 23032
rect 27479 23001 27491 23004
rect 27433 22995 27491 23001
rect 27522 22992 27528 23004
rect 27580 22992 27586 23044
rect 30377 23035 30435 23041
rect 30377 23001 30389 23035
rect 30423 23001 30435 23035
rect 31662 23032 31668 23044
rect 31602 23004 31668 23032
rect 30377 22995 30435 23001
rect 29270 22964 29276 22976
rect 27356 22936 29276 22964
rect 29270 22924 29276 22936
rect 29328 22924 29334 22976
rect 30392 22964 30420 22995
rect 31662 22992 31668 23004
rect 31720 23032 31726 23044
rect 32324 23032 32352 23063
rect 33686 23060 33692 23112
rect 33744 23060 33750 23112
rect 37645 23103 37703 23109
rect 37645 23100 37657 23103
rect 36464 23072 37657 23100
rect 32490 23032 32496 23044
rect 31720 23004 31892 23032
rect 32324 23004 32496 23032
rect 31720 22992 31726 23004
rect 31754 22964 31760 22976
rect 30392 22936 31760 22964
rect 31754 22924 31760 22936
rect 31812 22924 31818 22976
rect 31864 22964 31892 23004
rect 32490 22992 32496 23004
rect 32548 22992 32554 23044
rect 32582 22992 32588 23044
rect 32640 22992 32646 23044
rect 33594 22964 33600 22976
rect 31864 22936 33600 22964
rect 33594 22924 33600 22936
rect 33652 22964 33658 22976
rect 33704 22964 33732 23060
rect 35158 22992 35164 23044
rect 35216 22992 35222 23044
rect 35894 22992 35900 23044
rect 35952 22992 35958 23044
rect 33652 22936 33732 22964
rect 33652 22924 33658 22936
rect 35526 22924 35532 22976
rect 35584 22964 35590 22976
rect 36464 22964 36492 23072
rect 37645 23069 37657 23072
rect 37691 23069 37703 23103
rect 37645 23063 37703 23069
rect 38565 23103 38623 23109
rect 38565 23069 38577 23103
rect 38611 23100 38623 23103
rect 40221 23103 40279 23109
rect 40221 23100 40233 23103
rect 38611 23072 40233 23100
rect 38611 23069 38623 23072
rect 38565 23063 38623 23069
rect 40221 23069 40233 23072
rect 40267 23069 40279 23103
rect 40221 23063 40279 23069
rect 47670 23060 47676 23112
rect 47728 23100 47734 23112
rect 47949 23103 48007 23109
rect 47949 23100 47961 23103
rect 47728 23072 47961 23100
rect 47728 23060 47734 23072
rect 47949 23069 47961 23072
rect 47995 23069 48007 23103
rect 47949 23063 48007 23069
rect 37458 22992 37464 23044
rect 37516 23032 37522 23044
rect 38657 23035 38715 23041
rect 38657 23032 38669 23035
rect 37516 23004 38669 23032
rect 37516 22992 37522 23004
rect 38657 23001 38669 23004
rect 38703 23001 38715 23035
rect 38657 22995 38715 23001
rect 49142 22992 49148 23044
rect 49200 22992 49206 23044
rect 35584 22936 36492 22964
rect 38197 22967 38255 22973
rect 35584 22924 35590 22936
rect 38197 22933 38209 22967
rect 38243 22964 38255 22967
rect 38286 22964 38292 22976
rect 38243 22936 38292 22964
rect 38243 22933 38255 22936
rect 38197 22927 38255 22933
rect 38286 22924 38292 22936
rect 38344 22924 38350 22976
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 17773 22763 17831 22769
rect 17773 22729 17785 22763
rect 17819 22760 17831 22763
rect 19429 22763 19487 22769
rect 19429 22760 19441 22763
rect 17819 22732 19441 22760
rect 17819 22729 17831 22732
rect 17773 22723 17831 22729
rect 19429 22729 19441 22732
rect 19475 22729 19487 22763
rect 19429 22723 19487 22729
rect 19797 22763 19855 22769
rect 19797 22729 19809 22763
rect 19843 22760 19855 22763
rect 22278 22760 22284 22772
rect 19843 22732 22284 22760
rect 19843 22729 19855 22732
rect 19797 22723 19855 22729
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 23658 22720 23664 22772
rect 23716 22720 23722 22772
rect 24946 22720 24952 22772
rect 25004 22760 25010 22772
rect 30009 22763 30067 22769
rect 30009 22760 30021 22763
rect 25004 22732 30021 22760
rect 25004 22720 25010 22732
rect 30009 22729 30021 22732
rect 30055 22729 30067 22763
rect 30009 22723 30067 22729
rect 30101 22763 30159 22769
rect 30101 22729 30113 22763
rect 30147 22760 30159 22763
rect 30374 22760 30380 22772
rect 30147 22732 30380 22760
rect 30147 22729 30159 22732
rect 30101 22723 30159 22729
rect 30374 22720 30380 22732
rect 30432 22720 30438 22772
rect 31021 22763 31079 22769
rect 31021 22729 31033 22763
rect 31067 22760 31079 22763
rect 32674 22760 32680 22772
rect 31067 22732 32680 22760
rect 31067 22729 31079 22732
rect 31021 22723 31079 22729
rect 32674 22720 32680 22732
rect 32732 22720 32738 22772
rect 34057 22763 34115 22769
rect 34057 22729 34069 22763
rect 34103 22760 34115 22763
rect 34514 22760 34520 22772
rect 34103 22732 34520 22760
rect 34103 22729 34115 22732
rect 34057 22723 34115 22729
rect 34514 22720 34520 22732
rect 34572 22720 34578 22772
rect 37550 22720 37556 22772
rect 37608 22760 37614 22772
rect 38562 22760 38568 22772
rect 37608 22732 38568 22760
rect 37608 22720 37614 22732
rect 38562 22720 38568 22732
rect 38620 22720 38626 22772
rect 17402 22652 17408 22704
rect 17460 22692 17466 22704
rect 21177 22695 21235 22701
rect 17460 22664 20024 22692
rect 17460 22652 17466 22664
rect 16482 22584 16488 22636
rect 16540 22624 16546 22636
rect 18874 22624 18880 22636
rect 16540 22596 18880 22624
rect 16540 22584 16546 22596
rect 17972 22565 18000 22596
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 17865 22559 17923 22565
rect 17865 22525 17877 22559
rect 17911 22525 17923 22559
rect 17865 22519 17923 22525
rect 17957 22559 18015 22565
rect 17957 22525 17969 22559
rect 18003 22525 18015 22559
rect 17957 22519 18015 22525
rect 17880 22488 17908 22519
rect 19886 22516 19892 22568
rect 19944 22516 19950 22568
rect 19996 22565 20024 22664
rect 21177 22661 21189 22695
rect 21223 22692 21235 22695
rect 23382 22692 23388 22704
rect 21223 22664 23388 22692
rect 21223 22661 21235 22664
rect 21177 22655 21235 22661
rect 23382 22652 23388 22664
rect 23440 22652 23446 22704
rect 23676 22692 23704 22720
rect 23753 22695 23811 22701
rect 23753 22692 23765 22695
rect 23676 22664 23765 22692
rect 23753 22661 23765 22664
rect 23799 22692 23811 22695
rect 26878 22692 26884 22704
rect 23799 22664 26884 22692
rect 23799 22661 23811 22664
rect 23753 22655 23811 22661
rect 26878 22652 26884 22664
rect 26936 22652 26942 22704
rect 28810 22652 28816 22704
rect 28868 22692 28874 22704
rect 28868 22664 30420 22692
rect 28868 22652 28874 22664
rect 30392 22636 30420 22664
rect 30466 22652 30472 22704
rect 30524 22692 30530 22704
rect 31481 22695 31539 22701
rect 31481 22692 31493 22695
rect 30524 22664 31493 22692
rect 30524 22652 30530 22664
rect 31481 22661 31493 22664
rect 31527 22692 31539 22695
rect 31527 22664 34100 22692
rect 31527 22661 31539 22664
rect 31481 22655 31539 22661
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22624 21143 22627
rect 23290 22624 23296 22636
rect 21131 22596 23296 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 23290 22584 23296 22596
rect 23348 22584 23354 22636
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22624 23719 22627
rect 24762 22624 24768 22636
rect 23707 22596 24768 22624
rect 23707 22593 23719 22596
rect 23661 22587 23719 22593
rect 24762 22584 24768 22596
rect 24820 22584 24826 22636
rect 24949 22627 25007 22633
rect 24949 22593 24961 22627
rect 24995 22624 25007 22627
rect 25961 22627 26019 22633
rect 25961 22624 25973 22627
rect 24995 22596 25973 22624
rect 24995 22593 25007 22596
rect 24949 22587 25007 22593
rect 25961 22593 25973 22596
rect 26007 22593 26019 22627
rect 25961 22587 26019 22593
rect 27154 22584 27160 22636
rect 27212 22584 27218 22636
rect 28534 22584 28540 22636
rect 28592 22584 28598 22636
rect 28920 22596 30236 22624
rect 19981 22559 20039 22565
rect 19981 22525 19993 22559
rect 20027 22556 20039 22559
rect 21174 22556 21180 22568
rect 20027 22528 21180 22556
rect 20027 22525 20039 22528
rect 19981 22519 20039 22525
rect 21174 22516 21180 22528
rect 21232 22556 21238 22568
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 21232 22528 21281 22556
rect 21232 22516 21238 22528
rect 21269 22525 21281 22528
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 23937 22559 23995 22565
rect 23937 22525 23949 22559
rect 23983 22556 23995 22559
rect 25041 22559 25099 22565
rect 23983 22528 24992 22556
rect 23983 22525 23995 22528
rect 23937 22519 23995 22525
rect 20717 22491 20775 22497
rect 20717 22488 20729 22491
rect 17880 22460 20729 22488
rect 20717 22457 20729 22460
rect 20763 22457 20775 22491
rect 20717 22451 20775 22457
rect 21358 22448 21364 22500
rect 21416 22488 21422 22500
rect 24581 22491 24639 22497
rect 24581 22488 24593 22491
rect 21416 22460 24593 22488
rect 21416 22448 21422 22460
rect 24581 22457 24593 22460
rect 24627 22457 24639 22491
rect 24964 22488 24992 22528
rect 25041 22525 25053 22559
rect 25087 22556 25099 22559
rect 25225 22559 25283 22565
rect 25087 22528 25176 22556
rect 25087 22525 25099 22528
rect 25041 22519 25099 22525
rect 25148 22488 25176 22528
rect 25225 22525 25237 22559
rect 25271 22556 25283 22559
rect 25498 22556 25504 22568
rect 25271 22528 25504 22556
rect 25271 22525 25283 22528
rect 25225 22519 25283 22525
rect 25498 22516 25504 22528
rect 25556 22516 25562 22568
rect 27522 22516 27528 22568
rect 27580 22556 27586 22568
rect 28920 22565 28948 22596
rect 30208 22565 30236 22596
rect 30374 22584 30380 22636
rect 30432 22584 30438 22636
rect 31389 22627 31447 22633
rect 31389 22593 31401 22627
rect 31435 22624 31447 22627
rect 32493 22627 32551 22633
rect 32493 22624 32505 22627
rect 31435 22596 32505 22624
rect 31435 22593 31447 22596
rect 31389 22587 31447 22593
rect 32493 22593 32505 22596
rect 32539 22593 32551 22627
rect 34072 22624 34100 22664
rect 34146 22652 34152 22704
rect 34204 22652 34210 22704
rect 37366 22624 37372 22636
rect 34072 22596 37372 22624
rect 32493 22587 32551 22593
rect 37366 22584 37372 22596
rect 37424 22584 37430 22636
rect 37568 22633 37596 22720
rect 39574 22692 39580 22704
rect 39054 22678 39580 22692
rect 39040 22664 39580 22678
rect 37553 22627 37611 22633
rect 37553 22593 37565 22627
rect 37599 22593 37611 22627
rect 37553 22587 37611 22593
rect 39040 22568 39068 22664
rect 39574 22652 39580 22664
rect 39632 22652 39638 22704
rect 42794 22652 42800 22704
rect 42852 22692 42858 22704
rect 44269 22695 44327 22701
rect 44269 22692 44281 22695
rect 42852 22664 44281 22692
rect 42852 22652 42858 22664
rect 44269 22661 44281 22664
rect 44315 22661 44327 22695
rect 44269 22655 44327 22661
rect 28905 22559 28963 22565
rect 28905 22556 28917 22559
rect 27580 22528 28917 22556
rect 27580 22516 27586 22528
rect 28905 22525 28917 22528
rect 28951 22525 28963 22559
rect 28905 22519 28963 22525
rect 30193 22559 30251 22565
rect 30193 22525 30205 22559
rect 30239 22525 30251 22559
rect 30193 22519 30251 22525
rect 31665 22559 31723 22565
rect 31665 22525 31677 22559
rect 31711 22556 31723 22559
rect 32858 22556 32864 22568
rect 31711 22528 32864 22556
rect 31711 22525 31723 22528
rect 31665 22519 31723 22525
rect 32858 22516 32864 22528
rect 32916 22516 32922 22568
rect 34238 22516 34244 22568
rect 34296 22516 34302 22568
rect 37826 22516 37832 22568
rect 37884 22516 37890 22568
rect 39022 22516 39028 22568
rect 39080 22516 39086 22568
rect 39482 22516 39488 22568
rect 39540 22556 39546 22568
rect 39577 22559 39635 22565
rect 39577 22556 39589 22559
rect 39540 22528 39589 22556
rect 39540 22516 39546 22528
rect 39577 22525 39589 22528
rect 39623 22525 39635 22559
rect 39577 22519 39635 22525
rect 26510 22488 26516 22500
rect 24964 22460 25084 22488
rect 25148 22460 26516 22488
rect 24581 22451 24639 22457
rect 25056 22432 25084 22460
rect 26510 22448 26516 22460
rect 26568 22448 26574 22500
rect 29641 22491 29699 22497
rect 29641 22457 29653 22491
rect 29687 22488 29699 22491
rect 36906 22488 36912 22500
rect 29687 22460 36912 22488
rect 29687 22457 29699 22460
rect 29641 22451 29699 22457
rect 36906 22448 36912 22460
rect 36964 22448 36970 22500
rect 44453 22491 44511 22497
rect 44453 22457 44465 22491
rect 44499 22488 44511 22491
rect 46750 22488 46756 22500
rect 44499 22460 46756 22488
rect 44499 22457 44511 22460
rect 44453 22451 44511 22457
rect 46750 22448 46756 22460
rect 46808 22448 46814 22500
rect 13354 22380 13360 22432
rect 13412 22420 13418 22432
rect 16574 22420 16580 22432
rect 13412 22392 16580 22420
rect 13412 22380 13418 22392
rect 16574 22380 16580 22392
rect 16632 22380 16638 22432
rect 17402 22380 17408 22432
rect 17460 22380 17466 22432
rect 21174 22380 21180 22432
rect 21232 22420 21238 22432
rect 23293 22423 23351 22429
rect 23293 22420 23305 22423
rect 21232 22392 23305 22420
rect 21232 22380 21238 22392
rect 23293 22389 23305 22392
rect 23339 22389 23351 22423
rect 23293 22383 23351 22389
rect 25038 22380 25044 22432
rect 25096 22380 25102 22432
rect 25222 22380 25228 22432
rect 25280 22420 25286 22432
rect 27420 22423 27478 22429
rect 27420 22420 27432 22423
rect 25280 22392 27432 22420
rect 25280 22380 25286 22392
rect 27420 22389 27432 22392
rect 27466 22420 27478 22423
rect 31294 22420 31300 22432
rect 27466 22392 31300 22420
rect 27466 22389 27478 22392
rect 27420 22383 27478 22389
rect 31294 22380 31300 22392
rect 31352 22380 31358 22432
rect 32306 22380 32312 22432
rect 32364 22420 32370 22432
rect 33689 22423 33747 22429
rect 33689 22420 33701 22423
rect 32364 22392 33701 22420
rect 32364 22380 32370 22392
rect 33689 22389 33701 22392
rect 33735 22389 33747 22423
rect 33689 22383 33747 22389
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 12897 22219 12955 22225
rect 12897 22185 12909 22219
rect 12943 22216 12955 22219
rect 13354 22216 13360 22228
rect 12943 22188 13360 22216
rect 12943 22185 12955 22188
rect 12897 22179 12955 22185
rect 13354 22176 13360 22188
rect 13412 22176 13418 22228
rect 15086 22219 15144 22225
rect 15086 22216 15098 22219
rect 14936 22188 15098 22216
rect 5534 22108 5540 22160
rect 5592 22108 5598 22160
rect 14090 22108 14096 22160
rect 14148 22148 14154 22160
rect 14936 22148 14964 22188
rect 15086 22185 15098 22188
rect 15132 22185 15144 22219
rect 15086 22179 15144 22185
rect 23290 22176 23296 22228
rect 23348 22176 23354 22228
rect 23676 22188 24900 22216
rect 14148 22120 14964 22148
rect 14148 22108 14154 22120
rect 16482 22108 16488 22160
rect 16540 22108 16546 22160
rect 21082 22108 21088 22160
rect 21140 22148 21146 22160
rect 21140 22120 21496 22148
rect 21140 22108 21146 22120
rect 16500 22080 16528 22108
rect 21468 22089 21496 22120
rect 22554 22108 22560 22160
rect 22612 22148 22618 22160
rect 22612 22120 22692 22148
rect 22612 22108 22618 22120
rect 22664 22089 22692 22120
rect 13740 22052 16528 22080
rect 21453 22083 21511 22089
rect 9122 21972 9128 22024
rect 9180 22012 9186 22024
rect 9180 21984 12572 22012
rect 9180 21972 9186 21984
rect 5353 21947 5411 21953
rect 5353 21913 5365 21947
rect 5399 21944 5411 21947
rect 10226 21944 10232 21956
rect 5399 21916 10232 21944
rect 5399 21913 5411 21916
rect 5353 21907 5411 21913
rect 10226 21904 10232 21916
rect 10284 21904 10290 21956
rect 12544 21944 12572 21984
rect 12618 21972 12624 22024
rect 12676 21972 12682 22024
rect 13740 22021 13768 22052
rect 21453 22049 21465 22083
rect 21499 22049 21511 22083
rect 21453 22043 21511 22049
rect 22649 22083 22707 22089
rect 22649 22049 22661 22083
rect 22695 22049 22707 22083
rect 22649 22043 22707 22049
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 21981 13783 22015
rect 13725 21975 13783 21981
rect 14826 21972 14832 22024
rect 14884 21972 14890 22024
rect 16206 21972 16212 22024
rect 16264 21972 16270 22024
rect 16408 22012 16528 22022
rect 23676 22012 23704 22188
rect 24872 22148 24900 22188
rect 25038 22176 25044 22228
rect 25096 22216 25102 22228
rect 26602 22216 26608 22228
rect 25096 22188 26608 22216
rect 25096 22176 25102 22188
rect 26602 22176 26608 22188
rect 26660 22176 26666 22228
rect 31754 22216 31760 22228
rect 26712 22188 31760 22216
rect 25133 22151 25191 22157
rect 25133 22148 25145 22151
rect 24872 22120 25145 22148
rect 25133 22117 25145 22120
rect 25179 22117 25191 22151
rect 25133 22111 25191 22117
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22080 23995 22083
rect 24210 22080 24216 22092
rect 23983 22052 24216 22080
rect 23983 22049 23995 22052
rect 23937 22043 23995 22049
rect 24210 22040 24216 22052
rect 24268 22040 24274 22092
rect 25148 22080 25176 22111
rect 25222 22108 25228 22160
rect 25280 22148 25286 22160
rect 25590 22148 25596 22160
rect 25280 22120 25596 22148
rect 25280 22108 25286 22120
rect 25590 22108 25596 22120
rect 25648 22108 25654 22160
rect 26712 22148 26740 22188
rect 31754 22176 31760 22188
rect 31812 22216 31818 22228
rect 32674 22216 32680 22228
rect 31812 22188 32680 22216
rect 31812 22176 31818 22188
rect 32674 22176 32680 22188
rect 32732 22176 32738 22228
rect 34238 22176 34244 22228
rect 34296 22216 34302 22228
rect 35602 22219 35660 22225
rect 35602 22216 35614 22219
rect 34296 22188 35614 22216
rect 34296 22176 34302 22188
rect 35602 22185 35614 22188
rect 35648 22185 35660 22219
rect 35602 22179 35660 22185
rect 26528 22120 26740 22148
rect 25774 22080 25780 22092
rect 25148 22052 25780 22080
rect 25774 22040 25780 22052
rect 25832 22080 25838 22092
rect 26053 22083 26111 22089
rect 26053 22080 26065 22083
rect 25832 22052 26065 22080
rect 25832 22040 25838 22052
rect 26053 22049 26065 22052
rect 26099 22049 26111 22083
rect 26053 22043 26111 22049
rect 26237 22083 26295 22089
rect 26237 22049 26249 22083
rect 26283 22080 26295 22083
rect 26528 22080 26556 22120
rect 26878 22108 26884 22160
rect 26936 22148 26942 22160
rect 26936 22120 29040 22148
rect 26936 22108 26942 22120
rect 26283 22052 26556 22080
rect 26283 22049 26295 22052
rect 26237 22043 26295 22049
rect 27798 22040 27804 22092
rect 27856 22080 27862 22092
rect 29012 22089 29040 22120
rect 30374 22108 30380 22160
rect 30432 22148 30438 22160
rect 31662 22148 31668 22160
rect 30432 22120 31668 22148
rect 30432 22108 30438 22120
rect 31662 22108 31668 22120
rect 31720 22108 31726 22160
rect 33502 22108 33508 22160
rect 33560 22148 33566 22160
rect 34422 22148 34428 22160
rect 33560 22120 34428 22148
rect 33560 22108 33566 22120
rect 34422 22108 34428 22120
rect 34480 22108 34486 22160
rect 28997 22083 29055 22089
rect 27856 22052 28580 22080
rect 27856 22040 27862 22052
rect 16408 21994 23704 22012
rect 12544 21916 15516 21944
rect 9306 21836 9312 21888
rect 9364 21876 9370 21888
rect 13081 21879 13139 21885
rect 13081 21876 13093 21879
rect 9364 21848 13093 21876
rect 9364 21836 9370 21848
rect 13081 21845 13093 21848
rect 13127 21845 13139 21879
rect 13081 21839 13139 21845
rect 13538 21836 13544 21888
rect 13596 21836 13602 21888
rect 15488 21876 15516 21916
rect 16408 21876 16436 21994
rect 16500 21984 23704 21994
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 22012 23811 22015
rect 25961 22015 26019 22021
rect 23799 21984 25912 22012
rect 23799 21981 23811 21984
rect 23753 21975 23811 21981
rect 16482 21904 16488 21956
rect 16540 21944 16546 21956
rect 17402 21944 17408 21956
rect 16540 21916 17408 21944
rect 16540 21904 16546 21916
rect 17402 21904 17408 21916
rect 17460 21904 17466 21956
rect 20714 21904 20720 21956
rect 20772 21944 20778 21956
rect 20990 21944 20996 21956
rect 20772 21916 20996 21944
rect 20772 21904 20778 21916
rect 20990 21904 20996 21916
rect 21048 21944 21054 21956
rect 21269 21947 21327 21953
rect 21269 21944 21281 21947
rect 21048 21916 21281 21944
rect 21048 21904 21054 21916
rect 21269 21913 21281 21916
rect 21315 21913 21327 21947
rect 21269 21907 21327 21913
rect 21361 21947 21419 21953
rect 21361 21913 21373 21947
rect 21407 21944 21419 21947
rect 22278 21944 22284 21956
rect 21407 21916 22284 21944
rect 21407 21913 21419 21916
rect 21361 21907 21419 21913
rect 22278 21904 22284 21916
rect 22336 21904 22342 21956
rect 22465 21947 22523 21953
rect 22465 21913 22477 21947
rect 22511 21944 22523 21947
rect 23566 21944 23572 21956
rect 22511 21916 23572 21944
rect 22511 21913 22523 21916
rect 22465 21907 22523 21913
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 23661 21947 23719 21953
rect 23661 21913 23673 21947
rect 23707 21944 23719 21947
rect 23842 21944 23848 21956
rect 23707 21916 23848 21944
rect 23707 21913 23719 21916
rect 23661 21907 23719 21913
rect 23842 21904 23848 21916
rect 23900 21904 23906 21956
rect 25884 21944 25912 21984
rect 25961 21981 25973 22015
rect 26007 22012 26019 22015
rect 28442 22012 28448 22024
rect 26007 21984 28448 22012
rect 26007 21981 26019 21984
rect 25961 21975 26019 21981
rect 28442 21972 28448 21984
rect 28500 21972 28506 22024
rect 28552 22012 28580 22052
rect 28997 22049 29009 22083
rect 29043 22049 29055 22083
rect 28997 22043 29055 22049
rect 29840 22052 30052 22080
rect 29840 22012 29868 22052
rect 28552 21984 29868 22012
rect 29914 21972 29920 22024
rect 29972 21972 29978 22024
rect 30024 22012 30052 22052
rect 31110 22040 31116 22092
rect 31168 22080 31174 22092
rect 37093 22083 37151 22089
rect 31168 22052 36860 22080
rect 31168 22040 31174 22052
rect 30024 21984 32615 22012
rect 26786 21944 26792 21956
rect 25884 21916 26792 21944
rect 26786 21904 26792 21916
rect 26844 21904 26850 21956
rect 28813 21947 28871 21953
rect 28813 21913 28825 21947
rect 28859 21944 28871 21947
rect 32587 21944 32615 21984
rect 32858 21972 32864 22024
rect 32916 22012 32922 22024
rect 35345 22015 35403 22021
rect 35345 22012 35357 22015
rect 32916 21984 35357 22012
rect 32916 21972 32922 21984
rect 35345 21981 35357 21984
rect 35391 21981 35403 22015
rect 36832 22012 36860 22052
rect 37093 22049 37105 22083
rect 37139 22080 37151 22083
rect 37458 22080 37464 22092
rect 37139 22052 37464 22080
rect 37139 22049 37151 22052
rect 37093 22043 37151 22049
rect 37458 22040 37464 22052
rect 37516 22040 37522 22092
rect 37829 22015 37887 22021
rect 37829 22012 37841 22015
rect 36832 21984 37841 22012
rect 35345 21975 35403 21981
rect 37829 21981 37841 21984
rect 37875 21981 37887 22015
rect 37829 21975 37887 21981
rect 47578 21972 47584 22024
rect 47636 22012 47642 22024
rect 47949 22015 48007 22021
rect 47949 22012 47961 22015
rect 47636 21984 47961 22012
rect 47636 21972 47642 21984
rect 47949 21981 47961 21984
rect 47995 21981 48007 22015
rect 47949 21975 48007 21981
rect 49142 21972 49148 22024
rect 49200 21972 49206 22024
rect 35250 21944 35256 21956
rect 28859 21916 30328 21944
rect 32587 21916 35256 21944
rect 28859 21913 28871 21916
rect 28813 21907 28871 21913
rect 15488 21848 16436 21876
rect 16574 21836 16580 21888
rect 16632 21836 16638 21888
rect 20898 21836 20904 21888
rect 20956 21836 20962 21888
rect 22094 21836 22100 21888
rect 22152 21836 22158 21888
rect 22557 21879 22615 21885
rect 22557 21845 22569 21879
rect 22603 21876 22615 21879
rect 24946 21876 24952 21888
rect 22603 21848 24952 21876
rect 22603 21845 22615 21848
rect 22557 21839 22615 21845
rect 24946 21836 24952 21848
rect 25004 21836 25010 21888
rect 25590 21836 25596 21888
rect 25648 21836 25654 21888
rect 26418 21836 26424 21888
rect 26476 21876 26482 21888
rect 28445 21879 28503 21885
rect 28445 21876 28457 21879
rect 26476 21848 28457 21876
rect 26476 21836 26482 21848
rect 28445 21845 28457 21848
rect 28491 21845 28503 21879
rect 28445 21839 28503 21845
rect 28718 21836 28724 21888
rect 28776 21876 28782 21888
rect 28905 21879 28963 21885
rect 28905 21876 28917 21879
rect 28776 21848 28917 21876
rect 28776 21836 28782 21848
rect 28905 21845 28917 21848
rect 28951 21845 28963 21879
rect 30300 21876 30328 21916
rect 35250 21904 35256 21916
rect 35308 21904 35314 21956
rect 36078 21904 36084 21956
rect 36136 21904 36142 21956
rect 32122 21876 32128 21888
rect 30300 21848 32128 21876
rect 28905 21839 28963 21845
rect 32122 21836 32128 21848
rect 32180 21836 32186 21888
rect 37645 21879 37703 21885
rect 37645 21845 37657 21879
rect 37691 21876 37703 21879
rect 44174 21876 44180 21888
rect 37691 21848 44180 21876
rect 37691 21845 37703 21848
rect 37645 21839 37703 21845
rect 44174 21836 44180 21848
rect 44232 21836 44238 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 10226 21632 10232 21684
rect 10284 21632 10290 21684
rect 12158 21632 12164 21684
rect 12216 21672 12222 21684
rect 14277 21675 14335 21681
rect 14277 21672 14289 21675
rect 12216 21644 14289 21672
rect 12216 21632 12222 21644
rect 14277 21641 14289 21644
rect 14323 21641 14335 21675
rect 14277 21635 14335 21641
rect 23566 21632 23572 21684
rect 23624 21672 23630 21684
rect 25133 21675 25191 21681
rect 25133 21672 25145 21675
rect 23624 21644 25145 21672
rect 23624 21632 23630 21644
rect 25133 21641 25145 21644
rect 25179 21641 25191 21675
rect 25133 21635 25191 21641
rect 25501 21675 25559 21681
rect 25501 21641 25513 21675
rect 25547 21672 25559 21675
rect 25866 21672 25872 21684
rect 25547 21644 25872 21672
rect 25547 21641 25559 21644
rect 25501 21635 25559 21641
rect 25866 21632 25872 21644
rect 25924 21632 25930 21684
rect 28997 21675 29055 21681
rect 28997 21641 29009 21675
rect 29043 21672 29055 21675
rect 29914 21672 29920 21684
rect 29043 21644 29920 21672
rect 29043 21641 29055 21644
rect 28997 21635 29055 21641
rect 29914 21632 29920 21644
rect 29972 21632 29978 21684
rect 30466 21632 30472 21684
rect 30524 21672 30530 21684
rect 31573 21675 31631 21681
rect 30524 21644 31432 21672
rect 30524 21632 30530 21644
rect 19610 21604 19616 21616
rect 19260 21576 19616 21604
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 13538 21536 13544 21548
rect 9631 21508 13544 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 13538 21496 13544 21508
rect 13596 21496 13602 21548
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21505 14519 21539
rect 14461 21499 14519 21505
rect 9766 21428 9772 21480
rect 9824 21428 9830 21480
rect 14476 21468 14504 21499
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 19260 21545 19288 21576
rect 19610 21564 19616 21576
rect 19668 21564 19674 21616
rect 20806 21604 20812 21616
rect 20746 21576 20812 21604
rect 20806 21564 20812 21576
rect 20864 21564 20870 21616
rect 23474 21564 23480 21616
rect 23532 21564 23538 21616
rect 25590 21564 25596 21616
rect 25648 21604 25654 21616
rect 29089 21607 29147 21613
rect 29089 21604 29101 21607
rect 25648 21576 29101 21604
rect 25648 21564 25654 21576
rect 29089 21573 29101 21576
rect 29135 21573 29147 21607
rect 30190 21604 30196 21616
rect 29089 21567 29147 21573
rect 29840 21576 30196 21604
rect 19245 21539 19303 21545
rect 19245 21536 19257 21539
rect 14884 21508 19257 21536
rect 14884 21496 14890 21508
rect 19245 21505 19257 21508
rect 19291 21505 19303 21539
rect 19245 21499 19303 21505
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 28169 21539 28227 21545
rect 25188 21508 25728 21536
rect 25188 21496 25194 21508
rect 16022 21468 16028 21480
rect 14476 21440 16028 21468
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 19521 21471 19579 21477
rect 19521 21437 19533 21471
rect 19567 21468 19579 21471
rect 19567 21440 22094 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 19518 21292 19524 21344
rect 19576 21332 19582 21344
rect 20993 21335 21051 21341
rect 20993 21332 21005 21335
rect 19576 21304 21005 21332
rect 19576 21292 19582 21304
rect 20993 21301 21005 21304
rect 21039 21301 21051 21335
rect 22066 21332 22094 21440
rect 22462 21428 22468 21480
rect 22520 21428 22526 21480
rect 22741 21471 22799 21477
rect 22741 21437 22753 21471
rect 22787 21468 22799 21471
rect 22830 21468 22836 21480
rect 22787 21440 22836 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 25590 21428 25596 21480
rect 25648 21428 25654 21480
rect 25700 21477 25728 21508
rect 28169 21505 28181 21539
rect 28215 21536 28227 21539
rect 28626 21536 28632 21548
rect 28215 21508 28632 21536
rect 28215 21505 28227 21508
rect 28169 21499 28227 21505
rect 28626 21496 28632 21508
rect 28684 21496 28690 21548
rect 29840 21536 29868 21576
rect 30190 21564 30196 21576
rect 30248 21564 30254 21616
rect 31404 21604 31432 21644
rect 31573 21641 31585 21675
rect 31619 21672 31631 21675
rect 31754 21672 31760 21684
rect 31619 21644 31760 21672
rect 31619 21641 31631 21644
rect 31573 21635 31631 21641
rect 31754 21632 31760 21644
rect 31812 21672 31818 21684
rect 32582 21672 32588 21684
rect 31812 21644 32588 21672
rect 31812 21632 31818 21644
rect 32582 21632 32588 21644
rect 32640 21632 32646 21684
rect 33152 21644 36032 21672
rect 33152 21604 33180 21644
rect 31404 21576 33180 21604
rect 33502 21564 33508 21616
rect 33560 21564 33566 21616
rect 31662 21536 31668 21548
rect 28966 21508 29868 21536
rect 31234 21508 31668 21536
rect 25685 21471 25743 21477
rect 25685 21437 25697 21471
rect 25731 21437 25743 21471
rect 25685 21431 25743 21437
rect 25774 21428 25780 21480
rect 25832 21468 25838 21480
rect 28966 21468 28994 21508
rect 31662 21496 31668 21508
rect 31720 21496 31726 21548
rect 32490 21496 32496 21548
rect 32548 21496 32554 21548
rect 35250 21496 35256 21548
rect 35308 21496 35314 21548
rect 36004 21545 36032 21644
rect 38746 21564 38752 21616
rect 38804 21564 38810 21616
rect 38838 21564 38844 21616
rect 38896 21604 38902 21616
rect 39022 21604 39028 21616
rect 38896 21576 39028 21604
rect 38896 21564 38902 21576
rect 39022 21564 39028 21576
rect 39080 21604 39086 21616
rect 39080 21576 39238 21604
rect 39080 21564 39086 21576
rect 35989 21539 36047 21545
rect 35989 21505 36001 21539
rect 36035 21505 36047 21539
rect 35989 21499 36047 21505
rect 38470 21496 38476 21548
rect 38528 21496 38534 21548
rect 46290 21496 46296 21548
rect 46348 21536 46354 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 46348 21508 47961 21536
rect 46348 21496 46354 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 25832 21440 28994 21468
rect 29273 21471 29331 21477
rect 25832 21428 25838 21440
rect 29273 21437 29285 21471
rect 29319 21437 29331 21471
rect 29273 21431 29331 21437
rect 29288 21400 29316 21431
rect 29822 21428 29828 21480
rect 29880 21428 29886 21480
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29932 21440 30113 21468
rect 29932 21400 29960 21440
rect 30101 21437 30113 21440
rect 30147 21468 30159 21471
rect 31846 21468 31852 21480
rect 30147 21440 31852 21468
rect 30147 21437 30159 21440
rect 30101 21431 30159 21437
rect 31846 21428 31852 21440
rect 31904 21428 31910 21480
rect 32214 21428 32220 21480
rect 32272 21468 32278 21480
rect 32769 21471 32827 21477
rect 32769 21468 32781 21471
rect 32272 21440 32781 21468
rect 32272 21428 32278 21440
rect 32769 21437 32781 21440
rect 32815 21468 32827 21471
rect 34054 21468 34060 21480
rect 32815 21440 34060 21468
rect 32815 21437 32827 21440
rect 32769 21431 32827 21437
rect 34054 21428 34060 21440
rect 34112 21428 34118 21480
rect 37826 21428 37832 21480
rect 37884 21468 37890 21480
rect 40221 21471 40279 21477
rect 40221 21468 40233 21471
rect 37884 21440 40233 21468
rect 37884 21428 37890 21440
rect 40221 21437 40233 21440
rect 40267 21437 40279 21471
rect 40221 21431 40279 21437
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 36814 21400 36820 21412
rect 29288 21372 29960 21400
rect 33796 21372 36820 21400
rect 23934 21332 23940 21344
rect 22066 21304 23940 21332
rect 20993 21295 21051 21301
rect 23934 21292 23940 21304
rect 23992 21292 23998 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 24762 21332 24768 21344
rect 24268 21304 24768 21332
rect 24268 21292 24274 21304
rect 24762 21292 24768 21304
rect 24820 21292 24826 21344
rect 27798 21292 27804 21344
rect 27856 21332 27862 21344
rect 27985 21335 28043 21341
rect 27985 21332 27997 21335
rect 27856 21304 27997 21332
rect 27856 21292 27862 21304
rect 27985 21301 27997 21304
rect 28031 21301 28043 21335
rect 27985 21295 28043 21301
rect 28629 21335 28687 21341
rect 28629 21301 28641 21335
rect 28675 21332 28687 21335
rect 30650 21332 30656 21344
rect 28675 21304 30656 21332
rect 28675 21301 28687 21304
rect 28629 21295 28687 21301
rect 30650 21292 30656 21304
rect 30708 21292 30714 21344
rect 32122 21292 32128 21344
rect 32180 21332 32186 21344
rect 33796 21332 33824 21372
rect 36814 21360 36820 21372
rect 36872 21360 36878 21412
rect 40144 21372 41414 21400
rect 32180 21304 33824 21332
rect 32180 21292 32186 21304
rect 34238 21292 34244 21344
rect 34296 21292 34302 21344
rect 35066 21292 35072 21344
rect 35124 21292 35130 21344
rect 35805 21335 35863 21341
rect 35805 21301 35817 21335
rect 35851 21332 35863 21335
rect 40144 21332 40172 21372
rect 35851 21304 40172 21332
rect 41386 21332 41414 21372
rect 43346 21332 43352 21344
rect 41386 21304 43352 21332
rect 35851 21301 35863 21304
rect 35805 21295 35863 21301
rect 43346 21292 43352 21304
rect 43404 21292 43410 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 9674 21088 9680 21140
rect 9732 21088 9738 21140
rect 19429 21131 19487 21137
rect 19429 21097 19441 21131
rect 19475 21128 19487 21131
rect 19886 21128 19892 21140
rect 19475 21100 19892 21128
rect 19475 21097 19487 21100
rect 19429 21091 19487 21097
rect 19886 21088 19892 21100
rect 19944 21088 19950 21140
rect 32490 21088 32496 21140
rect 32548 21128 32554 21140
rect 32858 21128 32864 21140
rect 32548 21100 32864 21128
rect 32548 21088 32554 21100
rect 32858 21088 32864 21100
rect 32916 21088 32922 21140
rect 35066 21088 35072 21140
rect 35124 21128 35130 21140
rect 42794 21128 42800 21140
rect 35124 21100 42800 21128
rect 35124 21088 35130 21100
rect 42794 21088 42800 21100
rect 42852 21088 42858 21140
rect 36633 21063 36691 21069
rect 36633 21029 36645 21063
rect 36679 21060 36691 21063
rect 43714 21060 43720 21072
rect 36679 21032 43720 21060
rect 36679 21029 36691 21032
rect 36633 21023 36691 21029
rect 43714 21020 43720 21032
rect 43772 21020 43778 21072
rect 9125 20995 9183 21001
rect 9125 20961 9137 20995
rect 9171 20992 9183 20995
rect 10962 20992 10968 21004
rect 9171 20964 10968 20992
rect 9171 20961 9183 20964
rect 9125 20955 9183 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 19702 20952 19708 21004
rect 19760 20992 19766 21004
rect 20073 20995 20131 21001
rect 20073 20992 20085 20995
rect 19760 20964 20085 20992
rect 19760 20952 19766 20964
rect 20073 20961 20085 20964
rect 20119 20992 20131 20995
rect 24210 20992 24216 21004
rect 20119 20964 24216 20992
rect 20119 20961 20131 20964
rect 20073 20955 20131 20961
rect 24210 20952 24216 20964
rect 24268 20952 24274 21004
rect 30929 20995 30987 21001
rect 30929 20961 30941 20995
rect 30975 20992 30987 20995
rect 31754 20992 31760 21004
rect 30975 20964 31760 20992
rect 30975 20961 30987 20964
rect 30929 20955 30987 20961
rect 31754 20952 31760 20964
rect 31812 20952 31818 21004
rect 34790 20992 34796 21004
rect 32324 20964 34796 20992
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 7834 20924 7840 20936
rect 4203 20896 7840 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19518 20924 19524 20936
rect 19392 20896 19524 20924
rect 19392 20884 19398 20896
rect 19518 20884 19524 20896
rect 19576 20924 19582 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19576 20896 19809 20924
rect 19576 20884 19582 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 30650 20884 30656 20936
rect 30708 20884 30714 20936
rect 30742 20884 30748 20936
rect 30800 20924 30806 20936
rect 32324 20933 32352 20964
rect 34790 20952 34796 20964
rect 34848 20952 34854 21004
rect 37826 20952 37832 21004
rect 37884 20992 37890 21004
rect 38381 20995 38439 21001
rect 38381 20992 38393 20995
rect 37884 20964 38393 20992
rect 37884 20952 37890 20964
rect 38381 20961 38393 20964
rect 38427 20961 38439 20995
rect 38381 20955 38439 20961
rect 31665 20927 31723 20933
rect 31665 20924 31677 20927
rect 30800 20896 31677 20924
rect 30800 20884 30806 20896
rect 31665 20893 31677 20896
rect 31711 20893 31723 20927
rect 31665 20887 31723 20893
rect 32309 20927 32367 20933
rect 32309 20893 32321 20927
rect 32355 20893 32367 20927
rect 32309 20887 32367 20893
rect 34698 20884 34704 20936
rect 34756 20924 34762 20936
rect 36817 20927 36875 20933
rect 36817 20924 36829 20927
rect 34756 20896 36829 20924
rect 34756 20884 34762 20896
rect 36817 20893 36829 20896
rect 36863 20893 36875 20927
rect 36817 20887 36875 20893
rect 38197 20927 38255 20933
rect 38197 20893 38209 20927
rect 38243 20924 38255 20927
rect 38286 20924 38292 20936
rect 38243 20896 38292 20924
rect 38243 20893 38255 20896
rect 38197 20887 38255 20893
rect 38286 20884 38292 20896
rect 38344 20884 38350 20936
rect 43806 20884 43812 20936
rect 43864 20884 43870 20936
rect 47026 20884 47032 20936
rect 47084 20924 47090 20936
rect 47949 20927 48007 20933
rect 47949 20924 47961 20927
rect 47084 20896 47961 20924
rect 47084 20884 47090 20896
rect 47949 20893 47961 20896
rect 47995 20893 48007 20927
rect 47949 20887 48007 20893
rect 43993 20859 44051 20865
rect 43993 20825 44005 20859
rect 44039 20856 44051 20859
rect 45186 20856 45192 20868
rect 44039 20828 45192 20856
rect 44039 20825 44051 20828
rect 43993 20819 44051 20825
rect 45186 20816 45192 20828
rect 45244 20816 45250 20868
rect 49142 20816 49148 20868
rect 49200 20816 49206 20868
rect 2866 20748 2872 20800
rect 2924 20788 2930 20800
rect 4249 20791 4307 20797
rect 4249 20788 4261 20791
rect 2924 20760 4261 20788
rect 2924 20748 2930 20760
rect 4249 20757 4261 20760
rect 4295 20757 4307 20791
rect 4249 20751 4307 20757
rect 19886 20748 19892 20800
rect 19944 20748 19950 20800
rect 30282 20748 30288 20800
rect 30340 20748 30346 20800
rect 30745 20791 30803 20797
rect 30745 20757 30757 20791
rect 30791 20788 30803 20791
rect 31386 20788 31392 20800
rect 30791 20760 31392 20788
rect 30791 20757 30803 20760
rect 30745 20751 30803 20757
rect 31386 20748 31392 20760
rect 31444 20748 31450 20800
rect 32122 20748 32128 20800
rect 32180 20748 32186 20800
rect 36446 20748 36452 20800
rect 36504 20788 36510 20800
rect 37829 20791 37887 20797
rect 37829 20788 37841 20791
rect 36504 20760 37841 20788
rect 36504 20748 36510 20760
rect 37829 20757 37841 20760
rect 37875 20757 37887 20791
rect 37829 20751 37887 20757
rect 38289 20791 38347 20797
rect 38289 20757 38301 20791
rect 38335 20788 38347 20791
rect 38378 20788 38384 20800
rect 38335 20760 38384 20788
rect 38335 20757 38347 20760
rect 38289 20751 38347 20757
rect 38378 20748 38384 20760
rect 38436 20748 38442 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 21174 20544 21180 20596
rect 21232 20544 21238 20596
rect 24857 20587 24915 20593
rect 24857 20553 24869 20587
rect 24903 20584 24915 20587
rect 25130 20584 25136 20596
rect 24903 20556 25136 20584
rect 24903 20553 24915 20556
rect 24857 20547 24915 20553
rect 25130 20544 25136 20556
rect 25188 20544 25194 20596
rect 26142 20544 26148 20596
rect 26200 20584 26206 20596
rect 26237 20587 26295 20593
rect 26237 20584 26249 20587
rect 26200 20556 26249 20584
rect 26200 20544 26206 20556
rect 26237 20553 26249 20556
rect 26283 20553 26295 20587
rect 26237 20547 26295 20553
rect 30009 20587 30067 20593
rect 30009 20553 30021 20587
rect 30055 20553 30067 20587
rect 30009 20547 30067 20553
rect 23290 20476 23296 20528
rect 23348 20516 23354 20528
rect 23385 20519 23443 20525
rect 23385 20516 23397 20519
rect 23348 20488 23397 20516
rect 23348 20476 23354 20488
rect 23385 20485 23397 20488
rect 23431 20485 23443 20519
rect 23385 20479 23443 20485
rect 23474 20476 23480 20528
rect 23532 20516 23538 20528
rect 23532 20488 23874 20516
rect 23532 20476 23538 20488
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 2774 20448 2780 20460
rect 1811 20420 2780 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 2774 20408 2780 20420
rect 2832 20408 2838 20460
rect 20806 20408 20812 20460
rect 20864 20448 20870 20460
rect 21085 20451 21143 20457
rect 21085 20448 21097 20451
rect 20864 20420 21097 20448
rect 20864 20408 20870 20420
rect 21085 20417 21097 20420
rect 21131 20448 21143 20451
rect 22370 20448 22376 20460
rect 21131 20420 22376 20448
rect 21131 20417 21143 20420
rect 21085 20411 21143 20417
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 22462 20408 22468 20460
rect 22520 20448 22526 20460
rect 23109 20451 23167 20457
rect 23109 20448 23121 20451
rect 22520 20420 23121 20448
rect 22520 20408 22526 20420
rect 23109 20417 23121 20420
rect 23155 20417 23167 20451
rect 23109 20411 23167 20417
rect 26142 20408 26148 20460
rect 26200 20408 26206 20460
rect 30024 20448 30052 20547
rect 30466 20544 30472 20596
rect 30524 20544 30530 20596
rect 32858 20544 32864 20596
rect 32916 20544 32922 20596
rect 30377 20519 30435 20525
rect 30377 20485 30389 20519
rect 30423 20516 30435 20519
rect 30742 20516 30748 20528
rect 30423 20488 30748 20516
rect 30423 20485 30435 20488
rect 30377 20479 30435 20485
rect 30742 20476 30748 20488
rect 30800 20476 30806 20528
rect 32769 20519 32827 20525
rect 32769 20516 32781 20519
rect 31726 20488 32781 20516
rect 31726 20448 31754 20488
rect 32769 20485 32781 20488
rect 32815 20485 32827 20519
rect 32769 20479 32827 20485
rect 30024 20420 31754 20448
rect 36906 20408 36912 20460
rect 36964 20408 36970 20460
rect 47854 20408 47860 20460
rect 47912 20448 47918 20460
rect 47949 20451 48007 20457
rect 47949 20448 47961 20451
rect 47912 20420 47961 20448
rect 47912 20408 47918 20420
rect 47949 20417 47961 20420
rect 47995 20417 48007 20451
rect 47949 20411 48007 20417
rect 1302 20340 1308 20392
rect 1360 20380 1366 20392
rect 2041 20383 2099 20389
rect 2041 20380 2053 20383
rect 1360 20352 2053 20380
rect 1360 20340 1366 20352
rect 2041 20349 2053 20352
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20380 21419 20383
rect 21910 20380 21916 20392
rect 21407 20352 21916 20380
rect 21407 20349 21419 20352
rect 21361 20343 21419 20349
rect 21910 20340 21916 20352
rect 21968 20340 21974 20392
rect 25498 20340 25504 20392
rect 25556 20380 25562 20392
rect 26421 20383 26479 20389
rect 26421 20380 26433 20383
rect 25556 20352 26433 20380
rect 25556 20340 25562 20352
rect 26421 20349 26433 20352
rect 26467 20380 26479 20383
rect 26602 20380 26608 20392
rect 26467 20352 26608 20380
rect 26467 20349 26479 20352
rect 26421 20343 26479 20349
rect 26602 20340 26608 20352
rect 26660 20340 26666 20392
rect 30653 20383 30711 20389
rect 30653 20349 30665 20383
rect 30699 20380 30711 20383
rect 32214 20380 32220 20392
rect 30699 20352 32220 20380
rect 30699 20349 30711 20352
rect 30653 20343 30711 20349
rect 32214 20340 32220 20352
rect 32272 20340 32278 20392
rect 33045 20383 33103 20389
rect 33045 20349 33057 20383
rect 33091 20380 33103 20383
rect 34238 20380 34244 20392
rect 33091 20352 34244 20380
rect 33091 20349 33103 20352
rect 33045 20343 33103 20349
rect 34238 20340 34244 20352
rect 34296 20340 34302 20392
rect 49142 20340 49148 20392
rect 49200 20340 49206 20392
rect 18598 20272 18604 20324
rect 18656 20312 18662 20324
rect 18656 20284 22094 20312
rect 18656 20272 18662 20284
rect 20717 20247 20775 20253
rect 20717 20213 20729 20247
rect 20763 20244 20775 20247
rect 21174 20244 21180 20256
rect 20763 20216 21180 20244
rect 20763 20213 20775 20216
rect 20717 20207 20775 20213
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 22066 20244 22094 20284
rect 27154 20272 27160 20324
rect 27212 20312 27218 20324
rect 34974 20312 34980 20324
rect 27212 20284 34980 20312
rect 27212 20272 27218 20284
rect 34974 20272 34980 20284
rect 35032 20312 35038 20324
rect 37182 20312 37188 20324
rect 35032 20284 37188 20312
rect 35032 20272 35038 20284
rect 37182 20272 37188 20284
rect 37240 20272 37246 20324
rect 24578 20244 24584 20256
rect 22066 20216 24584 20244
rect 24578 20204 24584 20216
rect 24636 20204 24642 20256
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 25777 20247 25835 20253
rect 25777 20244 25789 20247
rect 24912 20216 25789 20244
rect 24912 20204 24918 20216
rect 25777 20213 25789 20216
rect 25823 20213 25835 20247
rect 25777 20207 25835 20213
rect 32401 20247 32459 20253
rect 32401 20213 32413 20247
rect 32447 20244 32459 20247
rect 32582 20244 32588 20256
rect 32447 20216 32588 20244
rect 32447 20213 32459 20216
rect 32401 20207 32459 20213
rect 32582 20204 32588 20216
rect 32640 20204 32646 20256
rect 36725 20247 36783 20253
rect 36725 20213 36737 20247
rect 36771 20244 36783 20247
rect 44450 20244 44456 20256
rect 36771 20216 44456 20244
rect 36771 20213 36783 20216
rect 36725 20207 36783 20213
rect 44450 20204 44456 20216
rect 44508 20204 44514 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 10962 20000 10968 20052
rect 11020 20040 11026 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 11020 20012 14289 20040
rect 11020 20000 11026 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 18141 20043 18199 20049
rect 18141 20009 18153 20043
rect 18187 20040 18199 20043
rect 19978 20040 19984 20052
rect 18187 20012 19984 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 20530 20000 20536 20052
rect 20588 20040 20594 20052
rect 22084 20043 22142 20049
rect 22084 20040 22096 20043
rect 20588 20012 22096 20040
rect 20588 20000 20594 20012
rect 22084 20009 22096 20012
rect 22130 20040 22142 20043
rect 22130 20012 24900 20040
rect 22130 20009 22142 20012
rect 22084 20003 22142 20009
rect 24872 19972 24900 20012
rect 24946 20000 24952 20052
rect 25004 20040 25010 20052
rect 25225 20043 25283 20049
rect 25225 20040 25237 20043
rect 25004 20012 25237 20040
rect 25004 20000 25010 20012
rect 25225 20009 25237 20012
rect 25271 20009 25283 20043
rect 25225 20003 25283 20009
rect 26786 20000 26792 20052
rect 26844 20000 26850 20052
rect 31754 20000 31760 20052
rect 31812 20040 31818 20052
rect 35621 20043 35679 20049
rect 35621 20040 35633 20043
rect 31812 20012 35633 20040
rect 31812 20000 31818 20012
rect 35621 20009 35633 20012
rect 35667 20009 35679 20043
rect 35621 20003 35679 20009
rect 25498 19972 25504 19984
rect 24872 19944 25504 19972
rect 25498 19932 25504 19944
rect 25556 19932 25562 19984
rect 27062 19932 27068 19984
rect 27120 19972 27126 19984
rect 44910 19972 44916 19984
rect 27120 19944 44916 19972
rect 27120 19932 27126 19944
rect 44910 19932 44916 19944
rect 44968 19932 44974 19984
rect 18598 19864 18604 19916
rect 18656 19864 18662 19916
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 19426 19904 19432 19916
rect 18831 19876 19432 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 21821 19907 21879 19913
rect 21821 19904 21833 19907
rect 19668 19876 21833 19904
rect 19668 19864 19674 19876
rect 21821 19873 21833 19876
rect 21867 19904 21879 19907
rect 22462 19904 22468 19916
rect 21867 19876 22468 19904
rect 21867 19873 21879 19876
rect 21821 19867 21879 19873
rect 22462 19864 22468 19876
rect 22520 19864 22526 19916
rect 25130 19864 25136 19916
rect 25188 19904 25194 19916
rect 25777 19907 25835 19913
rect 25777 19904 25789 19907
rect 25188 19876 25789 19904
rect 25188 19864 25194 19876
rect 25777 19873 25789 19876
rect 25823 19873 25835 19907
rect 27433 19907 27491 19913
rect 25777 19867 25835 19873
rect 25884 19876 27292 19904
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19836 14519 19839
rect 15654 19836 15660 19848
rect 14507 19808 15660 19836
rect 14507 19805 14519 19808
rect 14461 19799 14519 19805
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 17310 19796 17316 19848
rect 17368 19836 17374 19848
rect 17678 19836 17684 19848
rect 17368 19808 17684 19836
rect 17368 19796 17374 19808
rect 17678 19796 17684 19808
rect 17736 19836 17742 19848
rect 18509 19839 18567 19845
rect 18509 19836 18521 19839
rect 17736 19808 18521 19836
rect 17736 19796 17742 19808
rect 18509 19805 18521 19808
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 19444 19768 19472 19864
rect 23934 19796 23940 19848
rect 23992 19836 23998 19848
rect 25884 19836 25912 19876
rect 23992 19808 25912 19836
rect 23992 19796 23998 19808
rect 27154 19796 27160 19848
rect 27212 19796 27218 19848
rect 27264 19836 27292 19876
rect 27433 19873 27445 19907
rect 27479 19904 27491 19907
rect 27522 19904 27528 19916
rect 27479 19876 27528 19904
rect 27479 19873 27491 19876
rect 27433 19867 27491 19873
rect 27522 19864 27528 19876
rect 27580 19864 27586 19916
rect 32674 19864 32680 19916
rect 32732 19904 32738 19916
rect 35342 19904 35348 19916
rect 32732 19876 35348 19904
rect 32732 19864 32738 19876
rect 35342 19864 35348 19876
rect 35400 19864 35406 19916
rect 27798 19836 27804 19848
rect 27264 19808 27804 19836
rect 27798 19796 27804 19808
rect 27856 19796 27862 19848
rect 31938 19796 31944 19848
rect 31996 19836 32002 19848
rect 32214 19836 32220 19848
rect 31996 19808 32220 19836
rect 31996 19796 32002 19808
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 32306 19796 32312 19848
rect 32364 19796 32370 19848
rect 33137 19839 33195 19845
rect 33137 19805 33149 19839
rect 33183 19836 33195 19839
rect 33318 19836 33324 19848
rect 33183 19808 33324 19836
rect 33183 19805 33195 19808
rect 33137 19799 33195 19805
rect 33318 19796 33324 19808
rect 33376 19796 33382 19848
rect 33873 19839 33931 19845
rect 33873 19805 33885 19839
rect 33919 19836 33931 19839
rect 33962 19836 33968 19848
rect 33919 19808 33968 19836
rect 33919 19805 33931 19808
rect 33873 19799 33931 19805
rect 33962 19796 33968 19808
rect 34020 19796 34026 19848
rect 34977 19839 35035 19845
rect 34977 19805 34989 19839
rect 35023 19836 35035 19839
rect 35434 19836 35440 19848
rect 35023 19808 35440 19836
rect 35023 19805 35035 19808
rect 34977 19799 35035 19805
rect 35434 19796 35440 19808
rect 35492 19796 35498 19848
rect 35805 19839 35863 19845
rect 35805 19805 35817 19839
rect 35851 19836 35863 19839
rect 36354 19836 36360 19848
rect 35851 19808 36360 19836
rect 35851 19805 35863 19808
rect 35805 19799 35863 19805
rect 36354 19796 36360 19808
rect 36412 19796 36418 19848
rect 44082 19796 44088 19848
rect 44140 19836 44146 19848
rect 44177 19839 44235 19845
rect 44177 19836 44189 19839
rect 44140 19808 44189 19836
rect 44140 19796 44146 19808
rect 44177 19805 44189 19808
rect 44223 19805 44235 19839
rect 44177 19799 44235 19805
rect 19794 19768 19800 19780
rect 19444 19740 19800 19768
rect 19794 19728 19800 19740
rect 19852 19728 19858 19780
rect 19889 19771 19947 19777
rect 19889 19737 19901 19771
rect 19935 19737 19947 19771
rect 19889 19731 19947 19737
rect 19904 19700 19932 19731
rect 20898 19728 20904 19780
rect 20956 19728 20962 19780
rect 23474 19768 23480 19780
rect 23322 19740 23480 19768
rect 23474 19728 23480 19740
rect 23532 19768 23538 19780
rect 24210 19768 24216 19780
rect 23532 19740 24216 19768
rect 23532 19728 23538 19740
rect 24210 19728 24216 19740
rect 24268 19728 24274 19780
rect 25593 19771 25651 19777
rect 25593 19737 25605 19771
rect 25639 19768 25651 19771
rect 27338 19768 27344 19780
rect 25639 19740 27344 19768
rect 25639 19737 25651 19740
rect 25593 19731 25651 19737
rect 27338 19728 27344 19740
rect 27396 19728 27402 19780
rect 34057 19771 34115 19777
rect 34057 19737 34069 19771
rect 34103 19768 34115 19771
rect 34330 19768 34336 19780
rect 34103 19740 34336 19768
rect 34103 19737 34115 19740
rect 34057 19731 34115 19737
rect 34330 19728 34336 19740
rect 34388 19728 34394 19780
rect 44361 19771 44419 19777
rect 44361 19737 44373 19771
rect 44407 19768 44419 19771
rect 46198 19768 46204 19780
rect 44407 19740 46204 19768
rect 44407 19737 44419 19740
rect 44361 19731 44419 19737
rect 46198 19728 46204 19740
rect 46256 19728 46262 19780
rect 21266 19700 21272 19712
rect 19904 19672 21272 19700
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 21361 19703 21419 19709
rect 21361 19669 21373 19703
rect 21407 19700 21419 19703
rect 21450 19700 21456 19712
rect 21407 19672 21456 19700
rect 21407 19669 21419 19672
rect 21361 19663 21419 19669
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 23566 19660 23572 19712
rect 23624 19660 23630 19712
rect 25685 19703 25743 19709
rect 25685 19669 25697 19703
rect 25731 19700 25743 19703
rect 26510 19700 26516 19712
rect 25731 19672 26516 19700
rect 25731 19669 25743 19672
rect 25685 19663 25743 19669
rect 26510 19660 26516 19672
rect 26568 19660 26574 19712
rect 27246 19660 27252 19712
rect 27304 19660 27310 19712
rect 31938 19660 31944 19712
rect 31996 19700 32002 19712
rect 32401 19703 32459 19709
rect 32401 19700 32413 19703
rect 31996 19672 32413 19700
rect 31996 19660 32002 19672
rect 32401 19669 32413 19672
rect 32447 19669 32459 19703
rect 32401 19663 32459 19669
rect 33229 19703 33287 19709
rect 33229 19669 33241 19703
rect 33275 19700 33287 19703
rect 33318 19700 33324 19712
rect 33275 19672 33324 19700
rect 33275 19669 33287 19672
rect 33229 19663 33287 19669
rect 33318 19660 33324 19672
rect 33376 19660 33382 19712
rect 34974 19660 34980 19712
rect 35032 19700 35038 19712
rect 35069 19703 35127 19709
rect 35069 19700 35081 19703
rect 35032 19672 35081 19700
rect 35032 19660 35038 19672
rect 35069 19669 35081 19672
rect 35115 19669 35127 19703
rect 35069 19663 35127 19669
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 16022 19456 16028 19508
rect 16080 19496 16086 19508
rect 19521 19499 19579 19505
rect 19521 19496 19533 19499
rect 16080 19468 19533 19496
rect 16080 19456 16086 19468
rect 19521 19465 19533 19468
rect 19567 19465 19579 19499
rect 19521 19459 19579 19465
rect 19889 19499 19947 19505
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 19935 19468 20729 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 20717 19465 20729 19468
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 21085 19499 21143 19505
rect 21085 19465 21097 19499
rect 21131 19496 21143 19499
rect 21358 19496 21364 19508
rect 21131 19468 21364 19496
rect 21131 19465 21143 19468
rect 21085 19459 21143 19465
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 38470 19496 38476 19508
rect 22020 19468 28304 19496
rect 20070 19388 20076 19440
rect 20128 19428 20134 19440
rect 21177 19431 21235 19437
rect 21177 19428 21189 19431
rect 20128 19400 21189 19428
rect 20128 19388 20134 19400
rect 21177 19397 21189 19400
rect 21223 19397 21235 19431
rect 21177 19391 21235 19397
rect 21726 19388 21732 19440
rect 21784 19428 21790 19440
rect 22020 19437 22048 19468
rect 22005 19431 22063 19437
rect 22005 19428 22017 19431
rect 21784 19400 22017 19428
rect 21784 19388 21790 19400
rect 22005 19397 22017 19400
rect 22051 19397 22063 19431
rect 22005 19391 22063 19397
rect 22462 19388 22468 19440
rect 22520 19428 22526 19440
rect 22741 19431 22799 19437
rect 22741 19428 22753 19431
rect 22520 19400 22753 19428
rect 22520 19388 22526 19400
rect 22741 19397 22753 19400
rect 22787 19397 22799 19431
rect 22741 19391 22799 19397
rect 23290 19388 23296 19440
rect 23348 19428 23354 19440
rect 23348 19400 23520 19428
rect 23348 19388 23354 19400
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19360 20039 19363
rect 20990 19360 20996 19372
rect 20027 19332 20996 19360
rect 20027 19329 20039 19332
rect 19981 19323 20039 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 21450 19360 21456 19372
rect 21192 19332 21456 19360
rect 20165 19295 20223 19301
rect 20165 19261 20177 19295
rect 20211 19292 20223 19295
rect 21192 19292 21220 19332
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 22278 19320 22284 19372
rect 22336 19360 22342 19372
rect 22336 19332 23428 19360
rect 22336 19320 22342 19332
rect 20211 19264 21220 19292
rect 20211 19261 20223 19264
rect 20165 19255 20223 19261
rect 21266 19252 21272 19304
rect 21324 19252 21330 19304
rect 21542 19252 21548 19304
rect 21600 19292 21606 19304
rect 23290 19292 23296 19304
rect 21600 19264 23296 19292
rect 21600 19252 21606 19264
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 21284 19156 21312 19252
rect 23400 19233 23428 19332
rect 23492 19292 23520 19400
rect 23658 19388 23664 19440
rect 23716 19428 23722 19440
rect 23845 19431 23903 19437
rect 23845 19428 23857 19431
rect 23716 19400 23857 19428
rect 23716 19388 23722 19400
rect 23845 19397 23857 19400
rect 23891 19428 23903 19431
rect 24118 19428 24124 19440
rect 23891 19400 24124 19428
rect 23891 19397 23903 19400
rect 23845 19391 23903 19397
rect 24118 19388 24124 19400
rect 24176 19388 24182 19440
rect 24210 19388 24216 19440
rect 24268 19428 24274 19440
rect 28276 19437 28304 19468
rect 33796 19468 36216 19496
rect 28261 19431 28319 19437
rect 24268 19400 25346 19428
rect 24268 19388 24274 19400
rect 28261 19397 28273 19431
rect 28307 19428 28319 19431
rect 28350 19428 28356 19440
rect 28307 19400 28356 19428
rect 28307 19397 28319 19400
rect 28261 19391 28319 19397
rect 28350 19388 28356 19400
rect 28408 19428 28414 19440
rect 29641 19431 29699 19437
rect 29641 19428 29653 19431
rect 28408 19400 29653 19428
rect 28408 19388 28414 19400
rect 29641 19397 29653 19400
rect 29687 19397 29699 19431
rect 33796 19428 33824 19468
rect 36078 19428 36084 19440
rect 29641 19391 29699 19397
rect 33704 19400 33824 19428
rect 35190 19400 36084 19428
rect 23753 19363 23811 19369
rect 23753 19329 23765 19363
rect 23799 19360 23811 19363
rect 23934 19360 23940 19372
rect 23799 19332 23940 19360
rect 23799 19329 23811 19332
rect 23753 19323 23811 19329
rect 23934 19320 23940 19332
rect 23992 19320 23998 19372
rect 24394 19320 24400 19372
rect 24452 19360 24458 19372
rect 24570 19363 24628 19369
rect 24570 19360 24582 19363
rect 24452 19332 24582 19360
rect 24452 19320 24458 19332
rect 24570 19329 24582 19332
rect 24616 19329 24628 19363
rect 24570 19323 24628 19329
rect 26602 19320 26608 19372
rect 26660 19360 26666 19372
rect 26786 19360 26792 19372
rect 26660 19332 26792 19360
rect 26660 19320 26666 19332
rect 26786 19320 26792 19332
rect 26844 19320 26850 19372
rect 28442 19320 28448 19372
rect 28500 19360 28506 19372
rect 29730 19360 29736 19372
rect 28500 19332 29736 19360
rect 28500 19320 28506 19332
rect 29730 19320 29736 19332
rect 29788 19320 29794 19372
rect 33704 19369 33732 19400
rect 36078 19388 36084 19400
rect 36136 19388 36142 19440
rect 33689 19363 33747 19369
rect 33689 19329 33701 19363
rect 33735 19329 33747 19363
rect 33689 19323 33747 19329
rect 35342 19320 35348 19372
rect 35400 19360 35406 19372
rect 35400 19332 35480 19360
rect 35400 19320 35406 19332
rect 24029 19295 24087 19301
rect 24029 19292 24041 19295
rect 23492 19264 24041 19292
rect 24029 19261 24041 19264
rect 24075 19292 24087 19295
rect 24857 19295 24915 19301
rect 24857 19292 24869 19295
rect 24075 19264 24532 19292
rect 24075 19261 24087 19264
rect 24029 19255 24087 19261
rect 23385 19227 23443 19233
rect 23385 19193 23397 19227
rect 23431 19193 23443 19227
rect 23385 19187 23443 19193
rect 23566 19156 23572 19168
rect 21284 19128 23572 19156
rect 23566 19116 23572 19128
rect 23624 19116 23630 19168
rect 24504 19156 24532 19264
rect 24688 19264 24869 19292
rect 24578 19184 24584 19236
rect 24636 19224 24642 19236
rect 24688 19224 24716 19264
rect 24857 19261 24869 19264
rect 24903 19292 24915 19295
rect 27890 19292 27896 19304
rect 24903 19264 27896 19292
rect 24903 19261 24915 19264
rect 24857 19255 24915 19261
rect 27890 19252 27896 19264
rect 27948 19252 27954 19304
rect 28810 19252 28816 19304
rect 28868 19292 28874 19304
rect 28997 19295 29055 19301
rect 28997 19292 29009 19295
rect 28868 19264 29009 19292
rect 28868 19252 28874 19264
rect 28997 19261 29009 19264
rect 29043 19261 29055 19295
rect 28997 19255 29055 19261
rect 29822 19252 29828 19304
rect 29880 19292 29886 19304
rect 35452 19301 35480 19332
rect 30377 19295 30435 19301
rect 30377 19292 30389 19295
rect 29880 19264 30389 19292
rect 29880 19252 29886 19264
rect 30377 19261 30389 19264
rect 30423 19261 30435 19295
rect 30377 19255 30435 19261
rect 33965 19295 34023 19301
rect 33965 19261 33977 19295
rect 34011 19292 34023 19295
rect 35437 19295 35495 19301
rect 34011 19264 35388 19292
rect 34011 19261 34023 19264
rect 33965 19255 34023 19261
rect 24636 19196 24716 19224
rect 35360 19224 35388 19264
rect 35437 19261 35449 19295
rect 35483 19261 35495 19295
rect 36188 19292 36216 19468
rect 37476 19468 38476 19496
rect 37274 19320 37280 19372
rect 37332 19360 37338 19372
rect 37476 19369 37504 19468
rect 38470 19456 38476 19468
rect 38528 19456 38534 19508
rect 38562 19456 38568 19508
rect 38620 19496 38626 19508
rect 39209 19499 39267 19505
rect 39209 19496 39221 19499
rect 38620 19468 39221 19496
rect 38620 19456 38626 19468
rect 39209 19465 39221 19468
rect 39255 19465 39267 19499
rect 39209 19459 39267 19465
rect 38746 19388 38752 19440
rect 38804 19388 38810 19440
rect 37461 19363 37519 19369
rect 37461 19360 37473 19363
rect 37332 19332 37473 19360
rect 37332 19320 37338 19332
rect 37461 19329 37473 19332
rect 37507 19329 37519 19363
rect 37461 19323 37519 19329
rect 45462 19320 45468 19372
rect 45520 19360 45526 19372
rect 47949 19363 48007 19369
rect 47949 19360 47961 19363
rect 45520 19332 47961 19360
rect 45520 19320 45526 19332
rect 47949 19329 47961 19332
rect 47995 19329 48007 19363
rect 47949 19323 48007 19329
rect 49142 19320 49148 19372
rect 49200 19320 49206 19372
rect 37292 19292 37320 19320
rect 37737 19295 37795 19301
rect 37737 19292 37749 19295
rect 36188 19264 37320 19292
rect 37476 19264 37749 19292
rect 35437 19255 35495 19261
rect 37476 19236 37504 19264
rect 37737 19261 37749 19264
rect 37783 19261 37795 19295
rect 37737 19255 37795 19261
rect 36630 19224 36636 19236
rect 35360 19196 36636 19224
rect 24636 19184 24642 19196
rect 36630 19184 36636 19196
rect 36688 19184 36694 19236
rect 37458 19184 37464 19236
rect 37516 19184 37522 19236
rect 26326 19156 26332 19168
rect 24504 19128 26332 19156
rect 26326 19116 26332 19128
rect 26384 19156 26390 19168
rect 27430 19156 27436 19168
rect 26384 19128 27436 19156
rect 26384 19116 26390 19128
rect 27430 19116 27436 19128
rect 27488 19116 27494 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18952 18199 18955
rect 18187 18924 19840 18952
rect 18187 18921 18199 18924
rect 18141 18915 18199 18921
rect 9766 18844 9772 18896
rect 9824 18884 9830 18896
rect 18325 18887 18383 18893
rect 18325 18884 18337 18887
rect 9824 18856 18337 18884
rect 9824 18844 9830 18856
rect 18325 18853 18337 18856
rect 18371 18853 18383 18887
rect 19812 18884 19840 18924
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 20533 18955 20591 18961
rect 20533 18952 20545 18955
rect 19944 18924 20545 18952
rect 19944 18912 19950 18924
rect 20533 18921 20545 18924
rect 20579 18921 20591 18955
rect 20533 18915 20591 18921
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 23293 18955 23351 18961
rect 23293 18952 23305 18955
rect 21048 18924 23305 18952
rect 21048 18912 21054 18924
rect 23293 18921 23305 18924
rect 23339 18921 23351 18955
rect 23293 18915 23351 18921
rect 23382 18912 23388 18964
rect 23440 18952 23446 18964
rect 24581 18955 24639 18961
rect 24581 18952 24593 18955
rect 23440 18924 24593 18952
rect 23440 18912 23446 18924
rect 24581 18921 24593 18924
rect 24627 18921 24639 18955
rect 24581 18915 24639 18921
rect 26142 18912 26148 18964
rect 26200 18952 26206 18964
rect 27157 18955 27215 18961
rect 27157 18952 27169 18955
rect 26200 18924 27169 18952
rect 26200 18912 26206 18924
rect 27157 18921 27169 18924
rect 27203 18921 27215 18955
rect 34974 18952 34980 18964
rect 27157 18915 27215 18921
rect 30944 18924 34980 18952
rect 24670 18884 24676 18896
rect 19812 18856 24676 18884
rect 18325 18847 18383 18853
rect 24670 18844 24676 18856
rect 24728 18844 24734 18896
rect 21177 18819 21235 18825
rect 21177 18785 21189 18819
rect 21223 18816 21235 18819
rect 22370 18816 22376 18828
rect 21223 18788 22376 18816
rect 21223 18785 21235 18788
rect 21177 18779 21235 18785
rect 22370 18776 22376 18788
rect 22428 18816 22434 18828
rect 22830 18816 22836 18828
rect 22428 18788 22836 18816
rect 22428 18776 22434 18788
rect 22830 18776 22836 18788
rect 22888 18776 22894 18828
rect 23566 18776 23572 18828
rect 23624 18816 23630 18828
rect 23845 18819 23903 18825
rect 23845 18816 23857 18819
rect 23624 18788 23857 18816
rect 23624 18776 23630 18788
rect 23845 18785 23857 18788
rect 23891 18785 23903 18819
rect 23845 18779 23903 18785
rect 24762 18776 24768 18828
rect 24820 18816 24826 18828
rect 25133 18819 25191 18825
rect 25133 18816 25145 18819
rect 24820 18788 25145 18816
rect 24820 18776 24826 18788
rect 25133 18785 25145 18788
rect 25179 18785 25191 18819
rect 25133 18779 25191 18785
rect 25590 18776 25596 18828
rect 25648 18816 25654 18828
rect 25648 18788 26372 18816
rect 25648 18776 25654 18788
rect 4617 18751 4675 18757
rect 4617 18717 4629 18751
rect 4663 18748 4675 18751
rect 9306 18748 9312 18760
rect 4663 18720 9312 18748
rect 4663 18717 4675 18720
rect 4617 18711 4675 18717
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 12676 18720 17877 18748
rect 12676 18708 12682 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 21726 18708 21732 18760
rect 21784 18708 21790 18760
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18748 23719 18751
rect 24854 18748 24860 18760
rect 23707 18720 24860 18748
rect 23707 18717 23719 18720
rect 23661 18711 23719 18717
rect 24854 18708 24860 18720
rect 24912 18708 24918 18760
rect 26234 18748 26240 18760
rect 24964 18720 26240 18748
rect 20901 18683 20959 18689
rect 20901 18649 20913 18683
rect 20947 18680 20959 18683
rect 22462 18680 22468 18692
rect 20947 18652 22468 18680
rect 20947 18649 20959 18652
rect 20901 18643 20959 18649
rect 22462 18640 22468 18652
rect 22520 18640 22526 18692
rect 22554 18640 22560 18692
rect 22612 18640 22618 18692
rect 23753 18683 23811 18689
rect 23753 18649 23765 18683
rect 23799 18680 23811 18683
rect 24964 18680 24992 18720
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 26344 18748 26372 18788
rect 26418 18776 26424 18828
rect 26476 18776 26482 18828
rect 26602 18776 26608 18828
rect 26660 18776 26666 18828
rect 27801 18819 27859 18825
rect 27801 18785 27813 18819
rect 27847 18816 27859 18819
rect 27890 18816 27896 18828
rect 27847 18788 27896 18816
rect 27847 18785 27859 18788
rect 27801 18779 27859 18785
rect 27890 18776 27896 18788
rect 27948 18816 27954 18828
rect 28626 18816 28632 18828
rect 27948 18788 28632 18816
rect 27948 18776 27954 18788
rect 28626 18776 28632 18788
rect 28684 18776 28690 18828
rect 28718 18776 28724 18828
rect 28776 18816 28782 18828
rect 28813 18819 28871 18825
rect 28813 18816 28825 18819
rect 28776 18788 28825 18816
rect 28776 18776 28782 18788
rect 28813 18785 28825 18788
rect 28859 18785 28871 18819
rect 28813 18779 28871 18785
rect 28902 18776 28908 18828
rect 28960 18776 28966 18828
rect 27525 18751 27583 18757
rect 26344 18720 27292 18748
rect 23799 18652 24992 18680
rect 25041 18683 25099 18689
rect 23799 18649 23811 18652
rect 23753 18643 23811 18649
rect 25041 18649 25053 18683
rect 25087 18680 25099 18683
rect 27154 18680 27160 18692
rect 25087 18652 27160 18680
rect 25087 18649 25099 18652
rect 25041 18643 25099 18649
rect 27154 18640 27160 18652
rect 27212 18640 27218 18692
rect 27264 18680 27292 18720
rect 27525 18717 27537 18751
rect 27571 18748 27583 18751
rect 27571 18720 28672 18748
rect 27571 18717 27583 18720
rect 27525 18711 27583 18717
rect 27264 18652 28396 18680
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 4709 18615 4767 18621
rect 4709 18612 4721 18615
rect 2832 18584 4721 18612
rect 2832 18572 2838 18584
rect 4709 18581 4721 18584
rect 4755 18581 4767 18615
rect 4709 18575 4767 18581
rect 20993 18615 21051 18621
rect 20993 18581 21005 18615
rect 21039 18612 21051 18615
rect 21358 18612 21364 18624
rect 21039 18584 21364 18612
rect 21039 18581 21051 18584
rect 20993 18575 21051 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 24946 18572 24952 18624
rect 25004 18572 25010 18624
rect 25958 18572 25964 18624
rect 26016 18572 26022 18624
rect 26326 18572 26332 18624
rect 26384 18572 26390 18624
rect 27246 18572 27252 18624
rect 27304 18612 27310 18624
rect 28368 18621 28396 18652
rect 27617 18615 27675 18621
rect 27617 18612 27629 18615
rect 27304 18584 27629 18612
rect 27304 18572 27310 18584
rect 27617 18581 27629 18584
rect 27663 18581 27675 18615
rect 27617 18575 27675 18581
rect 28353 18615 28411 18621
rect 28353 18581 28365 18615
rect 28399 18581 28411 18615
rect 28644 18612 28672 18720
rect 28721 18683 28779 18689
rect 28721 18649 28733 18683
rect 28767 18680 28779 18683
rect 30944 18680 30972 18924
rect 34974 18912 34980 18924
rect 35032 18912 35038 18964
rect 31021 18887 31079 18893
rect 31021 18853 31033 18887
rect 31067 18884 31079 18887
rect 32858 18884 32864 18896
rect 31067 18856 32864 18884
rect 31067 18853 31079 18856
rect 31021 18847 31079 18853
rect 32858 18844 32864 18856
rect 32916 18844 32922 18896
rect 31478 18776 31484 18828
rect 31536 18776 31542 18828
rect 31665 18819 31723 18825
rect 31665 18785 31677 18819
rect 31711 18816 31723 18819
rect 32490 18816 32496 18828
rect 31711 18788 32496 18816
rect 31711 18785 31723 18788
rect 31665 18779 31723 18785
rect 32490 18776 32496 18788
rect 32548 18776 32554 18828
rect 36909 18819 36967 18825
rect 36909 18785 36921 18819
rect 36955 18816 36967 18819
rect 37274 18816 37280 18828
rect 36955 18788 37280 18816
rect 36955 18785 36967 18788
rect 36909 18779 36967 18785
rect 37274 18776 37280 18788
rect 37332 18776 37338 18828
rect 31294 18708 31300 18760
rect 31352 18708 31358 18760
rect 34238 18708 34244 18760
rect 34296 18748 34302 18760
rect 36078 18748 36084 18760
rect 34296 18720 36084 18748
rect 34296 18708 34302 18720
rect 36078 18708 36084 18720
rect 36136 18708 36142 18760
rect 36170 18708 36176 18760
rect 36228 18748 36234 18760
rect 36265 18751 36323 18757
rect 36265 18748 36277 18751
rect 36228 18720 36277 18748
rect 36228 18708 36234 18720
rect 36265 18717 36277 18720
rect 36311 18717 36323 18751
rect 36265 18711 36323 18717
rect 44174 18708 44180 18760
rect 44232 18708 44238 18760
rect 44634 18708 44640 18760
rect 44692 18748 44698 18760
rect 47949 18751 48007 18757
rect 47949 18748 47961 18751
rect 44692 18720 47961 18748
rect 44692 18708 44698 18720
rect 47949 18717 47961 18720
rect 47995 18717 48007 18751
rect 47949 18711 48007 18717
rect 28767 18652 30972 18680
rect 31312 18680 31340 18708
rect 31389 18683 31447 18689
rect 31389 18680 31401 18683
rect 31312 18652 31401 18680
rect 28767 18649 28779 18652
rect 28721 18643 28779 18649
rect 31389 18649 31401 18652
rect 31435 18649 31447 18683
rect 31389 18643 31447 18649
rect 36449 18683 36507 18689
rect 36449 18649 36461 18683
rect 36495 18680 36507 18683
rect 36722 18680 36728 18692
rect 36495 18652 36728 18680
rect 36495 18649 36507 18652
rect 36449 18643 36507 18649
rect 36722 18640 36728 18652
rect 36780 18640 36786 18692
rect 37185 18683 37243 18689
rect 37185 18649 37197 18683
rect 37231 18649 37243 18683
rect 38746 18680 38752 18692
rect 38410 18652 38752 18680
rect 37185 18643 37243 18649
rect 34146 18612 34152 18624
rect 28644 18584 34152 18612
rect 28353 18575 28411 18581
rect 34146 18572 34152 18584
rect 34204 18612 34210 18624
rect 35158 18612 35164 18624
rect 34204 18584 35164 18612
rect 34204 18572 34210 18584
rect 35158 18572 35164 18584
rect 35216 18572 35222 18624
rect 37200 18612 37228 18643
rect 38746 18640 38752 18652
rect 38804 18640 38810 18692
rect 44361 18683 44419 18689
rect 44361 18649 44373 18683
rect 44407 18680 44419 18683
rect 47854 18680 47860 18692
rect 44407 18652 47860 18680
rect 44407 18649 44419 18652
rect 44361 18643 44419 18649
rect 47854 18640 47860 18652
rect 47912 18640 47918 18692
rect 49142 18640 49148 18692
rect 49200 18640 49206 18692
rect 37366 18612 37372 18624
rect 37200 18584 37372 18612
rect 37366 18572 37372 18584
rect 37424 18572 37430 18624
rect 37458 18572 37464 18624
rect 37516 18612 37522 18624
rect 38657 18615 38715 18621
rect 38657 18612 38669 18615
rect 37516 18584 38669 18612
rect 37516 18572 37522 18584
rect 38657 18581 38669 18584
rect 38703 18612 38715 18615
rect 39206 18612 39212 18624
rect 38703 18584 39212 18612
rect 38703 18581 38715 18584
rect 38657 18575 38715 18581
rect 39206 18572 39212 18584
rect 39264 18572 39270 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 19797 18411 19855 18417
rect 19797 18377 19809 18411
rect 19843 18408 19855 18411
rect 20717 18411 20775 18417
rect 20717 18408 20729 18411
rect 19843 18380 20729 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 20717 18377 20729 18380
rect 20763 18377 20775 18411
rect 20717 18371 20775 18377
rect 21174 18368 21180 18420
rect 21232 18368 21238 18420
rect 24302 18408 24308 18420
rect 23676 18380 24308 18408
rect 19889 18343 19947 18349
rect 19889 18309 19901 18343
rect 19935 18340 19947 18343
rect 21266 18340 21272 18352
rect 19935 18312 21272 18340
rect 19935 18309 19947 18312
rect 19889 18303 19947 18309
rect 21266 18300 21272 18312
rect 21324 18300 21330 18352
rect 21450 18300 21456 18352
rect 21508 18340 21514 18352
rect 23293 18343 23351 18349
rect 23293 18340 23305 18343
rect 21508 18312 23305 18340
rect 21508 18300 21514 18312
rect 23293 18309 23305 18312
rect 23339 18309 23351 18343
rect 23293 18303 23351 18309
rect 23566 18300 23572 18352
rect 23624 18340 23630 18352
rect 23676 18340 23704 18380
rect 24302 18368 24308 18380
rect 24360 18368 24366 18420
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 27341 18411 27399 18417
rect 27341 18408 27353 18411
rect 25004 18380 27353 18408
rect 25004 18368 25010 18380
rect 27341 18377 27353 18380
rect 27387 18377 27399 18411
rect 27341 18371 27399 18377
rect 27801 18411 27859 18417
rect 27801 18377 27813 18411
rect 27847 18408 27859 18411
rect 28442 18408 28448 18420
rect 27847 18380 28448 18408
rect 27847 18377 27859 18380
rect 27801 18371 27859 18377
rect 28442 18368 28448 18380
rect 28500 18368 28506 18420
rect 29825 18411 29883 18417
rect 29825 18377 29837 18411
rect 29871 18408 29883 18411
rect 33594 18408 33600 18420
rect 29871 18380 33600 18408
rect 29871 18377 29883 18380
rect 29825 18371 29883 18377
rect 33594 18368 33600 18380
rect 33652 18368 33658 18420
rect 34057 18411 34115 18417
rect 34057 18377 34069 18411
rect 34103 18408 34115 18411
rect 34790 18408 34796 18420
rect 34103 18380 34796 18408
rect 34103 18377 34115 18380
rect 34057 18371 34115 18377
rect 34790 18368 34796 18380
rect 34848 18368 34854 18420
rect 35066 18368 35072 18420
rect 35124 18408 35130 18420
rect 37829 18411 37887 18417
rect 37829 18408 37841 18411
rect 35124 18380 37841 18408
rect 35124 18368 35130 18380
rect 37829 18377 37841 18380
rect 37875 18377 37887 18411
rect 37829 18371 37887 18377
rect 37921 18411 37979 18417
rect 37921 18377 37933 18411
rect 37967 18408 37979 18411
rect 38654 18408 38660 18420
rect 37967 18380 38660 18408
rect 37967 18377 37979 18380
rect 37921 18371 37979 18377
rect 38654 18368 38660 18380
rect 38712 18368 38718 18420
rect 23624 18312 23782 18340
rect 23624 18300 23630 18312
rect 25038 18300 25044 18352
rect 25096 18300 25102 18352
rect 27246 18300 27252 18352
rect 27304 18340 27310 18352
rect 30193 18343 30251 18349
rect 30193 18340 30205 18343
rect 27304 18312 30205 18340
rect 27304 18300 27310 18312
rect 30193 18309 30205 18312
rect 30239 18309 30251 18343
rect 30193 18303 30251 18309
rect 30285 18343 30343 18349
rect 30285 18309 30297 18343
rect 30331 18340 30343 18343
rect 30834 18340 30840 18352
rect 30331 18312 30840 18340
rect 30331 18309 30343 18312
rect 30285 18303 30343 18309
rect 30834 18300 30840 18312
rect 30892 18300 30898 18352
rect 32490 18300 32496 18352
rect 32548 18340 32554 18352
rect 32585 18343 32643 18349
rect 32585 18340 32597 18343
rect 32548 18312 32597 18340
rect 32548 18300 32554 18312
rect 32585 18309 32597 18312
rect 32631 18309 32643 18343
rect 33870 18340 33876 18352
rect 33810 18312 33876 18340
rect 32585 18303 32643 18309
rect 33870 18300 33876 18312
rect 33928 18340 33934 18352
rect 34238 18340 34244 18352
rect 33928 18312 34244 18340
rect 33928 18300 33934 18312
rect 34238 18300 34244 18312
rect 34296 18300 34302 18352
rect 36078 18340 36084 18352
rect 36018 18312 36084 18340
rect 36078 18300 36084 18312
rect 36136 18340 36142 18352
rect 36538 18340 36544 18352
rect 36136 18312 36544 18340
rect 36136 18300 36142 18312
rect 36538 18300 36544 18312
rect 36596 18300 36602 18352
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2866 18272 2872 18284
rect 1811 18244 2872 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 2866 18232 2872 18244
rect 2924 18232 2930 18284
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18272 21143 18275
rect 22830 18272 22836 18284
rect 21131 18244 22836 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 27614 18232 27620 18284
rect 27672 18272 27678 18284
rect 27709 18275 27767 18281
rect 27709 18272 27721 18275
rect 27672 18244 27721 18272
rect 27672 18232 27678 18244
rect 27709 18241 27721 18244
rect 27755 18272 27767 18275
rect 31938 18272 31944 18284
rect 27755 18244 29040 18272
rect 27755 18241 27767 18244
rect 27709 18235 27767 18241
rect 1302 18164 1308 18216
rect 1360 18204 1366 18216
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 1360 18176 2053 18204
rect 1360 18164 1366 18176
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 20073 18207 20131 18213
rect 20073 18173 20085 18207
rect 20119 18204 20131 18207
rect 20990 18204 20996 18216
rect 20119 18176 20996 18204
rect 20119 18173 20131 18176
rect 20073 18167 20131 18173
rect 20990 18164 20996 18176
rect 21048 18164 21054 18216
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 20898 18096 20904 18148
rect 20956 18136 20962 18148
rect 21284 18136 21312 18167
rect 22554 18164 22560 18216
rect 22612 18204 22618 18216
rect 23017 18207 23075 18213
rect 23017 18204 23029 18207
rect 22612 18176 23029 18204
rect 22612 18164 22618 18176
rect 23017 18173 23029 18176
rect 23063 18173 23075 18207
rect 23017 18167 23075 18173
rect 27522 18164 27528 18216
rect 27580 18204 27586 18216
rect 27893 18207 27951 18213
rect 27893 18204 27905 18207
rect 27580 18176 27905 18204
rect 27580 18164 27586 18176
rect 27893 18173 27905 18176
rect 27939 18173 27951 18207
rect 29012 18204 29040 18244
rect 30300 18244 31944 18272
rect 30300 18204 30328 18244
rect 31938 18232 31944 18244
rect 31996 18232 32002 18284
rect 46750 18232 46756 18284
rect 46808 18272 46814 18284
rect 47949 18275 48007 18281
rect 47949 18272 47961 18275
rect 46808 18244 47961 18272
rect 46808 18232 46814 18244
rect 47949 18241 47961 18244
rect 47995 18241 48007 18275
rect 47949 18235 48007 18241
rect 29012 18176 30328 18204
rect 27893 18167 27951 18173
rect 30374 18164 30380 18216
rect 30432 18164 30438 18216
rect 32309 18207 32367 18213
rect 32309 18204 32321 18207
rect 31726 18176 32321 18204
rect 20956 18108 21312 18136
rect 20956 18096 20962 18108
rect 30190 18096 30196 18148
rect 30248 18136 30254 18148
rect 31726 18136 31754 18176
rect 32309 18173 32321 18176
rect 32355 18173 32367 18207
rect 32309 18167 32367 18173
rect 34517 18207 34575 18213
rect 34517 18173 34529 18207
rect 34563 18204 34575 18207
rect 34563 18176 34652 18204
rect 34563 18173 34575 18176
rect 34517 18167 34575 18173
rect 30248 18108 31754 18136
rect 30248 18096 30254 18108
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 19429 18071 19487 18077
rect 19429 18068 19441 18071
rect 15712 18040 19441 18068
rect 15712 18028 15718 18040
rect 19429 18037 19441 18040
rect 19475 18037 19487 18071
rect 19429 18031 19487 18037
rect 22462 18028 22468 18080
rect 22520 18068 22526 18080
rect 27890 18068 27896 18080
rect 22520 18040 27896 18068
rect 22520 18028 22526 18040
rect 27890 18028 27896 18040
rect 27948 18028 27954 18080
rect 34624 18068 34652 18176
rect 34790 18164 34796 18216
rect 34848 18204 34854 18216
rect 35342 18204 35348 18216
rect 34848 18176 35348 18204
rect 34848 18164 34854 18176
rect 35342 18164 35348 18176
rect 35400 18164 35406 18216
rect 38010 18164 38016 18216
rect 38068 18204 38074 18216
rect 38105 18207 38163 18213
rect 38105 18204 38117 18207
rect 38068 18176 38117 18204
rect 38068 18164 38074 18176
rect 38105 18173 38117 18176
rect 38151 18204 38163 18207
rect 38562 18204 38568 18216
rect 38151 18176 38568 18204
rect 38151 18173 38163 18176
rect 38105 18167 38163 18173
rect 38562 18164 38568 18176
rect 38620 18164 38626 18216
rect 49142 18164 49148 18216
rect 49200 18164 49206 18216
rect 34882 18068 34888 18080
rect 34624 18040 34888 18068
rect 34882 18028 34888 18040
rect 34940 18028 34946 18080
rect 35894 18028 35900 18080
rect 35952 18068 35958 18080
rect 36265 18071 36323 18077
rect 36265 18068 36277 18071
rect 35952 18040 36277 18068
rect 35952 18028 35958 18040
rect 36265 18037 36277 18040
rect 36311 18037 36323 18071
rect 36265 18031 36323 18037
rect 37461 18071 37519 18077
rect 37461 18037 37473 18071
rect 37507 18068 37519 18071
rect 39758 18068 39764 18080
rect 37507 18040 39764 18068
rect 37507 18037 37519 18040
rect 37461 18031 37519 18037
rect 39758 18028 39764 18040
rect 39816 18028 39822 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 19889 17867 19947 17873
rect 19889 17833 19901 17867
rect 19935 17864 19947 17867
rect 20070 17864 20076 17876
rect 19935 17836 20076 17864
rect 19935 17833 19947 17836
rect 19889 17827 19947 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 27338 17824 27344 17876
rect 27396 17824 27402 17876
rect 32401 17867 32459 17873
rect 32401 17833 32413 17867
rect 32447 17864 32459 17867
rect 32490 17864 32496 17876
rect 32447 17836 32496 17864
rect 32447 17833 32459 17836
rect 32401 17827 32459 17833
rect 32490 17824 32496 17836
rect 32548 17824 32554 17876
rect 37277 17867 37335 17873
rect 33060 17836 36860 17864
rect 27430 17756 27436 17808
rect 27488 17796 27494 17808
rect 28902 17796 28908 17808
rect 27488 17768 28908 17796
rect 27488 17756 27494 17768
rect 20530 17688 20536 17740
rect 20588 17688 20594 17740
rect 20990 17688 20996 17740
rect 21048 17728 21054 17740
rect 21361 17731 21419 17737
rect 21361 17728 21373 17731
rect 21048 17700 21373 17728
rect 21048 17688 21054 17700
rect 21361 17697 21373 17700
rect 21407 17728 21419 17731
rect 21450 17728 21456 17740
rect 21407 17700 21456 17728
rect 21407 17697 21419 17700
rect 21361 17691 21419 17697
rect 21450 17688 21456 17700
rect 21508 17688 21514 17740
rect 22370 17688 22376 17740
rect 22428 17728 22434 17740
rect 23109 17731 23167 17737
rect 23109 17728 23121 17731
rect 22428 17700 23121 17728
rect 22428 17688 22434 17700
rect 23109 17697 23121 17700
rect 23155 17728 23167 17731
rect 27522 17728 27528 17740
rect 23155 17700 27528 17728
rect 23155 17697 23167 17700
rect 23109 17691 23167 17697
rect 27522 17688 27528 17700
rect 27580 17688 27586 17740
rect 27908 17737 27936 17768
rect 28902 17756 28908 17768
rect 28960 17756 28966 17808
rect 27893 17731 27951 17737
rect 27893 17697 27905 17731
rect 27939 17697 27951 17731
rect 27893 17691 27951 17697
rect 29730 17688 29736 17740
rect 29788 17728 29794 17740
rect 30190 17728 30196 17740
rect 29788 17700 30196 17728
rect 29788 17688 29794 17700
rect 30190 17688 30196 17700
rect 30248 17728 30254 17740
rect 30653 17731 30711 17737
rect 30653 17728 30665 17731
rect 30248 17700 30665 17728
rect 30248 17688 30254 17700
rect 30653 17697 30665 17700
rect 30699 17697 30711 17731
rect 30653 17691 30711 17697
rect 31018 17688 31024 17740
rect 31076 17728 31082 17740
rect 32214 17728 32220 17740
rect 31076 17700 32220 17728
rect 31076 17688 31082 17700
rect 32214 17688 32220 17700
rect 32272 17728 32278 17740
rect 33060 17728 33088 17836
rect 36832 17796 36860 17836
rect 37277 17833 37289 17867
rect 37323 17864 37335 17867
rect 37366 17864 37372 17876
rect 37323 17836 37372 17864
rect 37323 17833 37335 17836
rect 37277 17827 37335 17833
rect 37366 17824 37372 17836
rect 37424 17824 37430 17876
rect 38194 17864 38200 17876
rect 37476 17836 38200 17864
rect 37476 17796 37504 17836
rect 38194 17824 38200 17836
rect 38252 17824 38258 17876
rect 36832 17768 37504 17796
rect 32272 17700 33088 17728
rect 32272 17688 32278 17700
rect 33778 17688 33784 17740
rect 33836 17688 33842 17740
rect 33965 17731 34023 17737
rect 33965 17697 33977 17731
rect 34011 17697 34023 17731
rect 33965 17691 34023 17697
rect 35529 17731 35587 17737
rect 35529 17697 35541 17731
rect 35575 17728 35587 17731
rect 35802 17728 35808 17740
rect 35575 17700 35808 17728
rect 35575 17697 35587 17700
rect 35529 17691 35587 17697
rect 19242 17620 19248 17672
rect 19300 17660 19306 17672
rect 21085 17663 21143 17669
rect 21085 17660 21097 17663
rect 19300 17632 21097 17660
rect 19300 17620 19306 17632
rect 21085 17629 21097 17632
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 23198 17620 23204 17672
rect 23256 17660 23262 17672
rect 23753 17663 23811 17669
rect 23753 17660 23765 17663
rect 23256 17632 23765 17660
rect 23256 17620 23262 17632
rect 23753 17629 23765 17632
rect 23799 17629 23811 17663
rect 23753 17623 23811 17629
rect 27614 17620 27620 17672
rect 27672 17660 27678 17672
rect 27709 17663 27767 17669
rect 27709 17660 27721 17663
rect 27672 17632 27721 17660
rect 27672 17620 27678 17632
rect 27709 17629 27721 17632
rect 27755 17629 27767 17663
rect 27709 17623 27767 17629
rect 27801 17663 27859 17669
rect 27801 17629 27813 17663
rect 27847 17660 27859 17663
rect 28442 17660 28448 17672
rect 27847 17632 28448 17660
rect 27847 17629 27859 17632
rect 27801 17623 27859 17629
rect 28442 17620 28448 17632
rect 28500 17660 28506 17672
rect 28626 17660 28632 17672
rect 28500 17632 28632 17660
rect 28500 17620 28506 17632
rect 28626 17620 28632 17632
rect 28684 17620 28690 17672
rect 33870 17660 33876 17672
rect 32062 17646 33876 17660
rect 32048 17632 33876 17646
rect 23290 17592 23296 17604
rect 22586 17564 23296 17592
rect 23290 17552 23296 17564
rect 23348 17592 23354 17604
rect 23566 17592 23572 17604
rect 23348 17564 23572 17592
rect 23348 17552 23354 17564
rect 23566 17552 23572 17564
rect 23624 17552 23630 17604
rect 30009 17595 30067 17601
rect 30009 17561 30021 17595
rect 30055 17592 30067 17595
rect 30282 17592 30288 17604
rect 30055 17564 30288 17592
rect 30055 17561 30067 17564
rect 30009 17555 30067 17561
rect 30282 17552 30288 17564
rect 30340 17552 30346 17604
rect 30926 17552 30932 17604
rect 30984 17552 30990 17604
rect 19978 17484 19984 17536
rect 20036 17524 20042 17536
rect 20257 17527 20315 17533
rect 20257 17524 20269 17527
rect 20036 17496 20269 17524
rect 20036 17484 20042 17496
rect 20257 17493 20269 17496
rect 20303 17493 20315 17527
rect 20257 17487 20315 17493
rect 20349 17527 20407 17533
rect 20349 17493 20361 17527
rect 20395 17524 20407 17527
rect 22738 17524 22744 17536
rect 20395 17496 22744 17524
rect 20395 17493 20407 17496
rect 20349 17487 20407 17493
rect 22738 17484 22744 17496
rect 22796 17484 22802 17536
rect 29362 17484 29368 17536
rect 29420 17524 29426 17536
rect 30101 17527 30159 17533
rect 30101 17524 30113 17527
rect 29420 17496 30113 17524
rect 29420 17484 29426 17496
rect 30101 17493 30113 17496
rect 30147 17493 30159 17527
rect 30101 17487 30159 17493
rect 30558 17484 30564 17536
rect 30616 17524 30622 17536
rect 32048 17524 32076 17632
rect 33870 17620 33876 17632
rect 33928 17620 33934 17672
rect 33980 17592 34008 17691
rect 35802 17688 35808 17700
rect 35860 17728 35866 17740
rect 37274 17728 37280 17740
rect 35860 17700 37280 17728
rect 35860 17688 35866 17700
rect 37274 17688 37280 17700
rect 37332 17728 37338 17740
rect 37737 17731 37795 17737
rect 37737 17728 37749 17731
rect 37332 17700 37749 17728
rect 37332 17688 37338 17700
rect 37737 17697 37749 17700
rect 37783 17697 37795 17731
rect 37737 17691 37795 17697
rect 38010 17688 38016 17740
rect 38068 17688 38074 17740
rect 44637 17731 44695 17737
rect 44637 17697 44649 17731
rect 44683 17728 44695 17731
rect 44683 17700 45048 17728
rect 44683 17697 44695 17700
rect 44637 17691 44695 17697
rect 42794 17620 42800 17672
rect 42852 17660 42858 17672
rect 42981 17663 43039 17669
rect 42981 17660 42993 17663
rect 42852 17632 42993 17660
rect 42852 17620 42858 17632
rect 42981 17629 42993 17632
rect 43027 17629 43039 17663
rect 42981 17623 43039 17629
rect 43346 17620 43352 17672
rect 43404 17660 43410 17672
rect 43717 17663 43775 17669
rect 43717 17660 43729 17663
rect 43404 17632 43729 17660
rect 43404 17620 43410 17632
rect 43717 17629 43729 17632
rect 43763 17629 43775 17663
rect 43717 17623 43775 17629
rect 43901 17663 43959 17669
rect 43901 17629 43913 17663
rect 43947 17660 43959 17663
rect 43947 17632 44680 17660
rect 43947 17629 43959 17632
rect 43901 17623 43959 17629
rect 35805 17595 35863 17601
rect 35805 17592 35817 17595
rect 33336 17564 33916 17592
rect 33980 17564 35817 17592
rect 33336 17533 33364 17564
rect 30616 17496 32076 17524
rect 33321 17527 33379 17533
rect 30616 17484 30622 17496
rect 33321 17493 33333 17527
rect 33367 17493 33379 17527
rect 33321 17487 33379 17493
rect 33686 17484 33692 17536
rect 33744 17484 33750 17536
rect 33888 17524 33916 17564
rect 35805 17561 35817 17564
rect 35851 17592 35863 17595
rect 35894 17592 35900 17604
rect 35851 17564 35900 17592
rect 35851 17561 35863 17564
rect 35805 17555 35863 17561
rect 35894 17552 35900 17564
rect 35952 17552 35958 17604
rect 36538 17552 36544 17604
rect 36596 17552 36602 17604
rect 37090 17552 37096 17604
rect 37148 17592 37154 17604
rect 37148 17564 37872 17592
rect 37148 17552 37154 17564
rect 37734 17524 37740 17536
rect 33888 17496 37740 17524
rect 37734 17484 37740 17496
rect 37792 17484 37798 17536
rect 37844 17524 37872 17564
rect 38654 17552 38660 17604
rect 38712 17552 38718 17604
rect 44450 17552 44456 17604
rect 44508 17552 44514 17604
rect 39485 17527 39543 17533
rect 39485 17524 39497 17527
rect 37844 17496 39497 17524
rect 39485 17493 39497 17496
rect 39531 17493 39543 17527
rect 39485 17487 39543 17493
rect 43073 17527 43131 17533
rect 43073 17493 43085 17527
rect 43119 17524 43131 17527
rect 44542 17524 44548 17536
rect 43119 17496 44548 17524
rect 43119 17493 43131 17496
rect 43073 17487 43131 17493
rect 44542 17484 44548 17496
rect 44600 17484 44606 17536
rect 44652 17524 44680 17632
rect 45020 17592 45048 17700
rect 45186 17620 45192 17672
rect 45244 17660 45250 17672
rect 47949 17663 48007 17669
rect 47949 17660 47961 17663
rect 45244 17632 47961 17660
rect 45244 17620 45250 17632
rect 47949 17629 47961 17632
rect 47995 17629 48007 17663
rect 47949 17623 48007 17629
rect 46842 17592 46848 17604
rect 45020 17564 46848 17592
rect 46842 17552 46848 17564
rect 46900 17552 46906 17604
rect 49142 17552 49148 17604
rect 49200 17552 49206 17604
rect 46658 17524 46664 17536
rect 44652 17496 46664 17524
rect 46658 17484 46664 17496
rect 46716 17484 46722 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 20898 17320 20904 17332
rect 19996 17292 20904 17320
rect 19996 17261 20024 17292
rect 20898 17280 20904 17292
rect 20956 17320 20962 17332
rect 20956 17292 21404 17320
rect 20956 17280 20962 17292
rect 19981 17255 20039 17261
rect 19981 17221 19993 17255
rect 20027 17221 20039 17255
rect 21376 17252 21404 17292
rect 21450 17280 21456 17332
rect 21508 17280 21514 17332
rect 22830 17280 22836 17332
rect 22888 17280 22894 17332
rect 23198 17280 23204 17332
rect 23256 17280 23262 17332
rect 24397 17323 24455 17329
rect 24397 17289 24409 17323
rect 24443 17320 24455 17323
rect 25958 17320 25964 17332
rect 24443 17292 25964 17320
rect 24443 17289 24455 17292
rect 24397 17283 24455 17289
rect 25958 17280 25964 17292
rect 26016 17280 26022 17332
rect 26326 17280 26332 17332
rect 26384 17320 26390 17332
rect 27249 17323 27307 17329
rect 27249 17320 27261 17323
rect 26384 17292 27261 17320
rect 26384 17280 26390 17292
rect 27249 17289 27261 17292
rect 27295 17289 27307 17323
rect 27249 17283 27307 17289
rect 28813 17323 28871 17329
rect 28813 17289 28825 17323
rect 28859 17320 28871 17323
rect 31018 17320 31024 17332
rect 28859 17292 31024 17320
rect 28859 17289 28871 17292
rect 28813 17283 28871 17289
rect 31018 17280 31024 17292
rect 31076 17280 31082 17332
rect 31110 17280 31116 17332
rect 31168 17320 31174 17332
rect 33965 17323 34023 17329
rect 33965 17320 33977 17323
rect 31168 17292 33977 17320
rect 31168 17280 31174 17292
rect 33965 17289 33977 17292
rect 34011 17289 34023 17323
rect 33965 17283 34023 17289
rect 34057 17323 34115 17329
rect 34057 17289 34069 17323
rect 34103 17320 34115 17323
rect 34422 17320 34428 17332
rect 34103 17292 34428 17320
rect 34103 17289 34115 17292
rect 34057 17283 34115 17289
rect 34422 17280 34428 17292
rect 34480 17280 34486 17332
rect 36538 17280 36544 17332
rect 36596 17320 36602 17332
rect 38654 17320 38660 17332
rect 36596 17292 38660 17320
rect 36596 17280 36602 17292
rect 38654 17280 38660 17292
rect 38712 17280 38718 17332
rect 23382 17252 23388 17264
rect 21376 17224 23388 17252
rect 19981 17215 20039 17221
rect 23382 17212 23388 17224
rect 23440 17252 23446 17264
rect 23440 17224 24440 17252
rect 23440 17212 23446 17224
rect 21082 17144 21088 17196
rect 21140 17184 21146 17196
rect 23198 17184 23204 17196
rect 21140 17156 23204 17184
rect 21140 17144 21146 17156
rect 23198 17144 23204 17156
rect 23256 17144 23262 17196
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17184 23351 17187
rect 24026 17184 24032 17196
rect 23339 17156 24032 17184
rect 23339 17153 23351 17156
rect 23293 17147 23351 17153
rect 24026 17144 24032 17156
rect 24084 17184 24090 17196
rect 24302 17184 24308 17196
rect 24084 17156 24308 17184
rect 24084 17144 24090 17156
rect 24302 17144 24308 17156
rect 24360 17144 24366 17196
rect 19242 17076 19248 17128
rect 19300 17116 19306 17128
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19300 17088 19717 17116
rect 19300 17076 19306 17088
rect 19705 17085 19717 17088
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 21910 17076 21916 17128
rect 21968 17116 21974 17128
rect 23385 17119 23443 17125
rect 23385 17116 23397 17119
rect 21968 17088 23397 17116
rect 21968 17076 21974 17088
rect 23385 17085 23397 17088
rect 23431 17116 23443 17119
rect 24412 17116 24440 17224
rect 25038 17212 25044 17264
rect 25096 17252 25102 17264
rect 25096 17224 27844 17252
rect 25096 17212 25102 17224
rect 24489 17187 24547 17193
rect 24489 17153 24501 17187
rect 24535 17184 24547 17187
rect 25866 17184 25872 17196
rect 24535 17156 25872 17184
rect 24535 17153 24547 17156
rect 24489 17147 24547 17153
rect 25866 17144 25872 17156
rect 25924 17144 25930 17196
rect 27617 17187 27675 17193
rect 27617 17153 27629 17187
rect 27663 17153 27675 17187
rect 27617 17147 27675 17153
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 23431 17088 24348 17116
rect 24412 17088 24593 17116
rect 23431 17085 23443 17088
rect 23385 17079 23443 17085
rect 21266 17008 21272 17060
rect 21324 17048 21330 17060
rect 24029 17051 24087 17057
rect 24029 17048 24041 17051
rect 21324 17020 24041 17048
rect 21324 17008 21330 17020
rect 24029 17017 24041 17020
rect 24075 17017 24087 17051
rect 24320 17048 24348 17088
rect 24581 17085 24593 17088
rect 24627 17085 24639 17119
rect 24581 17079 24639 17085
rect 26602 17048 26608 17060
rect 24320 17020 26608 17048
rect 24029 17011 24087 17017
rect 26602 17008 26608 17020
rect 26660 17008 26666 17060
rect 27632 17048 27660 17147
rect 27706 17076 27712 17128
rect 27764 17076 27770 17128
rect 27816 17125 27844 17224
rect 30558 17212 30564 17264
rect 30616 17252 30622 17264
rect 37550 17252 37556 17264
rect 30616 17224 30774 17252
rect 33612 17224 37556 17252
rect 30616 17212 30622 17224
rect 28718 17144 28724 17196
rect 28776 17184 28782 17196
rect 29546 17184 29552 17196
rect 28776 17156 29552 17184
rect 28776 17144 28782 17156
rect 27801 17119 27859 17125
rect 27801 17085 27813 17119
rect 27847 17116 27859 17119
rect 28166 17116 28172 17128
rect 27847 17088 28172 17116
rect 27847 17085 27859 17088
rect 27801 17079 27859 17085
rect 28166 17076 28172 17088
rect 28224 17076 28230 17128
rect 28350 17076 28356 17128
rect 28408 17116 28414 17128
rect 29012 17125 29040 17156
rect 29546 17144 29552 17156
rect 29604 17144 29610 17196
rect 32398 17144 32404 17196
rect 32456 17184 32462 17196
rect 32493 17187 32551 17193
rect 32493 17184 32505 17187
rect 32456 17156 32505 17184
rect 32456 17144 32462 17156
rect 32493 17153 32505 17156
rect 32539 17153 32551 17187
rect 32493 17147 32551 17153
rect 28905 17119 28963 17125
rect 28905 17116 28917 17119
rect 28408 17088 28917 17116
rect 28408 17076 28414 17088
rect 28905 17085 28917 17088
rect 28951 17085 28963 17119
rect 28905 17079 28963 17085
rect 28997 17119 29055 17125
rect 28997 17085 29009 17119
rect 29043 17085 29055 17119
rect 28997 17079 29055 17085
rect 29730 17076 29736 17128
rect 29788 17116 29794 17128
rect 30009 17119 30067 17125
rect 30009 17116 30021 17119
rect 29788 17088 30021 17116
rect 29788 17076 29794 17088
rect 30009 17085 30021 17088
rect 30055 17085 30067 17119
rect 30009 17079 30067 17085
rect 30282 17076 30288 17128
rect 30340 17076 30346 17128
rect 30926 17076 30932 17128
rect 30984 17116 30990 17128
rect 31757 17119 31815 17125
rect 31757 17116 31769 17119
rect 30984 17088 31769 17116
rect 30984 17076 30990 17088
rect 31757 17085 31769 17088
rect 31803 17116 31815 17119
rect 33502 17116 33508 17128
rect 31803 17088 33508 17116
rect 31803 17085 31815 17088
rect 31757 17079 31815 17085
rect 33502 17076 33508 17088
rect 33560 17076 33566 17128
rect 33612 17057 33640 17224
rect 37550 17212 37556 17224
rect 37608 17212 37614 17264
rect 43714 17212 43720 17264
rect 43772 17212 43778 17264
rect 35161 17187 35219 17193
rect 33704 17156 34376 17184
rect 33597 17051 33655 17057
rect 27632 17020 29684 17048
rect 28442 16940 28448 16992
rect 28500 16940 28506 16992
rect 29656 16980 29684 17020
rect 33597 17017 33609 17051
rect 33643 17017 33655 17051
rect 33597 17011 33655 17017
rect 32122 16980 32128 16992
rect 29656 16952 32128 16980
rect 32122 16940 32128 16952
rect 32180 16940 32186 16992
rect 32306 16940 32312 16992
rect 32364 16940 32370 16992
rect 32858 16940 32864 16992
rect 32916 16980 32922 16992
rect 33704 16980 33732 17156
rect 34241 17119 34299 17125
rect 34241 17085 34253 17119
rect 34287 17085 34299 17119
rect 34348 17116 34376 17156
rect 35161 17153 35173 17187
rect 35207 17184 35219 17187
rect 36173 17187 36231 17193
rect 36173 17184 36185 17187
rect 35207 17156 36185 17184
rect 35207 17153 35219 17156
rect 35161 17147 35219 17153
rect 36173 17153 36185 17156
rect 36219 17153 36231 17187
rect 36173 17147 36231 17153
rect 35253 17119 35311 17125
rect 35253 17116 35265 17119
rect 34348 17088 35265 17116
rect 34241 17079 34299 17085
rect 35253 17085 35265 17088
rect 35299 17085 35311 17119
rect 35253 17079 35311 17085
rect 34256 17048 34284 17079
rect 35342 17076 35348 17128
rect 35400 17076 35406 17128
rect 35526 17048 35532 17060
rect 34256 17020 35532 17048
rect 35526 17008 35532 17020
rect 35584 17008 35590 17060
rect 39942 17048 39948 17060
rect 38028 17020 39948 17048
rect 32916 16952 33732 16980
rect 34793 16983 34851 16989
rect 32916 16940 32922 16952
rect 34793 16949 34805 16983
rect 34839 16980 34851 16983
rect 38028 16980 38056 17020
rect 39942 17008 39948 17020
rect 40000 17008 40006 17060
rect 43901 17051 43959 17057
rect 43901 17017 43913 17051
rect 43947 17048 43959 17051
rect 46750 17048 46756 17060
rect 43947 17020 46756 17048
rect 43947 17017 43959 17020
rect 43901 17011 43959 17017
rect 46750 17008 46756 17020
rect 46808 17008 46814 17060
rect 34839 16952 38056 16980
rect 34839 16949 34851 16952
rect 34793 16943 34851 16949
rect 38102 16940 38108 16992
rect 38160 16940 38166 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 22462 16776 22468 16788
rect 21652 16748 22468 16776
rect 18598 16600 18604 16652
rect 18656 16640 18662 16652
rect 19242 16640 19248 16652
rect 18656 16612 19248 16640
rect 18656 16600 18662 16612
rect 19242 16600 19248 16612
rect 19300 16640 19306 16652
rect 21652 16649 21680 16748
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 23382 16736 23388 16788
rect 23440 16736 23446 16788
rect 26513 16779 26571 16785
rect 26513 16745 26525 16779
rect 26559 16776 26571 16779
rect 26602 16776 26608 16788
rect 26559 16748 26608 16776
rect 26559 16745 26571 16748
rect 26513 16739 26571 16745
rect 26602 16736 26608 16748
rect 26660 16736 26666 16788
rect 27430 16736 27436 16788
rect 27488 16776 27494 16788
rect 31110 16776 31116 16788
rect 27488 16748 31116 16776
rect 27488 16736 27494 16748
rect 31110 16736 31116 16748
rect 31168 16736 31174 16788
rect 37090 16776 37096 16788
rect 34808 16748 37096 16776
rect 19429 16643 19487 16649
rect 19429 16640 19441 16643
rect 19300 16612 19441 16640
rect 19300 16600 19306 16612
rect 19429 16609 19441 16612
rect 19475 16640 19487 16643
rect 21637 16643 21695 16649
rect 21637 16640 21649 16643
rect 19475 16612 21649 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 21637 16609 21649 16612
rect 21683 16609 21695 16643
rect 21637 16603 21695 16609
rect 21910 16600 21916 16652
rect 21968 16600 21974 16652
rect 24394 16600 24400 16652
rect 24452 16640 24458 16652
rect 24762 16640 24768 16652
rect 24452 16612 24768 16640
rect 24452 16600 24458 16612
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 25038 16600 25044 16652
rect 25096 16600 25102 16652
rect 26786 16600 26792 16652
rect 26844 16640 26850 16652
rect 27709 16643 27767 16649
rect 27709 16640 27721 16643
rect 26844 16612 27721 16640
rect 26844 16600 26850 16612
rect 27709 16609 27721 16612
rect 27755 16609 27767 16643
rect 27709 16603 27767 16609
rect 28166 16600 28172 16652
rect 28224 16640 28230 16652
rect 28902 16640 28908 16652
rect 28224 16612 28908 16640
rect 28224 16600 28230 16612
rect 28902 16600 28908 16612
rect 28960 16600 28966 16652
rect 32030 16600 32036 16652
rect 32088 16640 32094 16652
rect 34057 16643 34115 16649
rect 34057 16640 34069 16643
rect 32088 16612 34069 16640
rect 32088 16600 32094 16612
rect 34057 16609 34069 16612
rect 34103 16609 34115 16643
rect 34057 16603 34115 16609
rect 34241 16643 34299 16649
rect 34241 16609 34253 16643
rect 34287 16640 34299 16643
rect 34808 16640 34836 16748
rect 37090 16736 37096 16748
rect 37148 16736 37154 16788
rect 34287 16612 34836 16640
rect 34287 16609 34299 16612
rect 34241 16603 34299 16609
rect 34882 16600 34888 16652
rect 34940 16600 34946 16652
rect 35161 16643 35219 16649
rect 35161 16609 35173 16643
rect 35207 16640 35219 16643
rect 35526 16640 35532 16652
rect 35207 16612 35532 16640
rect 35207 16609 35219 16612
rect 35161 16603 35219 16609
rect 35526 16600 35532 16612
rect 35584 16600 35590 16652
rect 37366 16600 37372 16652
rect 37424 16640 37430 16652
rect 38013 16643 38071 16649
rect 38013 16640 38025 16643
rect 37424 16612 38025 16640
rect 37424 16600 37430 16612
rect 38013 16609 38025 16612
rect 38059 16609 38071 16643
rect 38013 16603 38071 16609
rect 27525 16575 27583 16581
rect 27525 16541 27537 16575
rect 27571 16572 27583 16575
rect 28442 16572 28448 16584
rect 27571 16544 28448 16572
rect 27571 16541 27583 16544
rect 27525 16535 27583 16541
rect 28442 16532 28448 16544
rect 28500 16532 28506 16584
rect 30650 16532 30656 16584
rect 30708 16572 30714 16584
rect 33965 16575 34023 16581
rect 33965 16572 33977 16575
rect 30708 16544 33977 16572
rect 30708 16532 30714 16544
rect 33965 16541 33977 16544
rect 34011 16541 34023 16575
rect 33965 16535 34023 16541
rect 37829 16575 37887 16581
rect 37829 16541 37841 16575
rect 37875 16572 37887 16575
rect 38102 16572 38108 16584
rect 37875 16544 38108 16572
rect 37875 16541 37887 16544
rect 37829 16535 37887 16541
rect 38102 16532 38108 16544
rect 38160 16532 38166 16584
rect 46198 16532 46204 16584
rect 46256 16572 46262 16584
rect 47949 16575 48007 16581
rect 47949 16572 47961 16575
rect 46256 16544 47961 16572
rect 46256 16532 46262 16544
rect 47949 16541 47961 16544
rect 47995 16541 48007 16575
rect 47949 16535 48007 16541
rect 5537 16507 5595 16513
rect 5537 16473 5549 16507
rect 5583 16504 5595 16507
rect 9766 16504 9772 16516
rect 5583 16476 9772 16504
rect 5583 16473 5595 16476
rect 5537 16467 5595 16473
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 19705 16507 19763 16513
rect 19705 16473 19717 16507
rect 19751 16504 19763 16507
rect 19794 16504 19800 16516
rect 19751 16476 19800 16504
rect 19751 16473 19763 16476
rect 19705 16467 19763 16473
rect 19794 16464 19800 16476
rect 19852 16464 19858 16516
rect 23290 16504 23296 16516
rect 19904 16476 20194 16504
rect 23138 16476 23296 16504
rect 5626 16396 5632 16448
rect 5684 16396 5690 16448
rect 19242 16396 19248 16448
rect 19300 16436 19306 16448
rect 19904 16436 19932 16476
rect 23290 16464 23296 16476
rect 23348 16504 23354 16516
rect 24762 16504 24768 16516
rect 23348 16476 24768 16504
rect 23348 16464 23354 16476
rect 24762 16464 24768 16476
rect 24820 16504 24826 16516
rect 27617 16507 27675 16513
rect 24820 16476 25530 16504
rect 24820 16464 24826 16476
rect 27617 16473 27629 16507
rect 27663 16504 27675 16507
rect 28718 16504 28724 16516
rect 27663 16476 28724 16504
rect 27663 16473 27675 16476
rect 27617 16467 27675 16473
rect 28718 16464 28724 16476
rect 28776 16464 28782 16516
rect 35434 16504 35440 16516
rect 33612 16476 35440 16504
rect 21082 16436 21088 16448
rect 19300 16408 21088 16436
rect 19300 16396 19306 16408
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 21174 16396 21180 16448
rect 21232 16396 21238 16448
rect 26326 16396 26332 16448
rect 26384 16436 26390 16448
rect 27157 16439 27215 16445
rect 27157 16436 27169 16439
rect 26384 16408 27169 16436
rect 26384 16396 26390 16408
rect 27157 16405 27169 16408
rect 27203 16405 27215 16439
rect 27157 16399 27215 16405
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 28442 16436 28448 16448
rect 28316 16408 28448 16436
rect 28316 16396 28322 16408
rect 28442 16396 28448 16408
rect 28500 16396 28506 16448
rect 28810 16396 28816 16448
rect 28868 16436 28874 16448
rect 29730 16436 29736 16448
rect 28868 16408 29736 16436
rect 28868 16396 28874 16408
rect 29730 16396 29736 16408
rect 29788 16396 29794 16448
rect 33612 16445 33640 16476
rect 35434 16464 35440 16476
rect 35492 16464 35498 16516
rect 36538 16504 36544 16516
rect 36386 16476 36544 16504
rect 36538 16464 36544 16476
rect 36596 16464 36602 16516
rect 37734 16464 37740 16516
rect 37792 16504 37798 16516
rect 37921 16507 37979 16513
rect 37921 16504 37933 16507
rect 37792 16476 37933 16504
rect 37792 16464 37798 16476
rect 37921 16473 37933 16476
rect 37967 16473 37979 16507
rect 37921 16467 37979 16473
rect 49142 16464 49148 16516
rect 49200 16464 49206 16516
rect 33597 16439 33655 16445
rect 33597 16405 33609 16439
rect 33643 16405 33655 16439
rect 33597 16399 33655 16405
rect 36630 16396 36636 16448
rect 36688 16396 36694 16448
rect 37461 16439 37519 16445
rect 37461 16405 37473 16439
rect 37507 16436 37519 16439
rect 39482 16436 39488 16448
rect 37507 16408 39488 16436
rect 37507 16405 37519 16408
rect 37461 16399 37519 16405
rect 39482 16396 39488 16408
rect 39540 16396 39546 16448
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 19978 16192 19984 16244
rect 20036 16232 20042 16244
rect 25685 16235 25743 16241
rect 25685 16232 25697 16235
rect 20036 16204 25697 16232
rect 20036 16192 20042 16204
rect 25685 16201 25697 16204
rect 25731 16201 25743 16235
rect 25685 16195 25743 16201
rect 27154 16192 27160 16244
rect 27212 16192 27218 16244
rect 27430 16192 27436 16244
rect 27488 16232 27494 16244
rect 27617 16235 27675 16241
rect 27617 16232 27629 16235
rect 27488 16204 27629 16232
rect 27488 16192 27494 16204
rect 27617 16201 27629 16204
rect 27663 16201 27675 16235
rect 27617 16195 27675 16201
rect 28350 16192 28356 16244
rect 28408 16232 28414 16244
rect 33413 16235 33471 16241
rect 33413 16232 33425 16235
rect 28408 16204 33425 16232
rect 28408 16192 28414 16204
rect 33413 16201 33425 16204
rect 33459 16201 33471 16235
rect 33413 16195 33471 16201
rect 16574 16124 16580 16176
rect 16632 16164 16638 16176
rect 23017 16167 23075 16173
rect 23017 16164 23029 16167
rect 16632 16136 23029 16164
rect 16632 16124 16638 16136
rect 23017 16133 23029 16136
rect 23063 16133 23075 16167
rect 23017 16127 23075 16133
rect 24670 16124 24676 16176
rect 24728 16164 24734 16176
rect 24765 16167 24823 16173
rect 24765 16164 24777 16167
rect 24728 16136 24777 16164
rect 24728 16124 24734 16136
rect 24765 16133 24777 16136
rect 24811 16133 24823 16167
rect 24765 16127 24823 16133
rect 26878 16124 26884 16176
rect 26936 16164 26942 16176
rect 27525 16167 27583 16173
rect 27525 16164 27537 16167
rect 26936 16136 27537 16164
rect 26936 16124 26942 16136
rect 27525 16133 27537 16136
rect 27571 16164 27583 16167
rect 29362 16164 29368 16176
rect 27571 16136 29368 16164
rect 27571 16133 27583 16136
rect 27525 16127 27583 16133
rect 29362 16124 29368 16136
rect 29420 16124 29426 16176
rect 30466 16164 30472 16176
rect 30314 16136 30472 16164
rect 30466 16124 30472 16136
rect 30524 16124 30530 16176
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 2774 16096 2780 16108
rect 1811 16068 2780 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 33321 16099 33379 16105
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 22462 15988 22468 16040
rect 22520 16028 22526 16040
rect 22741 16031 22799 16037
rect 22741 16028 22753 16031
rect 22520 16000 22753 16028
rect 22520 15988 22526 16000
rect 22741 15997 22753 16000
rect 22787 15997 22799 16031
rect 24136 16028 24164 16082
rect 33321 16065 33333 16099
rect 33367 16096 33379 16099
rect 34333 16099 34391 16105
rect 34333 16096 34345 16099
rect 33367 16068 34345 16096
rect 33367 16065 33379 16068
rect 33321 16059 33379 16065
rect 34333 16065 34345 16068
rect 34379 16065 34391 16099
rect 34333 16059 34391 16065
rect 36265 16099 36323 16105
rect 36265 16065 36277 16099
rect 36311 16096 36323 16099
rect 36446 16096 36452 16108
rect 36311 16068 36452 16096
rect 36311 16065 36323 16068
rect 36265 16059 36323 16065
rect 36446 16056 36452 16068
rect 36504 16056 36510 16108
rect 38933 16099 38991 16105
rect 38933 16065 38945 16099
rect 38979 16096 38991 16099
rect 40034 16096 40040 16108
rect 38979 16068 40040 16096
rect 38979 16065 38991 16068
rect 38933 16059 38991 16065
rect 40034 16056 40040 16068
rect 40092 16056 40098 16108
rect 47854 16056 47860 16108
rect 47912 16096 47918 16108
rect 47949 16099 48007 16105
rect 47949 16096 47961 16099
rect 47912 16068 47961 16096
rect 47912 16056 47918 16068
rect 47949 16065 47961 16068
rect 47995 16065 48007 16099
rect 47949 16059 48007 16065
rect 24762 16028 24768 16040
rect 24136 16000 24768 16028
rect 22741 15991 22799 15997
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 25777 16031 25835 16037
rect 25777 15997 25789 16031
rect 25823 15997 25835 16031
rect 25777 15991 25835 15997
rect 25961 16031 26019 16037
rect 25961 15997 25973 16031
rect 26007 16028 26019 16031
rect 26142 16028 26148 16040
rect 26007 16000 26148 16028
rect 26007 15997 26019 16000
rect 25961 15991 26019 15997
rect 25792 15960 25820 15991
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 27522 15988 27528 16040
rect 27580 16028 27586 16040
rect 27709 16031 27767 16037
rect 27709 16028 27721 16031
rect 27580 16000 27721 16028
rect 27580 15988 27586 16000
rect 27709 15997 27721 16000
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 27798 15988 27804 16040
rect 27856 16028 27862 16040
rect 28810 16028 28816 16040
rect 27856 16000 28816 16028
rect 27856 15988 27862 16000
rect 28810 15988 28816 16000
rect 28868 15988 28874 16040
rect 29089 16031 29147 16037
rect 29089 15997 29101 16031
rect 29135 16028 29147 16031
rect 29454 16028 29460 16040
rect 29135 16000 29460 16028
rect 29135 15997 29147 16000
rect 29089 15991 29147 15997
rect 29454 15988 29460 16000
rect 29512 15988 29518 16040
rect 32490 16028 32496 16040
rect 30116 16000 32496 16028
rect 25792 15932 28856 15960
rect 25317 15895 25375 15901
rect 25317 15861 25329 15895
rect 25363 15892 25375 15895
rect 28258 15892 28264 15904
rect 25363 15864 28264 15892
rect 25363 15861 25375 15864
rect 25317 15855 25375 15861
rect 28258 15852 28264 15864
rect 28316 15852 28322 15904
rect 28828 15892 28856 15932
rect 29638 15892 29644 15904
rect 28828 15864 29644 15892
rect 29638 15852 29644 15864
rect 29696 15892 29702 15904
rect 30116 15892 30144 16000
rect 32490 15988 32496 16000
rect 32548 15988 32554 16040
rect 33597 16031 33655 16037
rect 33597 15997 33609 16031
rect 33643 16028 33655 16031
rect 37458 16028 37464 16040
rect 33643 16000 37464 16028
rect 33643 15997 33655 16000
rect 33597 15991 33655 15997
rect 37458 15988 37464 16000
rect 37516 15988 37522 16040
rect 49142 15988 49148 16040
rect 49200 15988 49206 16040
rect 32953 15963 33011 15969
rect 32953 15929 32965 15963
rect 32999 15960 33011 15963
rect 35066 15960 35072 15972
rect 32999 15932 35072 15960
rect 32999 15929 33011 15932
rect 32953 15923 33011 15929
rect 35066 15920 35072 15932
rect 35124 15920 35130 15972
rect 29696 15864 30144 15892
rect 29696 15852 29702 15864
rect 30558 15852 30564 15904
rect 30616 15892 30622 15904
rect 32858 15892 32864 15904
rect 30616 15864 32864 15892
rect 30616 15852 30622 15864
rect 32858 15852 32864 15864
rect 32916 15852 32922 15904
rect 33410 15852 33416 15904
rect 33468 15892 33474 15904
rect 34977 15895 35035 15901
rect 34977 15892 34989 15895
rect 33468 15864 34989 15892
rect 33468 15852 33474 15864
rect 34977 15861 34989 15864
rect 35023 15861 35035 15895
rect 34977 15855 35035 15861
rect 36081 15895 36139 15901
rect 36081 15861 36093 15895
rect 36127 15892 36139 15895
rect 36446 15892 36452 15904
rect 36127 15864 36452 15892
rect 36127 15861 36139 15864
rect 36081 15855 36139 15861
rect 36446 15852 36452 15864
rect 36504 15852 36510 15904
rect 37642 15852 37648 15904
rect 37700 15852 37706 15904
rect 38470 15852 38476 15904
rect 38528 15892 38534 15904
rect 38749 15895 38807 15901
rect 38749 15892 38761 15895
rect 38528 15864 38761 15892
rect 38528 15852 38534 15864
rect 38749 15861 38761 15864
rect 38795 15861 38807 15895
rect 38749 15855 38807 15861
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 26510 15648 26516 15700
rect 26568 15648 26574 15700
rect 28810 15648 28816 15700
rect 28868 15688 28874 15700
rect 29454 15688 29460 15700
rect 28868 15660 29460 15688
rect 28868 15648 28874 15660
rect 29454 15648 29460 15660
rect 29512 15648 29518 15700
rect 30190 15648 30196 15700
rect 30248 15688 30254 15700
rect 31481 15691 31539 15697
rect 31481 15688 31493 15691
rect 30248 15660 31493 15688
rect 30248 15648 30254 15660
rect 31481 15657 31493 15660
rect 31527 15657 31539 15691
rect 31481 15651 31539 15657
rect 33045 15691 33103 15697
rect 33045 15657 33057 15691
rect 33091 15688 33103 15691
rect 39114 15688 39120 15700
rect 33091 15660 39120 15688
rect 33091 15657 33103 15660
rect 33045 15651 33103 15657
rect 39114 15648 39120 15660
rect 39172 15648 39178 15700
rect 21358 15580 21364 15632
rect 21416 15620 21422 15632
rect 27709 15623 27767 15629
rect 21416 15592 22094 15620
rect 21416 15580 21422 15592
rect 22066 15484 22094 15592
rect 27709 15589 27721 15623
rect 27755 15620 27767 15623
rect 29638 15620 29644 15632
rect 27755 15592 28856 15620
rect 27755 15589 27767 15592
rect 27709 15583 27767 15589
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 26053 15555 26111 15561
rect 26053 15552 26065 15555
rect 24176 15524 26065 15552
rect 24176 15512 24182 15524
rect 26053 15521 26065 15524
rect 26099 15521 26111 15555
rect 26053 15515 26111 15521
rect 27157 15555 27215 15561
rect 27157 15521 27169 15555
rect 27203 15552 27215 15555
rect 27338 15552 27344 15564
rect 27203 15524 27344 15552
rect 27203 15521 27215 15524
rect 27157 15515 27215 15521
rect 27338 15512 27344 15524
rect 27396 15512 27402 15564
rect 27982 15512 27988 15564
rect 28040 15552 28046 15564
rect 28261 15555 28319 15561
rect 28261 15552 28273 15555
rect 28040 15524 28273 15552
rect 28040 15512 28046 15524
rect 28261 15521 28273 15524
rect 28307 15521 28319 15555
rect 28828 15552 28856 15592
rect 28966 15592 29644 15620
rect 28966 15552 28994 15592
rect 29638 15580 29644 15592
rect 29696 15580 29702 15632
rect 28828 15524 28994 15552
rect 28261 15515 28319 15521
rect 29730 15512 29736 15564
rect 29788 15512 29794 15564
rect 30009 15555 30067 15561
rect 30009 15521 30021 15555
rect 30055 15552 30067 15555
rect 30558 15552 30564 15564
rect 30055 15524 30564 15552
rect 30055 15521 30067 15524
rect 30009 15515 30067 15521
rect 30558 15512 30564 15524
rect 30616 15512 30622 15564
rect 33502 15512 33508 15564
rect 33560 15552 33566 15564
rect 33597 15555 33655 15561
rect 33597 15552 33609 15555
rect 33560 15524 33609 15552
rect 33560 15512 33566 15524
rect 33597 15521 33609 15524
rect 33643 15521 33655 15555
rect 33597 15515 33655 15521
rect 35802 15512 35808 15564
rect 35860 15512 35866 15564
rect 36081 15555 36139 15561
rect 36081 15521 36093 15555
rect 36127 15552 36139 15555
rect 37090 15552 37096 15564
rect 36127 15524 37096 15552
rect 36127 15521 36139 15524
rect 36081 15515 36139 15521
rect 37090 15512 37096 15524
rect 37148 15512 37154 15564
rect 28077 15487 28135 15493
rect 28077 15484 28089 15487
rect 22066 15456 28089 15484
rect 28077 15453 28089 15456
rect 28123 15453 28135 15487
rect 28077 15447 28135 15453
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15484 28227 15487
rect 28215 15456 29776 15484
rect 28215 15453 28227 15456
rect 28169 15447 28227 15453
rect 24673 15419 24731 15425
rect 24673 15385 24685 15419
rect 24719 15416 24731 15419
rect 25314 15416 25320 15428
rect 24719 15388 25320 15416
rect 24719 15385 24731 15388
rect 24673 15379 24731 15385
rect 25314 15376 25320 15388
rect 25372 15376 25378 15428
rect 25406 15376 25412 15428
rect 25464 15416 25470 15428
rect 25869 15419 25927 15425
rect 25869 15416 25881 15419
rect 25464 15388 25881 15416
rect 25464 15376 25470 15388
rect 25869 15385 25881 15388
rect 25915 15385 25927 15419
rect 25869 15379 25927 15385
rect 26878 15376 26884 15428
rect 26936 15376 26942 15428
rect 26973 15419 27031 15425
rect 26973 15385 26985 15419
rect 27019 15416 27031 15419
rect 27430 15416 27436 15428
rect 27019 15388 27436 15416
rect 27019 15385 27031 15388
rect 26973 15379 27031 15385
rect 27430 15376 27436 15388
rect 27488 15376 27494 15428
rect 28258 15376 28264 15428
rect 28316 15416 28322 15428
rect 28810 15416 28816 15428
rect 28316 15388 28816 15416
rect 28316 15376 28322 15388
rect 28810 15376 28816 15388
rect 28868 15376 28874 15428
rect 28997 15419 29055 15425
rect 28997 15385 29009 15419
rect 29043 15416 29055 15419
rect 29178 15416 29184 15428
rect 29043 15388 29184 15416
rect 29043 15385 29055 15388
rect 28997 15379 29055 15385
rect 29178 15376 29184 15388
rect 29236 15376 29242 15428
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 24765 15351 24823 15357
rect 24765 15348 24777 15351
rect 22704 15320 24777 15348
rect 22704 15308 22710 15320
rect 24765 15317 24777 15320
rect 24811 15317 24823 15351
rect 24765 15311 24823 15317
rect 27338 15308 27344 15360
rect 27396 15348 27402 15360
rect 29089 15351 29147 15357
rect 29089 15348 29101 15351
rect 27396 15320 29101 15348
rect 27396 15308 27402 15320
rect 29089 15317 29101 15320
rect 29135 15317 29147 15351
rect 29748 15348 29776 15456
rect 32582 15444 32588 15496
rect 32640 15444 32646 15496
rect 33410 15444 33416 15496
rect 33468 15444 33474 15496
rect 46842 15444 46848 15496
rect 46900 15484 46906 15496
rect 47949 15487 48007 15493
rect 47949 15484 47961 15487
rect 46900 15456 47961 15484
rect 46900 15444 46906 15456
rect 47949 15453 47961 15456
rect 47995 15453 48007 15487
rect 47949 15447 48007 15453
rect 30466 15376 30472 15428
rect 30524 15376 30530 15428
rect 33505 15419 33563 15425
rect 31404 15388 31754 15416
rect 31404 15348 31432 15388
rect 29748 15320 31432 15348
rect 31726 15348 31754 15388
rect 32324 15388 32536 15416
rect 32324 15348 32352 15388
rect 31726 15320 32352 15348
rect 29089 15311 29147 15317
rect 32398 15308 32404 15360
rect 32456 15308 32462 15360
rect 32508 15348 32536 15388
rect 33505 15385 33517 15419
rect 33551 15416 33563 15419
rect 33594 15416 33600 15428
rect 33551 15388 33600 15416
rect 33551 15385 33563 15388
rect 33505 15379 33563 15385
rect 33594 15376 33600 15388
rect 33652 15376 33658 15428
rect 36538 15376 36544 15428
rect 36596 15376 36602 15428
rect 49142 15376 49148 15428
rect 49200 15376 49206 15428
rect 34422 15348 34428 15360
rect 32508 15320 34428 15348
rect 34422 15308 34428 15320
rect 34480 15308 34486 15360
rect 37553 15351 37611 15357
rect 37553 15317 37565 15351
rect 37599 15348 37611 15351
rect 37734 15348 37740 15360
rect 37599 15320 37740 15348
rect 37599 15317 37611 15320
rect 37553 15311 37611 15317
rect 37734 15308 37740 15320
rect 37792 15308 37798 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 20070 15104 20076 15156
rect 20128 15144 20134 15156
rect 20993 15147 21051 15153
rect 20993 15144 21005 15147
rect 20128 15116 21005 15144
rect 20128 15104 20134 15116
rect 20993 15113 21005 15116
rect 21039 15113 21051 15147
rect 20993 15107 21051 15113
rect 24213 15147 24271 15153
rect 24213 15113 24225 15147
rect 24259 15144 24271 15147
rect 26142 15144 26148 15156
rect 24259 15116 26148 15144
rect 24259 15113 24271 15116
rect 24213 15107 24271 15113
rect 26142 15104 26148 15116
rect 26200 15104 26206 15156
rect 26329 15147 26387 15153
rect 26329 15113 26341 15147
rect 26375 15144 26387 15147
rect 28994 15144 29000 15156
rect 26375 15116 29000 15144
rect 26375 15113 26387 15116
rect 26329 15107 26387 15113
rect 28994 15104 29000 15116
rect 29052 15104 29058 15156
rect 29454 15104 29460 15156
rect 29512 15104 29518 15156
rect 29638 15104 29644 15156
rect 29696 15144 29702 15156
rect 32769 15147 32827 15153
rect 32769 15144 32781 15147
rect 29696 15116 32781 15144
rect 29696 15104 29702 15116
rect 32769 15113 32781 15116
rect 32815 15113 32827 15147
rect 32769 15107 32827 15113
rect 37642 15104 37648 15156
rect 37700 15144 37706 15156
rect 37829 15147 37887 15153
rect 37829 15144 37841 15147
rect 37700 15116 37841 15144
rect 37700 15104 37706 15116
rect 37829 15113 37841 15116
rect 37875 15113 37887 15147
rect 37829 15107 37887 15113
rect 24762 15076 24768 15088
rect 23966 15048 24768 15076
rect 24762 15036 24768 15048
rect 24820 15036 24826 15088
rect 30009 15079 30067 15085
rect 30009 15045 30021 15079
rect 30055 15076 30067 15079
rect 30098 15076 30104 15088
rect 30055 15048 30104 15076
rect 30055 15045 30067 15048
rect 30009 15039 30067 15045
rect 30098 15036 30104 15048
rect 30156 15036 30162 15088
rect 31570 15036 31576 15088
rect 31628 15036 31634 15088
rect 37550 15036 37556 15088
rect 37608 15076 37614 15088
rect 37921 15079 37979 15085
rect 37921 15076 37933 15079
rect 37608 15048 37933 15076
rect 37608 15036 37614 15048
rect 37921 15045 37933 15048
rect 37967 15045 37979 15079
rect 37921 15039 37979 15045
rect 17034 14968 17040 15020
rect 17092 15008 17098 15020
rect 20901 15011 20959 15017
rect 20901 15008 20913 15011
rect 17092 14980 20913 15008
rect 17092 14968 17098 14980
rect 20901 14977 20913 14980
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 22462 14968 22468 15020
rect 22520 14968 22526 15020
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 15008 26295 15011
rect 27614 15008 27620 15020
rect 26283 14980 27620 15008
rect 26283 14977 26295 14980
rect 26237 14971 26295 14977
rect 27614 14968 27620 14980
rect 27672 14968 27678 15020
rect 29086 14968 29092 15020
rect 29144 14968 29150 15020
rect 32214 14968 32220 15020
rect 32272 15008 32278 15020
rect 32677 15011 32735 15017
rect 32677 15008 32689 15011
rect 32272 14980 32689 15008
rect 32272 14968 32278 14980
rect 32677 14977 32689 14980
rect 32723 14977 32735 15011
rect 32677 14971 32735 14977
rect 39758 14968 39764 15020
rect 39816 15008 39822 15020
rect 41969 15011 42027 15017
rect 41969 15008 41981 15011
rect 39816 14980 41981 15008
rect 39816 14968 39822 14980
rect 41969 14977 41981 14980
rect 42015 14977 42027 15011
rect 41969 14971 42027 14977
rect 46750 14968 46756 15020
rect 46808 15008 46814 15020
rect 47949 15011 48007 15017
rect 47949 15008 47961 15011
rect 46808 14980 47961 15008
rect 46808 14968 46814 14980
rect 47949 14977 47961 14980
rect 47995 14977 48007 15011
rect 47949 14971 48007 14977
rect 21174 14900 21180 14952
rect 21232 14940 21238 14952
rect 22741 14943 22799 14949
rect 22741 14940 22753 14943
rect 21232 14912 22753 14940
rect 21232 14900 21238 14912
rect 22741 14909 22753 14912
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 26513 14943 26571 14949
rect 26513 14909 26525 14943
rect 26559 14940 26571 14943
rect 26602 14940 26608 14952
rect 26559 14912 26608 14940
rect 26559 14909 26571 14912
rect 26513 14903 26571 14909
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 27706 14900 27712 14952
rect 27764 14900 27770 14952
rect 27982 14900 27988 14952
rect 28040 14940 28046 14952
rect 30193 14943 30251 14949
rect 28040 14912 29040 14940
rect 28040 14900 28046 14912
rect 25866 14832 25872 14884
rect 25924 14832 25930 14884
rect 29012 14872 29040 14912
rect 30193 14909 30205 14943
rect 30239 14940 30251 14943
rect 31018 14940 31024 14952
rect 30239 14912 31024 14940
rect 30239 14909 30251 14912
rect 30193 14903 30251 14909
rect 31018 14900 31024 14912
rect 31076 14900 31082 14952
rect 32858 14900 32864 14952
rect 32916 14900 32922 14952
rect 36630 14900 36636 14952
rect 36688 14940 36694 14952
rect 38013 14943 38071 14949
rect 38013 14940 38025 14943
rect 36688 14912 38025 14940
rect 36688 14900 36694 14912
rect 38013 14909 38025 14912
rect 38059 14909 38071 14943
rect 38013 14903 38071 14909
rect 49142 14900 49148 14952
rect 49200 14900 49206 14952
rect 30282 14872 30288 14884
rect 29012 14844 30288 14872
rect 30282 14832 30288 14844
rect 30340 14832 30346 14884
rect 31757 14875 31815 14881
rect 31757 14841 31769 14875
rect 31803 14872 31815 14875
rect 33778 14872 33784 14884
rect 31803 14844 33784 14872
rect 31803 14841 31815 14844
rect 31757 14835 31815 14841
rect 33778 14832 33784 14844
rect 33836 14832 33842 14884
rect 20530 14764 20536 14816
rect 20588 14764 20594 14816
rect 30190 14764 30196 14816
rect 30248 14804 30254 14816
rect 30837 14807 30895 14813
rect 30837 14804 30849 14807
rect 30248 14776 30849 14804
rect 30248 14764 30254 14776
rect 30837 14773 30849 14776
rect 30883 14773 30895 14807
rect 30837 14767 30895 14773
rect 32309 14807 32367 14813
rect 32309 14773 32321 14807
rect 32355 14804 32367 14807
rect 37366 14804 37372 14816
rect 32355 14776 37372 14804
rect 32355 14773 32367 14776
rect 32309 14767 32367 14773
rect 37366 14764 37372 14776
rect 37424 14764 37430 14816
rect 37461 14807 37519 14813
rect 37461 14773 37473 14807
rect 37507 14804 37519 14807
rect 41322 14804 41328 14816
rect 37507 14776 41328 14804
rect 37507 14773 37519 14776
rect 37461 14767 37519 14773
rect 41322 14764 41328 14776
rect 41380 14764 41386 14816
rect 41785 14807 41843 14813
rect 41785 14773 41797 14807
rect 41831 14804 41843 14807
rect 44174 14804 44180 14816
rect 41831 14776 44180 14804
rect 41831 14773 41843 14776
rect 41785 14767 41843 14773
rect 44174 14764 44180 14776
rect 44232 14764 44238 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 20530 14560 20536 14612
rect 20588 14600 20594 14612
rect 30558 14600 30564 14612
rect 20588 14572 30564 14600
rect 20588 14560 20594 14572
rect 30558 14560 30564 14572
rect 30616 14560 30622 14612
rect 32214 14560 32220 14612
rect 32272 14560 32278 14612
rect 27617 14535 27675 14541
rect 27617 14501 27629 14535
rect 27663 14532 27675 14535
rect 27982 14532 27988 14544
rect 27663 14504 27988 14532
rect 27663 14501 27675 14504
rect 27617 14495 27675 14501
rect 27982 14492 27988 14504
rect 28040 14492 28046 14544
rect 29825 14535 29883 14541
rect 29825 14501 29837 14535
rect 29871 14532 29883 14535
rect 29871 14504 30144 14532
rect 29871 14501 29883 14504
rect 29825 14495 29883 14501
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 25869 14467 25927 14473
rect 25869 14464 25881 14467
rect 24912 14436 25881 14464
rect 24912 14424 24918 14436
rect 25869 14433 25881 14436
rect 25915 14464 25927 14467
rect 27706 14464 27712 14476
rect 25915 14436 27712 14464
rect 25915 14433 25927 14436
rect 25869 14427 25927 14433
rect 27706 14424 27712 14436
rect 27764 14424 27770 14476
rect 26142 14288 26148 14340
rect 26200 14288 26206 14340
rect 29086 14328 29092 14340
rect 27370 14300 29092 14328
rect 24762 14220 24768 14272
rect 24820 14260 24826 14272
rect 27448 14260 27476 14300
rect 29086 14288 29092 14300
rect 29144 14288 29150 14340
rect 30116 14328 30144 14504
rect 30282 14492 30288 14544
rect 30340 14492 30346 14544
rect 32677 14535 32735 14541
rect 32677 14501 32689 14535
rect 32723 14532 32735 14535
rect 34422 14532 34428 14544
rect 32723 14504 34428 14532
rect 32723 14501 32735 14504
rect 32677 14495 32735 14501
rect 34422 14492 34428 14504
rect 34480 14492 34486 14544
rect 37185 14535 37243 14541
rect 37185 14501 37197 14535
rect 37231 14532 37243 14535
rect 39758 14532 39764 14544
rect 37231 14504 39764 14532
rect 37231 14501 37243 14504
rect 37185 14495 37243 14501
rect 39758 14492 39764 14504
rect 39816 14492 39822 14544
rect 30300 14464 30328 14492
rect 30377 14467 30435 14473
rect 30377 14464 30389 14467
rect 30300 14436 30389 14464
rect 30377 14433 30389 14436
rect 30423 14433 30435 14467
rect 30377 14427 30435 14433
rect 32490 14424 32496 14476
rect 32548 14464 32554 14476
rect 33137 14467 33195 14473
rect 33137 14464 33149 14467
rect 32548 14436 33149 14464
rect 32548 14424 32554 14436
rect 33137 14433 33149 14436
rect 33183 14433 33195 14467
rect 33137 14427 33195 14433
rect 33321 14467 33379 14473
rect 33321 14433 33333 14467
rect 33367 14464 33379 14467
rect 33962 14464 33968 14476
rect 33367 14436 33968 14464
rect 33367 14433 33379 14436
rect 33321 14427 33379 14433
rect 33962 14424 33968 14436
rect 34020 14424 34026 14476
rect 35434 14424 35440 14476
rect 35492 14464 35498 14476
rect 37645 14467 37703 14473
rect 37645 14464 37657 14467
rect 35492 14436 37657 14464
rect 35492 14424 35498 14436
rect 37645 14433 37657 14436
rect 37691 14433 37703 14467
rect 37645 14427 37703 14433
rect 37734 14424 37740 14476
rect 37792 14424 37798 14476
rect 30190 14356 30196 14408
rect 30248 14356 30254 14408
rect 30282 14356 30288 14408
rect 30340 14396 30346 14408
rect 33045 14399 33103 14405
rect 33045 14396 33057 14399
rect 30340 14368 33057 14396
rect 30340 14356 30346 14368
rect 33045 14365 33057 14368
rect 33091 14365 33103 14399
rect 33045 14359 33103 14365
rect 34606 14356 34612 14408
rect 34664 14396 34670 14408
rect 34977 14399 35035 14405
rect 34977 14396 34989 14399
rect 34664 14368 34989 14396
rect 34664 14356 34670 14368
rect 34977 14365 34989 14368
rect 35023 14365 35035 14399
rect 34977 14359 35035 14365
rect 37553 14399 37611 14405
rect 37553 14365 37565 14399
rect 37599 14396 37611 14399
rect 38565 14399 38623 14405
rect 38565 14396 38577 14399
rect 37599 14368 38577 14396
rect 37599 14365 37611 14368
rect 37553 14359 37611 14365
rect 38565 14365 38577 14368
rect 38611 14365 38623 14399
rect 38565 14359 38623 14365
rect 39942 14356 39948 14408
rect 40000 14396 40006 14408
rect 40221 14399 40279 14405
rect 40221 14396 40233 14399
rect 40000 14368 40233 14396
rect 40000 14356 40006 14368
rect 40221 14365 40233 14368
rect 40267 14365 40279 14399
rect 40221 14359 40279 14365
rect 30116 14300 34376 14328
rect 24820 14232 27476 14260
rect 24820 14220 24826 14232
rect 28810 14220 28816 14272
rect 28868 14260 28874 14272
rect 30285 14263 30343 14269
rect 30285 14260 30297 14263
rect 28868 14232 30297 14260
rect 28868 14220 28874 14232
rect 30285 14229 30297 14232
rect 30331 14229 30343 14263
rect 34348 14260 34376 14300
rect 35158 14288 35164 14340
rect 35216 14288 35222 14340
rect 36906 14260 36912 14272
rect 34348 14232 36912 14260
rect 30285 14223 30343 14229
rect 36906 14220 36912 14232
rect 36964 14220 36970 14272
rect 40037 14263 40095 14269
rect 40037 14229 40049 14263
rect 40083 14260 40095 14263
rect 44082 14260 44088 14272
rect 40083 14232 44088 14260
rect 40083 14229 40095 14232
rect 40037 14223 40095 14229
rect 44082 14220 44088 14232
rect 44140 14220 44146 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 34790 14056 34796 14068
rect 33980 14028 34796 14056
rect 28997 13991 29055 13997
rect 28997 13957 29009 13991
rect 29043 13988 29055 13991
rect 29270 13988 29276 14000
rect 29043 13960 29276 13988
rect 29043 13957 29055 13960
rect 28997 13951 29055 13957
rect 29270 13948 29276 13960
rect 29328 13948 29334 14000
rect 33980 13988 34008 14028
rect 34790 14016 34796 14028
rect 34848 14056 34854 14068
rect 35802 14056 35808 14068
rect 34848 14028 35808 14056
rect 34848 14016 34854 14028
rect 35802 14016 35808 14028
rect 35860 14016 35866 14068
rect 36725 14059 36783 14065
rect 36725 14025 36737 14059
rect 36771 14056 36783 14059
rect 38562 14056 38568 14068
rect 36771 14028 38568 14056
rect 36771 14025 36783 14028
rect 36725 14019 36783 14025
rect 38562 14016 38568 14028
rect 38620 14016 38626 14068
rect 38933 14059 38991 14065
rect 38933 14025 38945 14059
rect 38979 14056 38991 14059
rect 42702 14056 42708 14068
rect 38979 14028 42708 14056
rect 38979 14025 38991 14028
rect 38933 14019 38991 14025
rect 42702 14016 42708 14028
rect 42760 14016 42766 14068
rect 33888 13960 34008 13988
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 5626 13920 5632 13932
rect 1811 13892 5632 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 30558 13880 30564 13932
rect 30616 13880 30622 13932
rect 33888 13929 33916 13960
rect 36814 13948 36820 14000
rect 36872 13988 36878 14000
rect 37553 13991 37611 13997
rect 37553 13988 37565 13991
rect 36872 13960 37565 13988
rect 36872 13948 36878 13960
rect 37553 13957 37565 13960
rect 37599 13957 37611 13991
rect 37553 13951 37611 13957
rect 37737 13991 37795 13997
rect 37737 13957 37749 13991
rect 37783 13988 37795 13991
rect 40034 13988 40040 14000
rect 37783 13960 40040 13988
rect 37783 13957 37795 13960
rect 37737 13951 37795 13957
rect 40034 13948 40040 13960
rect 40092 13948 40098 14000
rect 33873 13923 33931 13929
rect 33873 13889 33885 13923
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 35250 13880 35256 13932
rect 35308 13880 35314 13932
rect 35452 13892 35756 13920
rect 2774 13812 2780 13864
rect 2832 13812 2838 13864
rect 29181 13855 29239 13861
rect 29181 13821 29193 13855
rect 29227 13852 29239 13855
rect 29730 13852 29736 13864
rect 29227 13824 29736 13852
rect 29227 13821 29239 13824
rect 29181 13815 29239 13821
rect 29730 13812 29736 13824
rect 29788 13812 29794 13864
rect 35452 13852 35480 13892
rect 30392 13824 35480 13852
rect 30392 13793 30420 13824
rect 35526 13812 35532 13864
rect 35584 13852 35590 13864
rect 35621 13855 35679 13861
rect 35621 13852 35633 13855
rect 35584 13824 35633 13852
rect 35584 13812 35590 13824
rect 35621 13821 35633 13824
rect 35667 13821 35679 13855
rect 35728 13852 35756 13892
rect 36906 13880 36912 13932
rect 36964 13880 36970 13932
rect 37826 13880 37832 13932
rect 37884 13920 37890 13932
rect 38289 13923 38347 13929
rect 38289 13920 38301 13923
rect 37884 13892 38301 13920
rect 37884 13880 37890 13892
rect 38289 13889 38301 13892
rect 38335 13889 38347 13923
rect 38289 13883 38347 13889
rect 39114 13880 39120 13932
rect 39172 13880 39178 13932
rect 39482 13880 39488 13932
rect 39540 13920 39546 13932
rect 41969 13923 42027 13929
rect 41969 13920 41981 13923
rect 39540 13892 41981 13920
rect 39540 13880 39546 13892
rect 41969 13889 41981 13892
rect 42015 13889 42027 13923
rect 41969 13883 42027 13889
rect 46658 13880 46664 13932
rect 46716 13920 46722 13932
rect 47949 13923 48007 13929
rect 47949 13920 47961 13923
rect 46716 13892 47961 13920
rect 46716 13880 46722 13892
rect 47949 13889 47961 13892
rect 47995 13889 48007 13923
rect 47949 13883 48007 13889
rect 35728 13824 38332 13852
rect 35621 13815 35679 13821
rect 30377 13787 30435 13793
rect 30377 13753 30389 13787
rect 30423 13753 30435 13787
rect 38304 13784 38332 13824
rect 38378 13812 38384 13864
rect 38436 13852 38442 13864
rect 38473 13855 38531 13861
rect 38473 13852 38485 13855
rect 38436 13824 38485 13852
rect 38436 13812 38442 13824
rect 38473 13821 38485 13824
rect 38519 13821 38531 13855
rect 40678 13852 40684 13864
rect 38473 13815 38531 13821
rect 38580 13824 40684 13852
rect 38580 13784 38608 13824
rect 40678 13812 40684 13824
rect 40736 13812 40742 13864
rect 44358 13852 44364 13864
rect 41800 13824 44364 13852
rect 41800 13793 41828 13824
rect 44358 13812 44364 13824
rect 44416 13812 44422 13864
rect 49142 13812 49148 13864
rect 49200 13812 49206 13864
rect 38304 13756 38608 13784
rect 41785 13787 41843 13793
rect 30377 13747 30435 13753
rect 41785 13753 41797 13787
rect 41831 13753 41843 13787
rect 41785 13747 41843 13753
rect 34136 13719 34194 13725
rect 34136 13685 34148 13719
rect 34182 13716 34194 13719
rect 35434 13716 35440 13728
rect 34182 13688 35440 13716
rect 34182 13685 34194 13688
rect 34136 13679 34194 13685
rect 35434 13676 35440 13688
rect 35492 13676 35498 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 27614 13472 27620 13524
rect 27672 13512 27678 13524
rect 28261 13515 28319 13521
rect 28261 13512 28273 13515
rect 27672 13484 28273 13512
rect 27672 13472 27678 13484
rect 28261 13481 28273 13484
rect 28307 13481 28319 13515
rect 28261 13475 28319 13481
rect 33962 13472 33968 13524
rect 34020 13512 34026 13524
rect 36633 13515 36691 13521
rect 36633 13512 36645 13515
rect 34020 13484 36645 13512
rect 34020 13472 34026 13484
rect 36633 13481 36645 13484
rect 36679 13481 36691 13515
rect 36633 13475 36691 13481
rect 28902 13404 28908 13456
rect 28960 13404 28966 13456
rect 28813 13379 28871 13385
rect 28813 13345 28825 13379
rect 28859 13376 28871 13379
rect 28920 13376 28948 13404
rect 30558 13376 30564 13388
rect 28859 13348 30564 13376
rect 28859 13345 28871 13348
rect 28813 13339 28871 13345
rect 30558 13336 30564 13348
rect 30616 13336 30622 13388
rect 34790 13336 34796 13388
rect 34848 13376 34854 13388
rect 34885 13379 34943 13385
rect 34885 13376 34897 13379
rect 34848 13348 34897 13376
rect 34848 13336 34854 13348
rect 34885 13345 34897 13348
rect 34931 13345 34943 13379
rect 34885 13339 34943 13345
rect 35161 13379 35219 13385
rect 35161 13345 35173 13379
rect 35207 13376 35219 13379
rect 37734 13376 37740 13388
rect 35207 13348 37740 13376
rect 35207 13345 35219 13348
rect 35161 13339 35219 13345
rect 37734 13336 37740 13348
rect 37792 13336 37798 13388
rect 25222 13268 25228 13320
rect 25280 13308 25286 13320
rect 25685 13311 25743 13317
rect 25685 13308 25697 13311
rect 25280 13280 25697 13308
rect 25280 13268 25286 13280
rect 25685 13277 25697 13280
rect 25731 13277 25743 13311
rect 25685 13271 25743 13277
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13308 28779 13311
rect 28902 13308 28908 13320
rect 28767 13280 28908 13308
rect 28767 13277 28779 13280
rect 28721 13271 28779 13277
rect 28902 13268 28908 13280
rect 28960 13308 28966 13320
rect 33686 13308 33692 13320
rect 28960 13280 33692 13308
rect 28960 13268 28966 13280
rect 33686 13268 33692 13280
rect 33744 13268 33750 13320
rect 34146 13268 34152 13320
rect 34204 13268 34210 13320
rect 37182 13268 37188 13320
rect 37240 13268 37246 13320
rect 37366 13268 37372 13320
rect 37424 13308 37430 13320
rect 38105 13311 38163 13317
rect 38105 13308 38117 13311
rect 37424 13280 38117 13308
rect 37424 13268 37430 13280
rect 38105 13277 38117 13280
rect 38151 13277 38163 13311
rect 38105 13271 38163 13277
rect 40678 13268 40684 13320
rect 40736 13268 40742 13320
rect 44542 13268 44548 13320
rect 44600 13308 44606 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 44600 13280 47961 13308
rect 44600 13268 44606 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 28629 13243 28687 13249
rect 28629 13209 28641 13243
rect 28675 13240 28687 13243
rect 36538 13240 36544 13252
rect 28675 13212 31754 13240
rect 36386 13212 36544 13240
rect 28675 13209 28687 13212
rect 28629 13203 28687 13209
rect 31726 13184 31754 13212
rect 36538 13200 36544 13212
rect 36596 13200 36602 13252
rect 49142 13200 49148 13252
rect 49200 13200 49206 13252
rect 24578 13132 24584 13184
rect 24636 13172 24642 13184
rect 25777 13175 25835 13181
rect 25777 13172 25789 13175
rect 24636 13144 25789 13172
rect 24636 13132 24642 13144
rect 25777 13141 25789 13144
rect 25823 13141 25835 13175
rect 31726 13144 31760 13184
rect 25777 13135 25835 13141
rect 31754 13132 31760 13144
rect 31812 13172 31818 13184
rect 32306 13172 32312 13184
rect 31812 13144 32312 13172
rect 31812 13132 31818 13144
rect 32306 13132 32312 13144
rect 32364 13132 32370 13184
rect 34238 13132 34244 13184
rect 34296 13132 34302 13184
rect 37274 13132 37280 13184
rect 37332 13132 37338 13184
rect 37921 13175 37979 13181
rect 37921 13141 37933 13175
rect 37967 13172 37979 13175
rect 39850 13172 39856 13184
rect 37967 13144 39856 13172
rect 37967 13141 37979 13144
rect 37921 13135 37979 13141
rect 39850 13132 39856 13144
rect 39908 13132 39914 13184
rect 40773 13175 40831 13181
rect 40773 13141 40785 13175
rect 40819 13172 40831 13175
rect 46750 13172 46756 13184
rect 40819 13144 46756 13172
rect 40819 13141 40831 13144
rect 40773 13135 40831 13141
rect 46750 13132 46756 13144
rect 46808 13132 46814 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 28718 12928 28724 12980
rect 28776 12968 28782 12980
rect 28813 12971 28871 12977
rect 28813 12968 28825 12971
rect 28776 12940 28825 12968
rect 28776 12928 28782 12940
rect 28813 12937 28825 12940
rect 28859 12937 28871 12971
rect 28813 12931 28871 12937
rect 29270 12928 29276 12980
rect 29328 12968 29334 12980
rect 30282 12968 30288 12980
rect 29328 12940 30288 12968
rect 29328 12928 29334 12940
rect 30282 12928 30288 12940
rect 30340 12928 30346 12980
rect 30466 12928 30472 12980
rect 30524 12968 30530 12980
rect 30650 12968 30656 12980
rect 30524 12940 30656 12968
rect 30524 12928 30530 12940
rect 30650 12928 30656 12940
rect 30708 12928 30714 12980
rect 31938 12928 31944 12980
rect 31996 12968 32002 12980
rect 32306 12968 32312 12980
rect 31996 12940 32312 12968
rect 31996 12928 32002 12940
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 34882 12968 34888 12980
rect 33704 12940 34888 12968
rect 26694 12860 26700 12912
rect 26752 12900 26758 12912
rect 27249 12903 27307 12909
rect 27249 12900 27261 12903
rect 26752 12872 27261 12900
rect 26752 12860 26758 12872
rect 27249 12869 27261 12872
rect 27295 12869 27307 12903
rect 27249 12863 27307 12869
rect 27798 12860 27804 12912
rect 27856 12900 27862 12912
rect 27985 12903 28043 12909
rect 27985 12900 27997 12903
rect 27856 12872 27997 12900
rect 27856 12860 27862 12872
rect 27985 12869 27997 12872
rect 28031 12869 28043 12903
rect 27985 12863 28043 12869
rect 29181 12903 29239 12909
rect 29181 12869 29193 12903
rect 29227 12900 29239 12903
rect 32398 12900 32404 12912
rect 29227 12872 32404 12900
rect 29227 12869 29239 12872
rect 29181 12863 29239 12869
rect 32398 12860 32404 12872
rect 32456 12860 32462 12912
rect 33704 12841 33732 12940
rect 34882 12928 34888 12940
rect 34940 12928 34946 12980
rect 35434 12928 35440 12980
rect 35492 12928 35498 12980
rect 36170 12928 36176 12980
rect 36228 12968 36234 12980
rect 36538 12968 36544 12980
rect 36228 12940 36544 12968
rect 36228 12928 36234 12940
rect 36538 12928 36544 12940
rect 36596 12968 36602 12980
rect 46014 12968 46020 12980
rect 36596 12940 46020 12968
rect 36596 12928 36602 12940
rect 46014 12928 46020 12940
rect 46072 12928 46078 12980
rect 33962 12860 33968 12912
rect 34020 12860 34026 12912
rect 35452 12900 35480 12928
rect 35452 12872 36492 12900
rect 30377 12835 30435 12841
rect 30377 12801 30389 12835
rect 30423 12832 30435 12835
rect 33689 12835 33747 12841
rect 30423 12804 31754 12832
rect 30423 12801 30435 12804
rect 30377 12795 30435 12801
rect 27798 12724 27804 12776
rect 27856 12764 27862 12776
rect 28626 12764 28632 12776
rect 27856 12736 28632 12764
rect 27856 12724 27862 12736
rect 28626 12724 28632 12736
rect 28684 12724 28690 12776
rect 29457 12767 29515 12773
rect 29457 12733 29469 12767
rect 29503 12764 29515 12767
rect 29546 12764 29552 12776
rect 29503 12736 29552 12764
rect 29503 12733 29515 12736
rect 29457 12727 29515 12733
rect 29546 12724 29552 12736
rect 29604 12724 29610 12776
rect 30558 12724 30564 12776
rect 30616 12724 30622 12776
rect 27154 12656 27160 12708
rect 27212 12696 27218 12708
rect 28169 12699 28227 12705
rect 28169 12696 28181 12699
rect 27212 12668 28181 12696
rect 27212 12656 27218 12668
rect 28169 12665 28181 12668
rect 28215 12665 28227 12699
rect 28169 12659 28227 12665
rect 28994 12656 29000 12708
rect 29052 12696 29058 12708
rect 30009 12699 30067 12705
rect 30009 12696 30021 12699
rect 29052 12668 30021 12696
rect 29052 12656 29058 12668
rect 30009 12665 30021 12668
rect 30055 12665 30067 12699
rect 30009 12659 30067 12665
rect 25222 12588 25228 12640
rect 25280 12628 25286 12640
rect 27341 12631 27399 12637
rect 27341 12628 27353 12631
rect 25280 12600 27353 12628
rect 25280 12588 25286 12600
rect 27341 12597 27353 12600
rect 27387 12597 27399 12631
rect 31726 12628 31754 12804
rect 33689 12801 33701 12835
rect 33735 12801 33747 12835
rect 35250 12832 35256 12844
rect 35098 12804 35256 12832
rect 33689 12795 33747 12801
rect 35250 12792 35256 12804
rect 35308 12832 35314 12844
rect 36170 12832 36176 12844
rect 35308 12804 36176 12832
rect 35308 12792 35314 12804
rect 36170 12792 36176 12804
rect 36228 12792 36234 12844
rect 36262 12792 36268 12844
rect 36320 12792 36326 12844
rect 34422 12724 34428 12776
rect 34480 12764 34486 12776
rect 36464 12773 36492 12872
rect 38562 12860 38568 12912
rect 38620 12900 38626 12912
rect 43809 12903 43867 12909
rect 43809 12900 43821 12903
rect 38620 12872 43821 12900
rect 38620 12860 38626 12872
rect 43809 12869 43821 12872
rect 43855 12869 43867 12903
rect 43809 12863 43867 12869
rect 46750 12792 46756 12844
rect 46808 12832 46814 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 46808 12804 47961 12832
rect 46808 12792 46814 12804
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 36357 12767 36415 12773
rect 36357 12764 36369 12767
rect 34480 12736 36369 12764
rect 34480 12724 34486 12736
rect 36357 12733 36369 12736
rect 36403 12733 36415 12767
rect 36357 12727 36415 12733
rect 36449 12767 36507 12773
rect 36449 12733 36461 12767
rect 36495 12733 36507 12767
rect 36449 12727 36507 12733
rect 49142 12724 49148 12776
rect 49200 12724 49206 12776
rect 36538 12696 36544 12708
rect 34992 12668 36544 12696
rect 34992 12628 35020 12668
rect 36538 12656 36544 12668
rect 36596 12656 36602 12708
rect 43993 12699 44051 12705
rect 43993 12665 44005 12699
rect 44039 12696 44051 12699
rect 44726 12696 44732 12708
rect 44039 12668 44732 12696
rect 44039 12665 44051 12668
rect 43993 12659 44051 12665
rect 44726 12656 44732 12668
rect 44784 12656 44790 12708
rect 31726 12600 35020 12628
rect 35897 12631 35955 12637
rect 27341 12591 27399 12597
rect 35897 12597 35909 12631
rect 35943 12628 35955 12631
rect 39942 12628 39948 12640
rect 35943 12600 39948 12628
rect 35943 12597 35955 12600
rect 35897 12591 35955 12597
rect 39942 12588 39948 12600
rect 40000 12588 40006 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 36262 12384 36268 12436
rect 36320 12424 36326 12436
rect 36541 12427 36599 12433
rect 36541 12424 36553 12427
rect 36320 12396 36553 12424
rect 36320 12384 36326 12396
rect 36541 12393 36553 12396
rect 36587 12393 36599 12427
rect 36541 12387 36599 12393
rect 39850 12248 39856 12300
rect 39908 12288 39914 12300
rect 39908 12260 44496 12288
rect 39908 12248 39914 12260
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 9398 12220 9404 12232
rect 3476 12192 9404 12220
rect 3476 12180 3482 12192
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 28813 12223 28871 12229
rect 28813 12189 28825 12223
rect 28859 12220 28871 12223
rect 28902 12220 28908 12232
rect 28859 12192 28908 12220
rect 28859 12189 28871 12192
rect 28813 12183 28871 12189
rect 28902 12180 28908 12192
rect 28960 12180 28966 12232
rect 38286 12180 38292 12232
rect 38344 12220 38350 12232
rect 39025 12223 39083 12229
rect 39025 12220 39037 12223
rect 38344 12192 39037 12220
rect 38344 12180 38350 12192
rect 39025 12189 39037 12192
rect 39071 12189 39083 12223
rect 39025 12183 39083 12189
rect 41322 12180 41328 12232
rect 41380 12220 41386 12232
rect 44468 12229 44496 12260
rect 41417 12223 41475 12229
rect 41417 12220 41429 12223
rect 41380 12192 41429 12220
rect 41380 12180 41386 12192
rect 41417 12189 41429 12192
rect 41463 12189 41475 12223
rect 41417 12183 41475 12189
rect 44453 12223 44511 12229
rect 44453 12189 44465 12223
rect 44499 12189 44511 12223
rect 44453 12183 44511 12189
rect 44726 12180 44732 12232
rect 44784 12220 44790 12232
rect 47949 12223 48007 12229
rect 47949 12220 47961 12223
rect 44784 12192 47961 12220
rect 44784 12180 44790 12192
rect 47949 12189 47961 12192
rect 47995 12189 48007 12223
rect 47949 12183 48007 12189
rect 28997 12155 29055 12161
rect 28997 12121 29009 12155
rect 29043 12152 29055 12155
rect 29178 12152 29184 12164
rect 29043 12124 29184 12152
rect 29043 12121 29055 12124
rect 28997 12115 29055 12121
rect 29178 12112 29184 12124
rect 29236 12112 29242 12164
rect 39209 12155 39267 12161
rect 39209 12121 39221 12155
rect 39255 12152 39267 12155
rect 41874 12152 41880 12164
rect 39255 12124 41880 12152
rect 39255 12121 39267 12124
rect 39209 12115 39267 12121
rect 41874 12112 41880 12124
rect 41932 12112 41938 12164
rect 49142 12112 49148 12164
rect 49200 12112 49206 12164
rect 41233 12087 41291 12093
rect 41233 12053 41245 12087
rect 41279 12084 41291 12087
rect 43346 12084 43352 12096
rect 41279 12056 43352 12084
rect 41279 12053 41291 12056
rect 41233 12047 41291 12053
rect 43346 12044 43352 12056
rect 43404 12044 43410 12096
rect 44266 12044 44272 12096
rect 44324 12044 44330 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 44174 11772 44180 11824
rect 44232 11812 44238 11824
rect 46201 11815 46259 11821
rect 46201 11812 46213 11815
rect 44232 11784 46213 11812
rect 44232 11772 44238 11784
rect 46201 11781 46213 11784
rect 46247 11781 46259 11815
rect 46201 11775 46259 11781
rect 39758 11704 39764 11756
rect 39816 11744 39822 11756
rect 41693 11747 41751 11753
rect 41693 11744 41705 11747
rect 39816 11716 41705 11744
rect 39816 11704 39822 11716
rect 41693 11713 41705 11716
rect 41739 11713 41751 11747
rect 41693 11707 41751 11713
rect 42702 11704 42708 11756
rect 42760 11744 42766 11756
rect 44729 11747 44787 11753
rect 44729 11744 44741 11747
rect 42760 11716 44741 11744
rect 42760 11704 42766 11716
rect 44729 11713 44741 11716
rect 44775 11713 44787 11747
rect 45465 11747 45523 11753
rect 45465 11744 45477 11747
rect 44729 11707 44787 11713
rect 44836 11716 45477 11744
rect 44082 11636 44088 11688
rect 44140 11676 44146 11688
rect 44836 11676 44864 11716
rect 45465 11713 45477 11716
rect 45511 11713 45523 11747
rect 45465 11707 45523 11713
rect 44140 11648 44864 11676
rect 44913 11679 44971 11685
rect 44140 11636 44146 11648
rect 44913 11645 44925 11679
rect 44959 11676 44971 11679
rect 46750 11676 46756 11688
rect 44959 11648 46756 11676
rect 44959 11645 44971 11648
rect 44913 11639 44971 11645
rect 46750 11636 46756 11648
rect 46808 11636 46814 11688
rect 45649 11611 45707 11617
rect 45649 11577 45661 11611
rect 45695 11608 45707 11611
rect 46658 11608 46664 11620
rect 45695 11580 46664 11608
rect 45695 11577 45707 11580
rect 45649 11571 45707 11577
rect 46658 11568 46664 11580
rect 46716 11568 46722 11620
rect 41509 11543 41567 11549
rect 41509 11509 41521 11543
rect 41555 11540 41567 11543
rect 44174 11540 44180 11552
rect 41555 11512 44180 11540
rect 41555 11509 41567 11512
rect 41509 11503 41567 11509
rect 44174 11500 44180 11512
rect 44232 11500 44238 11552
rect 46290 11500 46296 11552
rect 46348 11500 46354 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 17034 11336 17040 11348
rect 13035 11308 17040 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 19794 11200 19800 11212
rect 13679 11172 19800 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13403 11104 14473 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 44266 11092 44272 11144
rect 44324 11132 44330 11144
rect 47949 11135 48007 11141
rect 47949 11132 47961 11135
rect 44324 11104 47961 11132
rect 44324 11092 44330 11104
rect 47949 11101 47961 11104
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 49142 11092 49148 11144
rect 49200 11092 49206 11144
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 12437 11067 12495 11073
rect 12437 11064 12449 11067
rect 7616 11036 12449 11064
rect 7616 11024 7622 11036
rect 12437 11033 12449 11036
rect 12483 11064 12495 11067
rect 13449 11067 13507 11073
rect 13449 11064 13461 11067
rect 12483 11036 13461 11064
rect 12483 11033 12495 11036
rect 12437 11027 12495 11033
rect 13449 11033 13461 11036
rect 13495 11033 13507 11067
rect 13449 11027 13507 11033
rect 44358 11024 44364 11076
rect 44416 11064 44422 11076
rect 46293 11067 46351 11073
rect 46293 11064 46305 11067
rect 44416 11036 46305 11064
rect 44416 11024 44422 11036
rect 46293 11033 46305 11036
rect 46339 11033 46351 11067
rect 46293 11027 46351 11033
rect 46474 11024 46480 11076
rect 46532 11024 46538 11076
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 24302 10684 24308 10736
rect 24360 10724 24366 10736
rect 24397 10727 24455 10733
rect 24397 10724 24409 10727
rect 24360 10696 24409 10724
rect 24360 10684 24366 10696
rect 24397 10693 24409 10696
rect 24443 10693 24455 10727
rect 24397 10687 24455 10693
rect 39942 10616 39948 10668
rect 40000 10656 40006 10668
rect 40865 10659 40923 10665
rect 40865 10656 40877 10659
rect 40000 10628 40877 10656
rect 40000 10616 40006 10628
rect 40865 10625 40877 10628
rect 40911 10625 40923 10659
rect 40865 10619 40923 10625
rect 47762 10616 47768 10668
rect 47820 10656 47826 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 47820 10628 47961 10656
rect 47820 10616 47826 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 49142 10548 49148 10600
rect 49200 10548 49206 10600
rect 24581 10523 24639 10529
rect 24581 10489 24593 10523
rect 24627 10520 24639 10523
rect 25130 10520 25136 10532
rect 24627 10492 25136 10520
rect 24627 10489 24639 10492
rect 24581 10483 24639 10489
rect 25130 10480 25136 10492
rect 25188 10480 25194 10532
rect 40681 10455 40739 10461
rect 40681 10421 40693 10455
rect 40727 10452 40739 10455
rect 42702 10452 42708 10464
rect 40727 10424 42708 10452
rect 40727 10421 40739 10424
rect 40681 10415 40739 10421
rect 42702 10412 42708 10424
rect 42760 10412 42766 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 28442 10004 28448 10056
rect 28500 10044 28506 10056
rect 28721 10047 28779 10053
rect 28721 10044 28733 10047
rect 28500 10016 28733 10044
rect 28500 10004 28506 10016
rect 28721 10013 28733 10016
rect 28767 10013 28779 10047
rect 28721 10007 28779 10013
rect 31846 10004 31852 10056
rect 31904 10004 31910 10056
rect 46750 10004 46756 10056
rect 46808 10044 46814 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 46808 10016 47961 10044
rect 46808 10004 46814 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 28905 9979 28963 9985
rect 28905 9945 28917 9979
rect 28951 9976 28963 9979
rect 30098 9976 30104 9988
rect 28951 9948 30104 9976
rect 28951 9945 28963 9948
rect 28905 9939 28963 9945
rect 30098 9936 30104 9948
rect 30156 9936 30162 9988
rect 49142 9936 49148 9988
rect 49200 9936 49206 9988
rect 29914 9868 29920 9920
rect 29972 9908 29978 9920
rect 31941 9911 31999 9917
rect 31941 9908 31953 9911
rect 29972 9880 31953 9908
rect 29972 9868 29978 9880
rect 31941 9877 31953 9880
rect 31987 9877 31999 9911
rect 31941 9871 31999 9877
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 32030 9596 32036 9648
rect 32088 9636 32094 9648
rect 32401 9639 32459 9645
rect 32401 9636 32413 9639
rect 32088 9608 32413 9636
rect 32088 9596 32094 9608
rect 32401 9605 32413 9608
rect 32447 9605 32459 9639
rect 32401 9599 32459 9605
rect 34974 9596 34980 9648
rect 35032 9636 35038 9648
rect 35989 9639 36047 9645
rect 35989 9636 36001 9639
rect 35032 9608 36001 9636
rect 35032 9596 35038 9608
rect 35989 9605 36001 9608
rect 36035 9605 36047 9639
rect 35989 9599 36047 9605
rect 44174 9528 44180 9580
rect 44232 9568 44238 9580
rect 46201 9571 46259 9577
rect 46201 9568 46213 9571
rect 44232 9540 46213 9568
rect 44232 9528 44238 9540
rect 46201 9537 46213 9540
rect 46247 9537 46259 9571
rect 46201 9531 46259 9537
rect 46658 9528 46664 9580
rect 46716 9568 46722 9580
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 46716 9540 47961 9568
rect 46716 9528 46722 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 49142 9460 49148 9512
rect 49200 9460 49206 9512
rect 32585 9435 32643 9441
rect 32585 9401 32597 9435
rect 32631 9432 32643 9435
rect 33962 9432 33968 9444
rect 32631 9404 33968 9432
rect 32631 9401 32643 9404
rect 32585 9395 32643 9401
rect 33962 9392 33968 9404
rect 34020 9392 34026 9444
rect 36173 9435 36231 9441
rect 36173 9401 36185 9435
rect 36219 9432 36231 9435
rect 37366 9432 37372 9444
rect 36219 9404 37372 9432
rect 36219 9401 36231 9404
rect 36173 9395 36231 9401
rect 37366 9392 37372 9404
rect 37424 9392 37430 9444
rect 46017 9367 46075 9373
rect 46017 9333 46029 9367
rect 46063 9364 46075 9367
rect 47854 9364 47860 9376
rect 46063 9336 47860 9364
rect 46063 9333 46075 9336
rect 46017 9327 46075 9333
rect 47854 9324 47860 9336
rect 47912 9324 47918 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 9582 9092 9588 9104
rect 3384 9064 9588 9092
rect 3384 9052 3390 9064
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 43346 8916 43352 8968
rect 43404 8956 43410 8968
rect 46017 8959 46075 8965
rect 46017 8956 46029 8959
rect 43404 8928 46029 8956
rect 43404 8916 43410 8928
rect 46017 8925 46029 8928
rect 46063 8925 46075 8959
rect 46017 8919 46075 8925
rect 46198 8848 46204 8900
rect 46256 8848 46262 8900
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 9140 8588 13676 8616
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 5592 8520 6914 8548
rect 5592 8508 5598 8520
rect 6886 8412 6914 8520
rect 9140 8489 9168 8588
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 13648 8480 13676 8588
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 19242 8548 19248 8560
rect 16540 8520 19248 8548
rect 16540 8508 16546 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 32306 8508 32312 8560
rect 32364 8548 32370 8560
rect 36541 8551 36599 8557
rect 36541 8548 36553 8551
rect 32364 8520 36553 8548
rect 32364 8508 32370 8520
rect 36541 8517 36553 8520
rect 36587 8517 36599 8551
rect 36541 8511 36599 8517
rect 37921 8551 37979 8557
rect 37921 8517 37933 8551
rect 37967 8548 37979 8551
rect 38470 8548 38476 8560
rect 37967 8520 38476 8548
rect 37967 8517 37979 8520
rect 37921 8511 37979 8517
rect 38470 8508 38476 8520
rect 38528 8508 38534 8560
rect 42702 8508 42708 8560
rect 42760 8548 42766 8560
rect 45741 8551 45799 8557
rect 45741 8548 45753 8551
rect 42760 8520 45753 8548
rect 42760 8508 42766 8520
rect 45741 8517 45753 8520
rect 45787 8517 45799 8551
rect 45741 8511 45799 8517
rect 18598 8480 18604 8492
rect 9125 8443 9183 8449
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 6886 8384 9413 8412
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 10520 8344 10548 8466
rect 13648 8452 18604 8480
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 46474 8440 46480 8492
rect 46532 8480 46538 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 46532 8452 47961 8480
rect 46532 8440 46538 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 21542 8412 21548 8424
rect 11195 8384 21548 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 36725 8415 36783 8421
rect 36725 8381 36737 8415
rect 36771 8412 36783 8415
rect 42610 8412 42616 8424
rect 36771 8384 42616 8412
rect 36771 8381 36783 8384
rect 36725 8375 36783 8381
rect 42610 8372 42616 8384
rect 42668 8372 42674 8424
rect 49142 8372 49148 8424
rect 49200 8372 49206 8424
rect 16482 8344 16488 8356
rect 10520 8316 16488 8344
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 37642 8304 37648 8356
rect 37700 8344 37706 8356
rect 38105 8347 38163 8353
rect 38105 8344 38117 8347
rect 37700 8316 38117 8344
rect 37700 8304 37706 8316
rect 38105 8313 38117 8316
rect 38151 8313 38163 8347
rect 38105 8307 38163 8313
rect 45922 8304 45928 8356
rect 45980 8304 45986 8356
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 46290 7828 46296 7880
rect 46348 7868 46354 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 46348 7840 47961 7868
rect 46348 7828 46354 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 49142 7760 49148 7812
rect 49200 7760 49206 7812
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 31754 7420 31760 7472
rect 31812 7460 31818 7472
rect 35805 7463 35863 7469
rect 35805 7460 35817 7463
rect 31812 7432 35817 7460
rect 31812 7420 31818 7432
rect 35805 7429 35817 7432
rect 35851 7429 35863 7463
rect 35805 7423 35863 7429
rect 29362 7352 29368 7404
rect 29420 7392 29426 7404
rect 37553 7395 37611 7401
rect 37553 7392 37565 7395
rect 29420 7364 37565 7392
rect 29420 7352 29426 7364
rect 37553 7361 37565 7364
rect 37599 7361 37611 7395
rect 37553 7355 37611 7361
rect 47854 7352 47860 7404
rect 47912 7392 47918 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 47912 7364 47961 7392
rect 47912 7352 47918 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 49142 7284 49148 7336
rect 49200 7284 49206 7336
rect 37737 7259 37795 7265
rect 37737 7225 37749 7259
rect 37783 7256 37795 7259
rect 45186 7256 45192 7268
rect 37783 7228 45192 7256
rect 37783 7225 37795 7228
rect 37737 7219 37795 7225
rect 45186 7216 45192 7228
rect 45244 7216 45250 7268
rect 35897 7191 35955 7197
rect 35897 7157 35909 7191
rect 35943 7188 35955 7191
rect 41414 7188 41420 7200
rect 35943 7160 41420 7188
rect 35943 7157 35955 7160
rect 35897 7151 35955 7157
rect 41414 7148 41420 7160
rect 41472 7148 41478 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 8938 6848 8944 6860
rect 3476 6820 8944 6848
rect 3476 6808 3482 6820
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 45922 6808 45928 6860
rect 45980 6848 45986 6860
rect 45980 6820 47992 6848
rect 45980 6808 45986 6820
rect 36538 6740 36544 6792
rect 36596 6780 36602 6792
rect 37737 6783 37795 6789
rect 36596 6752 37688 6780
rect 36596 6740 36602 6752
rect 32398 6672 32404 6724
rect 32456 6712 32462 6724
rect 37553 6715 37611 6721
rect 37553 6712 37565 6715
rect 32456 6684 37565 6712
rect 32456 6672 32462 6684
rect 37553 6681 37565 6684
rect 37599 6681 37611 6715
rect 37660 6712 37688 6752
rect 37737 6749 37749 6783
rect 37783 6780 37795 6783
rect 40126 6780 40132 6792
rect 37783 6752 40132 6780
rect 37783 6749 37795 6752
rect 37737 6743 37795 6749
rect 40126 6740 40132 6752
rect 40184 6740 40190 6792
rect 47394 6740 47400 6792
rect 47452 6740 47458 6792
rect 47964 6789 47992 6820
rect 47949 6783 48007 6789
rect 47949 6749 47961 6783
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 38289 6715 38347 6721
rect 38289 6712 38301 6715
rect 37660 6684 38301 6712
rect 37553 6675 37611 6681
rect 38289 6681 38301 6684
rect 38335 6681 38347 6715
rect 38289 6675 38347 6681
rect 38473 6715 38531 6721
rect 38473 6681 38485 6715
rect 38519 6712 38531 6715
rect 44450 6712 44456 6724
rect 38519 6684 44456 6712
rect 38519 6681 38531 6684
rect 38473 6675 38531 6681
rect 44450 6672 44456 6684
rect 44508 6672 44514 6724
rect 49142 6672 49148 6724
rect 49200 6672 49206 6724
rect 47213 6647 47271 6653
rect 47213 6613 47225 6647
rect 47259 6644 47271 6647
rect 47486 6644 47492 6656
rect 47259 6616 47492 6644
rect 47259 6613 47271 6616
rect 47213 6607 47271 6613
rect 47486 6604 47492 6616
rect 47544 6604 47550 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 48685 6307 48743 6313
rect 48685 6273 48697 6307
rect 48731 6304 48743 6307
rect 48774 6304 48780 6316
rect 48731 6276 48780 6304
rect 48731 6273 48743 6276
rect 48685 6267 48743 6273
rect 48774 6264 48780 6276
rect 48832 6264 48838 6316
rect 48314 6060 48320 6112
rect 48372 6100 48378 6112
rect 48777 6103 48835 6109
rect 48777 6100 48789 6103
rect 48372 6072 48789 6100
rect 48372 6060 48378 6072
rect 48777 6069 48789 6072
rect 48823 6069 48835 6103
rect 48777 6063 48835 6069
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 46198 5652 46204 5704
rect 46256 5692 46262 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 46256 5664 47961 5692
rect 46256 5652 46262 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 49142 5652 49148 5704
rect 49200 5652 49206 5704
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 29457 5219 29515 5225
rect 29457 5216 29469 5219
rect 10100 5188 29469 5216
rect 10100 5176 10106 5188
rect 29457 5185 29469 5188
rect 29503 5216 29515 5219
rect 30101 5219 30159 5225
rect 30101 5216 30113 5219
rect 29503 5188 30113 5216
rect 29503 5185 29515 5188
rect 29457 5179 29515 5185
rect 30101 5185 30113 5188
rect 30147 5185 30159 5219
rect 30101 5179 30159 5185
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 9030 5012 9036 5024
rect 3476 4984 9036 5012
rect 3476 4972 3482 4984
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 30193 5015 30251 5021
rect 30193 4981 30205 5015
rect 30239 5012 30251 5015
rect 47854 5012 47860 5024
rect 30239 4984 47860 5012
rect 30239 4981 30251 4984
rect 30193 4975 30251 4981
rect 47854 4972 47860 4984
rect 47912 4972 47918 5024
rect 49326 4972 49332 5024
rect 49384 4972 49390 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 24670 4564 24676 4616
rect 24728 4604 24734 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 24728 4576 47961 4604
rect 24728 4564 24734 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 49142 4496 49148 4548
rect 49200 4496 49206 4548
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 33962 4088 33968 4140
rect 34020 4088 34026 4140
rect 38378 4088 38384 4140
rect 38436 4128 38442 4140
rect 39117 4131 39175 4137
rect 39117 4128 39129 4131
rect 38436 4100 39129 4128
rect 38436 4088 38442 4100
rect 39117 4097 39129 4100
rect 39163 4097 39175 4131
rect 39117 4091 39175 4097
rect 40126 4088 40132 4140
rect 40184 4128 40190 4140
rect 43533 4131 43591 4137
rect 43533 4128 43545 4131
rect 40184 4100 43545 4128
rect 40184 4088 40190 4100
rect 43533 4097 43545 4100
rect 43579 4097 43591 4131
rect 43533 4091 43591 4097
rect 46014 4088 46020 4140
rect 46072 4088 46078 4140
rect 48774 4088 48780 4140
rect 48832 4088 48838 4140
rect 33870 4020 33876 4072
rect 33928 4060 33934 4072
rect 34425 4063 34483 4069
rect 34425 4060 34437 4063
rect 33928 4032 34437 4060
rect 33928 4020 33934 4032
rect 34425 4029 34437 4032
rect 34471 4029 34483 4063
rect 34425 4023 34483 4029
rect 39022 4020 39028 4072
rect 39080 4060 39086 4072
rect 39577 4063 39635 4069
rect 39577 4060 39589 4063
rect 39080 4032 39589 4060
rect 39080 4020 39086 4032
rect 39577 4029 39589 4032
rect 39623 4029 39635 4063
rect 39577 4023 39635 4029
rect 43438 4020 43444 4072
rect 43496 4060 43502 4072
rect 43993 4063 44051 4069
rect 43993 4060 44005 4063
rect 43496 4032 44005 4060
rect 43496 4020 43502 4032
rect 43993 4029 44005 4032
rect 44039 4029 44051 4063
rect 43993 4023 44051 4029
rect 48501 4063 48559 4069
rect 48501 4029 48513 4063
rect 48547 4060 48559 4063
rect 48590 4060 48596 4072
rect 48547 4032 48596 4060
rect 48547 4029 48559 4032
rect 48501 4023 48559 4029
rect 48590 4020 48596 4032
rect 48648 4020 48654 4072
rect 45833 3927 45891 3933
rect 45833 3893 45845 3927
rect 45879 3924 45891 3927
rect 47762 3924 47768 3936
rect 45879 3896 47768 3924
rect 45879 3893 45891 3896
rect 45833 3887 45891 3893
rect 47762 3884 47768 3896
rect 47820 3884 47826 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 5534 3720 5540 3732
rect 1627 3692 5540 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 25041 3587 25099 3593
rect 25041 3584 25053 3587
rect 24360 3556 25053 3584
rect 24360 3544 24366 3556
rect 25041 3553 25053 3556
rect 25087 3553 25099 3587
rect 25041 3547 25099 3553
rect 29454 3544 29460 3596
rect 29512 3584 29518 3596
rect 30193 3587 30251 3593
rect 30193 3584 30205 3587
rect 29512 3556 30205 3584
rect 29512 3544 29518 3556
rect 30193 3553 30205 3556
rect 30239 3553 30251 3587
rect 30193 3547 30251 3553
rect 30926 3544 30932 3596
rect 30984 3584 30990 3596
rect 32033 3587 32091 3593
rect 32033 3584 32045 3587
rect 30984 3556 32045 3584
rect 30984 3544 30990 3556
rect 32033 3553 32045 3556
rect 32079 3553 32091 3587
rect 32033 3547 32091 3553
rect 34606 3544 34612 3596
rect 34664 3584 34670 3596
rect 35345 3587 35403 3593
rect 35345 3584 35357 3587
rect 34664 3556 35357 3584
rect 34664 3544 34670 3556
rect 35345 3553 35357 3556
rect 35391 3553 35403 3587
rect 35345 3547 35403 3553
rect 36078 3544 36084 3596
rect 36136 3584 36142 3596
rect 37185 3587 37243 3593
rect 37185 3584 37197 3587
rect 36136 3556 37197 3584
rect 36136 3544 36142 3556
rect 37185 3553 37197 3556
rect 37231 3553 37243 3587
rect 37185 3547 37243 3553
rect 39758 3544 39764 3596
rect 39816 3584 39822 3596
rect 40497 3587 40555 3593
rect 40497 3584 40509 3587
rect 39816 3556 40509 3584
rect 39816 3544 39822 3556
rect 40497 3553 40509 3556
rect 40543 3553 40555 3587
rect 40497 3547 40555 3553
rect 41230 3544 41236 3596
rect 41288 3584 41294 3596
rect 42337 3587 42395 3593
rect 42337 3584 42349 3587
rect 41288 3556 42349 3584
rect 41288 3544 41294 3556
rect 42337 3553 42349 3556
rect 42383 3553 42395 3587
rect 42337 3547 42395 3553
rect 44174 3544 44180 3596
rect 44232 3584 44238 3596
rect 45649 3587 45707 3593
rect 45649 3584 45661 3587
rect 44232 3556 45661 3584
rect 44232 3544 44238 3556
rect 45649 3553 45661 3556
rect 45695 3553 45707 3587
rect 45649 3547 45707 3553
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3516 1823 3519
rect 2774 3516 2780 3528
rect 1811 3488 2780 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 24578 3476 24584 3528
rect 24636 3476 24642 3528
rect 29730 3476 29736 3528
rect 29788 3476 29794 3528
rect 30098 3476 30104 3528
rect 30156 3516 30162 3528
rect 31573 3519 31631 3525
rect 31573 3516 31585 3519
rect 30156 3488 31585 3516
rect 30156 3476 30162 3488
rect 31573 3485 31585 3488
rect 31619 3485 31631 3519
rect 31573 3479 31631 3485
rect 34238 3476 34244 3528
rect 34296 3516 34302 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34296 3488 34897 3516
rect 34296 3476 34302 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 36722 3476 36728 3528
rect 36780 3476 36786 3528
rect 37366 3476 37372 3528
rect 37424 3516 37430 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 37424 3488 40049 3516
rect 37424 3476 37430 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 41874 3476 41880 3528
rect 41932 3476 41938 3528
rect 45186 3476 45192 3528
rect 45244 3476 45250 3528
rect 48133 3519 48191 3525
rect 48133 3485 48145 3519
rect 48179 3516 48191 3519
rect 48314 3516 48320 3528
rect 48179 3488 48320 3516
rect 48179 3485 48191 3488
rect 48133 3479 48191 3485
rect 48314 3476 48320 3488
rect 48372 3476 48378 3528
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 21358 3448 21364 3460
rect 6972 3420 21364 3448
rect 6972 3408 6978 3420
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 49145 3451 49203 3457
rect 49145 3417 49157 3451
rect 49191 3448 49203 3451
rect 49326 3448 49332 3460
rect 49191 3420 49332 3448
rect 49191 3417 49203 3420
rect 49145 3411 49203 3417
rect 49326 3408 49332 3420
rect 49384 3408 49390 3460
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 27246 3380 27252 3392
rect 12860 3352 27252 3380
rect 12860 3340 12866 3352
rect 27246 3340 27252 3352
rect 27304 3340 27310 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 12802 3136 12808 3188
rect 12860 3136 12866 3188
rect 14277 3179 14335 3185
rect 14277 3145 14289 3179
rect 14323 3176 14335 3179
rect 17218 3176 17224 3188
rect 14323 3148 17224 3176
rect 14323 3145 14335 3148
rect 14277 3139 14335 3145
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 17954 3136 17960 3188
rect 18012 3136 18018 3188
rect 28350 3176 28356 3188
rect 20824 3148 28356 3176
rect 4065 3111 4123 3117
rect 4065 3077 4077 3111
rect 4111 3108 4123 3111
rect 19978 3108 19984 3120
rect 4111 3080 19984 3108
rect 4111 3077 4123 3080
rect 4065 3071 4123 3077
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1544 3012 1593 3040
rect 1544 3000 1550 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1581 3003 1639 3009
rect 1688 3012 2513 3040
rect 750 2932 756 2984
rect 808 2972 814 2984
rect 1688 2972 1716 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3752 3012 3893 3040
rect 3752 3000 3758 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5224 3012 5273 3040
rect 5224 3000 5230 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6696 3012 6837 3040
rect 6696 3000 6702 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10376 3012 10425 3040
rect 10376 3000 10382 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 12584 3012 12725 3040
rect 12584 3000 12590 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14093 3043 14151 3049
rect 14093 3040 14105 3043
rect 14056 3012 14105 3040
rect 14056 3000 14062 3012
rect 14093 3009 14105 3012
rect 14139 3009 14151 3043
rect 14093 3003 14151 3009
rect 17678 3000 17684 3052
rect 17736 3040 17742 3052
rect 17773 3043 17831 3049
rect 17773 3040 17785 3043
rect 17736 3012 17785 3040
rect 17736 3000 17742 3012
rect 17773 3009 17785 3012
rect 17819 3009 17831 3043
rect 17773 3003 17831 3009
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3040 19579 3043
rect 20824 3040 20852 3148
rect 28350 3136 28356 3148
rect 28408 3136 28414 3188
rect 27430 3108 27436 3120
rect 20916 3080 22232 3108
rect 20916 3049 20944 3080
rect 19567 3012 20852 3040
rect 20901 3043 20959 3049
rect 19567 3009 19579 3012
rect 19521 3003 19579 3009
rect 20901 3009 20913 3043
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 17310 2972 17316 2984
rect 808 2944 1716 2972
rect 1780 2944 17316 2972
rect 808 2932 814 2944
rect 1780 2913 1808 2944
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 19150 2932 19156 2984
rect 19208 2972 19214 2984
rect 19245 2975 19303 2981
rect 19245 2972 19257 2975
rect 19208 2944 19257 2972
rect 19208 2932 19214 2944
rect 19245 2941 19257 2944
rect 19291 2941 19303 2975
rect 19245 2935 19303 2941
rect 20622 2932 20628 2984
rect 20680 2932 20686 2984
rect 22005 2975 22063 2981
rect 22005 2941 22017 2975
rect 22051 2972 22063 2975
rect 22094 2972 22100 2984
rect 22051 2944 22100 2972
rect 22051 2941 22063 2944
rect 22005 2935 22063 2941
rect 22094 2932 22100 2944
rect 22152 2932 22158 2984
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2873 1823 2907
rect 1765 2867 1823 2873
rect 2317 2907 2375 2913
rect 2317 2873 2329 2907
rect 2363 2904 2375 2907
rect 2363 2876 4660 2904
rect 2363 2873 2375 2876
rect 2317 2867 2375 2873
rect 4632 2836 4660 2876
rect 5442 2864 5448 2916
rect 5500 2864 5506 2916
rect 7558 2904 7564 2916
rect 6886 2876 7564 2904
rect 6886 2836 6914 2876
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 10597 2907 10655 2913
rect 10597 2873 10609 2907
rect 10643 2904 10655 2907
rect 14458 2904 14464 2916
rect 10643 2876 14464 2904
rect 10643 2873 10655 2876
rect 10597 2867 10655 2873
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 22204 2904 22232 3080
rect 22296 3080 27436 3108
rect 22296 3049 22324 3080
rect 27430 3068 27436 3080
rect 27488 3068 27494 3120
rect 37274 3068 37280 3120
rect 37332 3108 37338 3120
rect 37332 3080 39344 3108
rect 37332 3068 37338 3080
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3009 22339 3043
rect 22281 3003 22339 3009
rect 23385 3043 23443 3049
rect 23385 3009 23397 3043
rect 23431 3040 23443 3043
rect 24118 3040 24124 3052
rect 23431 3012 24124 3040
rect 23431 3009 23443 3012
rect 23385 3003 23443 3009
rect 24118 3000 24124 3012
rect 24176 3000 24182 3052
rect 25130 3000 25136 3052
rect 25188 3000 25194 3052
rect 27338 3000 27344 3052
rect 27396 3000 27402 3052
rect 29178 3000 29184 3052
rect 29236 3000 29242 3052
rect 32493 3043 32551 3049
rect 32493 3009 32505 3043
rect 32539 3040 32551 3043
rect 33318 3040 33324 3052
rect 32539 3012 33324 3040
rect 32539 3009 32551 3012
rect 32493 3003 32551 3009
rect 33318 3000 33324 3012
rect 33376 3000 33382 3052
rect 34330 3000 34336 3052
rect 34388 3000 34394 3052
rect 37642 3000 37648 3052
rect 37700 3000 37706 3052
rect 39316 3049 39344 3080
rect 39301 3043 39359 3049
rect 39301 3009 39313 3043
rect 39347 3009 39359 3043
rect 39301 3003 39359 3009
rect 42610 3000 42616 3052
rect 42668 3000 42674 3052
rect 44450 3000 44456 3052
rect 44508 3000 44514 3052
rect 46661 3043 46719 3049
rect 46661 3009 46673 3043
rect 46707 3040 46719 3043
rect 47394 3040 47400 3052
rect 46707 3012 47400 3040
rect 46707 3009 46719 3012
rect 46661 3003 46719 3009
rect 47394 3000 47400 3012
rect 47452 3000 47458 3052
rect 47486 3000 47492 3052
rect 47544 3040 47550 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47544 3012 47961 3040
rect 47544 3000 47550 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23753 2975 23811 2981
rect 23753 2972 23765 2975
rect 23624 2944 23765 2972
rect 23624 2932 23630 2944
rect 23753 2941 23765 2944
rect 23799 2941 23811 2975
rect 23753 2935 23811 2941
rect 25038 2932 25044 2984
rect 25096 2972 25102 2984
rect 25593 2975 25651 2981
rect 25593 2972 25605 2975
rect 25096 2944 25605 2972
rect 25096 2932 25102 2944
rect 25593 2941 25605 2944
rect 25639 2941 25651 2975
rect 25593 2935 25651 2941
rect 27246 2932 27252 2984
rect 27304 2972 27310 2984
rect 27801 2975 27859 2981
rect 27801 2972 27813 2975
rect 27304 2944 27813 2972
rect 27304 2932 27310 2944
rect 27801 2941 27813 2944
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 29641 2975 29699 2981
rect 29641 2972 29653 2975
rect 28776 2944 29653 2972
rect 28776 2932 28782 2944
rect 29641 2941 29653 2944
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 31662 2932 31668 2984
rect 31720 2972 31726 2984
rect 32769 2975 32827 2981
rect 32769 2972 32781 2975
rect 31720 2944 32781 2972
rect 31720 2932 31726 2944
rect 32769 2941 32781 2944
rect 32815 2941 32827 2975
rect 32769 2935 32827 2941
rect 34609 2975 34667 2981
rect 34609 2941 34621 2975
rect 34655 2941 34667 2975
rect 34609 2935 34667 2941
rect 30466 2904 30472 2916
rect 22204 2876 30472 2904
rect 30466 2864 30472 2876
rect 30524 2864 30530 2916
rect 32398 2864 32404 2916
rect 32456 2904 32462 2916
rect 34624 2904 34652 2935
rect 36814 2932 36820 2984
rect 36872 2972 36878 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 36872 2944 37933 2972
rect 36872 2932 36878 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 39761 2975 39819 2981
rect 39761 2941 39773 2975
rect 39807 2941 39819 2975
rect 39761 2935 39819 2941
rect 32456 2876 34652 2904
rect 32456 2864 32462 2876
rect 37550 2864 37556 2916
rect 37608 2904 37614 2916
rect 39776 2904 39804 2935
rect 41966 2932 41972 2984
rect 42024 2972 42030 2984
rect 43073 2975 43131 2981
rect 43073 2972 43085 2975
rect 42024 2944 43085 2972
rect 42024 2932 42030 2944
rect 43073 2941 43085 2944
rect 43119 2941 43131 2975
rect 43073 2935 43131 2941
rect 44913 2975 44971 2981
rect 44913 2941 44925 2975
rect 44959 2941 44971 2975
rect 44913 2935 44971 2941
rect 46385 2975 46443 2981
rect 46385 2941 46397 2975
rect 46431 2972 46443 2975
rect 47118 2972 47124 2984
rect 46431 2944 47124 2972
rect 46431 2941 46443 2944
rect 46385 2935 46443 2941
rect 37608 2876 39804 2904
rect 37608 2864 37614 2876
rect 42702 2864 42708 2916
rect 42760 2904 42766 2916
rect 44928 2904 44956 2935
rect 47118 2932 47124 2944
rect 47176 2932 47182 2984
rect 47854 2932 47860 2984
rect 47912 2972 47918 2984
rect 48409 2975 48467 2981
rect 48409 2972 48421 2975
rect 47912 2944 48421 2972
rect 47912 2932 47918 2944
rect 48409 2941 48421 2944
rect 48455 2941 48467 2975
rect 48409 2935 48467 2941
rect 42760 2876 44956 2904
rect 42760 2864 42766 2876
rect 4632 2808 6914 2836
rect 46382 2796 46388 2848
rect 46440 2836 46446 2848
rect 48314 2836 48320 2848
rect 46440 2808 48320 2836
rect 46440 2796 46446 2808
rect 48314 2796 48320 2808
rect 48372 2796 48378 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 7561 2635 7619 2641
rect 7561 2601 7573 2635
rect 7607 2632 7619 2635
rect 14458 2632 14464 2644
rect 7607 2604 14464 2632
rect 7607 2601 7619 2604
rect 7561 2595 7619 2601
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 14553 2635 14611 2641
rect 14553 2601 14565 2635
rect 14599 2632 14611 2635
rect 18690 2632 18696 2644
rect 14599 2604 18696 2632
rect 14599 2601 14611 2604
rect 14553 2595 14611 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 20714 2632 20720 2644
rect 18800 2604 20720 2632
rect 9493 2567 9551 2573
rect 9493 2533 9505 2567
rect 9539 2564 9551 2567
rect 9539 2536 16528 2564
rect 9539 2533 9551 2536
rect 9493 2527 9551 2533
rect 4893 2499 4951 2505
rect 4893 2465 4905 2499
rect 4939 2496 4951 2499
rect 16390 2496 16396 2508
rect 4939 2468 16396 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2222 2428 2228 2440
rect 2179 2400 2228 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 7374 2428 7380 2440
rect 7331 2400 7380 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8619 2400 9536 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 3053 2363 3111 2369
rect 3053 2360 3065 2363
rect 3016 2332 3065 2360
rect 3016 2320 3022 2332
rect 3053 2329 3065 2332
rect 3099 2329 3111 2363
rect 3053 2323 3111 2329
rect 4430 2320 4436 2372
rect 4488 2360 4494 2372
rect 4617 2363 4675 2369
rect 4617 2360 4629 2363
rect 4488 2332 4629 2360
rect 4488 2320 4494 2332
rect 4617 2329 4629 2332
rect 4663 2329 4675 2363
rect 4617 2323 4675 2329
rect 5629 2363 5687 2369
rect 5629 2329 5641 2363
rect 5675 2360 5687 2363
rect 5902 2360 5908 2372
rect 5675 2332 5908 2360
rect 5675 2329 5687 2332
rect 5629 2323 5687 2329
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 5994 2320 6000 2372
rect 6052 2320 6058 2372
rect 7834 2320 7840 2372
rect 7892 2360 7898 2372
rect 8205 2363 8263 2369
rect 8205 2360 8217 2363
rect 7892 2332 8217 2360
rect 7892 2320 7898 2332
rect 8205 2329 8217 2332
rect 8251 2329 8263 2363
rect 8205 2323 8263 2329
rect 8846 2320 8852 2372
rect 8904 2360 8910 2372
rect 9217 2363 9275 2369
rect 9217 2360 9229 2363
rect 8904 2332 9229 2360
rect 8904 2320 8910 2332
rect 9217 2329 9229 2332
rect 9263 2329 9275 2363
rect 9508 2360 9536 2400
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 9640 2400 10241 2428
rect 9640 2388 9646 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 12342 2388 12348 2440
rect 12400 2388 12406 2440
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 14734 2428 14740 2440
rect 14415 2400 14740 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14734 2388 14740 2400
rect 14792 2388 14798 2440
rect 16500 2428 16528 2536
rect 16574 2524 16580 2576
rect 16632 2564 16638 2576
rect 18800 2564 18828 2604
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 20806 2592 20812 2644
rect 20864 2632 20870 2644
rect 22186 2632 22192 2644
rect 20864 2604 22192 2632
rect 20864 2592 20870 2604
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 46014 2592 46020 2644
rect 46072 2632 46078 2644
rect 46753 2635 46811 2641
rect 46753 2632 46765 2635
rect 46072 2604 46765 2632
rect 46072 2592 46078 2604
rect 46753 2601 46765 2604
rect 46799 2601 46811 2635
rect 46753 2595 46811 2601
rect 16632 2536 18828 2564
rect 20073 2567 20131 2573
rect 16632 2524 16638 2536
rect 20073 2533 20085 2567
rect 20119 2564 20131 2567
rect 27798 2564 27804 2576
rect 20119 2536 27804 2564
rect 20119 2533 20131 2536
rect 20073 2527 20131 2533
rect 27798 2524 27804 2536
rect 27856 2524 27862 2576
rect 18049 2499 18107 2505
rect 18049 2465 18061 2499
rect 18095 2496 18107 2499
rect 18414 2496 18420 2508
rect 18095 2468 18420 2496
rect 18095 2465 18107 2468
rect 18049 2459 18107 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 21358 2496 21364 2508
rect 20671 2468 21364 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 21358 2456 21364 2468
rect 21416 2456 21422 2508
rect 22830 2456 22836 2508
rect 22888 2496 22894 2508
rect 23109 2499 23167 2505
rect 23109 2496 23121 2499
rect 22888 2468 23121 2496
rect 22888 2456 22894 2468
rect 23109 2465 23121 2468
rect 23155 2465 23167 2499
rect 23109 2459 23167 2465
rect 25774 2456 25780 2508
rect 25832 2456 25838 2508
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26568 2468 27629 2496
rect 26568 2456 26574 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 28350 2456 28356 2508
rect 28408 2496 28414 2508
rect 30193 2499 30251 2505
rect 30193 2496 30205 2499
rect 28408 2468 30205 2496
rect 28408 2456 28414 2468
rect 30193 2465 30205 2468
rect 30239 2465 30251 2499
rect 30193 2459 30251 2465
rect 30282 2456 30288 2508
rect 30340 2496 30346 2508
rect 32769 2499 32827 2505
rect 32769 2496 32781 2499
rect 30340 2468 32781 2496
rect 30340 2456 30346 2468
rect 32769 2465 32781 2468
rect 32815 2465 32827 2499
rect 32769 2459 32827 2465
rect 35342 2456 35348 2508
rect 35400 2496 35406 2508
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 35400 2468 37933 2496
rect 35400 2456 35406 2468
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 38286 2456 38292 2508
rect 38344 2496 38350 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 38344 2468 40509 2496
rect 38344 2456 38350 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 40586 2456 40592 2508
rect 40644 2496 40650 2508
rect 43073 2499 43131 2505
rect 43073 2496 43085 2499
rect 40644 2468 43085 2496
rect 40644 2456 40650 2468
rect 43073 2465 43085 2468
rect 43119 2465 43131 2499
rect 43073 2459 43131 2465
rect 48314 2456 48320 2508
rect 48372 2456 48378 2508
rect 14844 2400 15608 2428
rect 16500 2400 17264 2428
rect 10781 2363 10839 2369
rect 9508 2332 10732 2360
rect 9217 2323 9275 2329
rect 2406 2252 2412 2304
rect 2464 2252 2470 2304
rect 3326 2252 3332 2304
rect 3384 2252 3390 2304
rect 10042 2252 10048 2304
rect 10100 2252 10106 2304
rect 10704 2292 10732 2332
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 11054 2360 11060 2372
rect 10827 2332 11060 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 11146 2320 11152 2372
rect 11204 2320 11210 2372
rect 11790 2320 11796 2372
rect 11848 2360 11854 2372
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 11848 2332 11989 2360
rect 11848 2320 11854 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 13262 2320 13268 2372
rect 13320 2360 13326 2372
rect 13357 2363 13415 2369
rect 13357 2360 13369 2363
rect 13320 2332 13369 2360
rect 13320 2320 13326 2332
rect 13357 2329 13369 2332
rect 13403 2329 13415 2363
rect 14844 2360 14872 2400
rect 13357 2323 13415 2329
rect 13556 2332 14872 2360
rect 15197 2363 15255 2369
rect 13556 2292 13584 2332
rect 15197 2329 15209 2363
rect 15243 2360 15255 2363
rect 15470 2360 15476 2372
rect 15243 2332 15476 2360
rect 15243 2329 15255 2332
rect 15197 2323 15255 2329
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 10704 2264 13584 2292
rect 13630 2252 13636 2304
rect 13688 2252 13694 2304
rect 15286 2252 15292 2304
rect 15344 2252 15350 2304
rect 15580 2292 15608 2400
rect 15933 2363 15991 2369
rect 15933 2329 15945 2363
rect 15979 2360 15991 2363
rect 16206 2360 16212 2372
rect 15979 2332 16212 2360
rect 15979 2329 15991 2332
rect 15933 2323 15991 2329
rect 16206 2320 16212 2332
rect 16264 2320 16270 2372
rect 16298 2320 16304 2372
rect 16356 2320 16362 2372
rect 16942 2320 16948 2372
rect 17000 2360 17006 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 17000 2332 17141 2360
rect 17000 2320 17006 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17236 2360 17264 2400
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 18322 2388 18328 2440
rect 18380 2388 18386 2440
rect 19797 2431 19855 2437
rect 19797 2397 19809 2431
rect 19843 2428 19855 2431
rect 19886 2428 19892 2440
rect 19843 2400 19892 2428
rect 19843 2397 19855 2400
rect 19797 2391 19855 2397
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 20898 2388 20904 2440
rect 20956 2388 20962 2440
rect 22646 2388 22652 2440
rect 22704 2388 22710 2440
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 29914 2388 29920 2440
rect 29972 2388 29978 2440
rect 31018 2388 31024 2440
rect 31076 2428 31082 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31076 2400 32321 2428
rect 31076 2388 31082 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 33836 2400 34897 2428
rect 33836 2388 33842 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35250 2388 35256 2440
rect 35308 2428 35314 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 35308 2400 37473 2428
rect 35308 2388 35314 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 40034 2388 40040 2440
rect 40092 2388 40098 2440
rect 41414 2388 41420 2440
rect 41472 2428 41478 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 41472 2400 42625 2428
rect 41472 2388 41478 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 47762 2388 47768 2440
rect 47820 2388 47826 2440
rect 23658 2360 23664 2372
rect 17236 2332 23664 2360
rect 17129 2323 17187 2329
rect 23658 2320 23664 2332
rect 23716 2320 23722 2372
rect 35805 2363 35863 2369
rect 35805 2329 35817 2363
rect 35851 2329 35863 2363
rect 35805 2323 35863 2329
rect 45465 2363 45523 2369
rect 45465 2329 45477 2363
rect 45511 2360 45523 2363
rect 45646 2360 45652 2372
rect 45511 2332 45652 2360
rect 45511 2329 45523 2332
rect 45465 2323 45523 2329
rect 20806 2292 20812 2304
rect 15580 2264 20812 2292
rect 20806 2252 20812 2264
rect 20864 2252 20870 2304
rect 20990 2252 20996 2304
rect 21048 2292 21054 2304
rect 23750 2292 23756 2304
rect 21048 2264 23756 2292
rect 21048 2252 21054 2264
rect 23750 2252 23756 2264
rect 23808 2252 23814 2304
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 35820 2292 35848 2323
rect 45646 2320 45652 2332
rect 45704 2320 45710 2372
rect 33192 2264 35848 2292
rect 33192 2252 33198 2264
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
rect 13630 2048 13636 2100
rect 13688 2088 13694 2100
rect 22554 2088 22560 2100
rect 13688 2060 22560 2088
rect 13688 2048 13694 2060
rect 22554 2048 22560 2060
rect 22612 2048 22618 2100
rect 14458 1980 14464 2032
rect 14516 2020 14522 2032
rect 20990 2020 20996 2032
rect 14516 1992 20996 2020
rect 14516 1980 14522 1992
rect 20990 1980 20996 1992
rect 21048 1980 21054 2032
rect 16298 1912 16304 1964
rect 16356 1952 16362 1964
rect 28534 1952 28540 1964
rect 16356 1924 28540 1952
rect 16356 1912 16362 1924
rect 28534 1912 28540 1924
rect 28592 1912 28598 1964
rect 18322 1844 18328 1896
rect 18380 1884 18386 1896
rect 28810 1884 28816 1896
rect 18380 1856 28816 1884
rect 18380 1844 18386 1856
rect 28810 1844 28816 1856
rect 28868 1844 28874 1896
rect 2406 1776 2412 1828
rect 2464 1816 2470 1828
rect 19518 1816 19524 1828
rect 2464 1788 19524 1816
rect 2464 1776 2470 1788
rect 19518 1776 19524 1788
rect 19576 1776 19582 1828
rect 20898 1776 20904 1828
rect 20956 1816 20962 1828
rect 29270 1816 29276 1828
rect 20956 1788 29276 1816
rect 20956 1776 20962 1788
rect 29270 1776 29276 1788
rect 29328 1776 29334 1828
rect 3326 1708 3332 1760
rect 3384 1748 3390 1760
rect 21082 1748 21088 1760
rect 3384 1720 21088 1748
rect 3384 1708 3390 1720
rect 21082 1708 21088 1720
rect 21140 1708 21146 1760
rect 17494 1640 17500 1692
rect 17552 1680 17558 1692
rect 26050 1680 26056 1692
rect 17552 1652 26056 1680
rect 17552 1640 17558 1652
rect 26050 1640 26056 1652
rect 26108 1640 26114 1692
<< via1 >>
rect 388 55700 440 55752
rect 2872 55700 2924 55752
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 27950 54374 28002 54426
rect 28014 54374 28066 54426
rect 28078 54374 28130 54426
rect 28142 54374 28194 54426
rect 28206 54374 28258 54426
rect 37950 54374 38002 54426
rect 38014 54374 38066 54426
rect 38078 54374 38130 54426
rect 38142 54374 38194 54426
rect 38206 54374 38258 54426
rect 47950 54374 48002 54426
rect 48014 54374 48066 54426
rect 48078 54374 48130 54426
rect 48142 54374 48194 54426
rect 48206 54374 48258 54426
rect 3332 54204 3384 54256
rect 2780 54136 2832 54188
rect 10048 54272 10100 54324
rect 28908 54272 28960 54324
rect 37740 54272 37792 54324
rect 6276 54204 6328 54256
rect 8484 54204 8536 54256
rect 11428 54204 11480 54256
rect 13636 54204 13688 54256
rect 16580 54204 16632 54256
rect 18788 54204 18840 54256
rect 20996 54247 21048 54256
rect 20996 54213 21005 54247
rect 21005 54213 21039 54247
rect 21039 54213 21048 54247
rect 20996 54204 21048 54213
rect 24676 54204 24728 54256
rect 28356 54204 28408 54256
rect 32772 54204 32824 54256
rect 33508 54204 33560 54256
rect 37188 54204 37240 54256
rect 42340 54204 42392 54256
rect 3976 53975 4028 53984
rect 3976 53941 3985 53975
rect 3985 53941 4019 53975
rect 4019 53941 4028 53975
rect 3976 53932 4028 53941
rect 11704 54136 11756 54188
rect 14556 54136 14608 54188
rect 17684 54179 17736 54188
rect 17684 54145 17693 54179
rect 17693 54145 17727 54179
rect 17727 54145 17736 54179
rect 17684 54136 17736 54145
rect 20352 54136 20404 54188
rect 22744 54179 22796 54188
rect 22744 54145 22753 54179
rect 22753 54145 22787 54179
rect 22787 54145 22796 54179
rect 22744 54136 22796 54145
rect 25412 54136 25464 54188
rect 26240 54136 26292 54188
rect 26884 54136 26936 54188
rect 27620 54136 27672 54188
rect 29828 54136 29880 54188
rect 30564 54136 30616 54188
rect 31300 54136 31352 54188
rect 34244 54136 34296 54188
rect 35716 54136 35768 54188
rect 36452 54136 36504 54188
rect 38660 54136 38712 54188
rect 39396 54136 39448 54188
rect 40132 54136 40184 54188
rect 40868 54136 40920 54188
rect 43076 54136 43128 54188
rect 44088 54136 44140 54188
rect 44548 54136 44600 54188
rect 47860 54136 47912 54188
rect 20168 54068 20220 54120
rect 22468 54068 22520 54120
rect 43996 54068 44048 54120
rect 48228 54068 48280 54120
rect 14648 54000 14700 54052
rect 25228 54000 25280 54052
rect 29644 54000 29696 54052
rect 33416 54000 33468 54052
rect 33968 54000 34020 54052
rect 40316 54000 40368 54052
rect 12348 53932 12400 53984
rect 26056 53932 26108 53984
rect 26240 53975 26292 53984
rect 26240 53941 26249 53975
rect 26249 53941 26283 53975
rect 26283 53941 26292 53975
rect 26240 53932 26292 53941
rect 27436 53932 27488 53984
rect 28540 53932 28592 53984
rect 30104 53975 30156 53984
rect 30104 53941 30113 53975
rect 30113 53941 30147 53975
rect 30147 53941 30156 53975
rect 30104 53932 30156 53941
rect 30472 53932 30524 53984
rect 35256 53932 35308 53984
rect 36544 53932 36596 53984
rect 37188 53932 37240 53984
rect 37648 53975 37700 53984
rect 37648 53941 37657 53975
rect 37657 53941 37691 53975
rect 37691 53941 37700 53975
rect 37648 53932 37700 53941
rect 38936 53975 38988 53984
rect 38936 53941 38945 53975
rect 38945 53941 38979 53975
rect 38979 53941 38988 53975
rect 38936 53932 38988 53941
rect 40408 53932 40460 53984
rect 41052 53932 41104 53984
rect 43444 54000 43496 54052
rect 45192 53975 45244 53984
rect 45192 53941 45201 53975
rect 45201 53941 45235 53975
rect 45235 53941 45244 53975
rect 45192 53932 45244 53941
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 32950 53830 33002 53882
rect 33014 53830 33066 53882
rect 33078 53830 33130 53882
rect 33142 53830 33194 53882
rect 33206 53830 33258 53882
rect 42950 53830 43002 53882
rect 43014 53830 43066 53882
rect 43078 53830 43130 53882
rect 43142 53830 43194 53882
rect 43206 53830 43258 53882
rect 15844 53660 15896 53712
rect 27068 53660 27120 53712
rect 1860 53592 1912 53644
rect 5540 53592 5592 53644
rect 7012 53592 7064 53644
rect 10692 53592 10744 53644
rect 12164 53592 12216 53644
rect 18328 53635 18380 53644
rect 18328 53601 18337 53635
rect 18337 53601 18371 53635
rect 18371 53601 18380 53635
rect 18328 53592 18380 53601
rect 20260 53592 20312 53644
rect 21732 53592 21784 53644
rect 46756 53592 46808 53644
rect 6276 53456 6328 53508
rect 8944 53524 8996 53576
rect 10416 53567 10468 53576
rect 10416 53533 10425 53567
rect 10425 53533 10459 53567
rect 10459 53533 10468 53567
rect 10416 53524 10468 53533
rect 14740 53524 14792 53576
rect 10784 53456 10836 53508
rect 18420 53524 18472 53576
rect 22836 53524 22888 53576
rect 23296 53524 23348 53576
rect 23940 53524 23992 53576
rect 29092 53524 29144 53576
rect 32036 53524 32088 53576
rect 34980 53524 35032 53576
rect 37832 53524 37884 53576
rect 41604 53524 41656 53576
rect 46204 53524 46256 53576
rect 22192 53456 22244 53508
rect 25780 53456 25832 53508
rect 20444 53388 20496 53440
rect 29736 53431 29788 53440
rect 29736 53397 29745 53431
rect 29745 53397 29779 53431
rect 29779 53397 29788 53431
rect 29736 53388 29788 53397
rect 32128 53431 32180 53440
rect 32128 53397 32137 53431
rect 32137 53397 32171 53431
rect 32171 53397 32180 53431
rect 32128 53388 32180 53397
rect 35348 53388 35400 53440
rect 37832 53388 37884 53440
rect 40684 53388 40736 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 27950 53286 28002 53338
rect 28014 53286 28066 53338
rect 28078 53286 28130 53338
rect 28142 53286 28194 53338
rect 28206 53286 28258 53338
rect 37950 53286 38002 53338
rect 38014 53286 38066 53338
rect 38078 53286 38130 53338
rect 38142 53286 38194 53338
rect 38206 53286 38258 53338
rect 47950 53286 48002 53338
rect 48014 53286 48066 53338
rect 48078 53286 48130 53338
rect 48142 53286 48194 53338
rect 48206 53286 48258 53338
rect 46204 53227 46256 53236
rect 46204 53193 46213 53227
rect 46213 53193 46247 53227
rect 46247 53193 46256 53227
rect 46204 53184 46256 53193
rect 940 53048 992 53100
rect 6368 53116 6420 53168
rect 9864 53116 9916 53168
rect 9036 53048 9088 53100
rect 9772 53091 9824 53100
rect 9772 53057 9781 53091
rect 9781 53057 9815 53091
rect 9815 53057 9824 53091
rect 9772 53048 9824 53057
rect 16948 53116 17000 53168
rect 15200 53048 15252 53100
rect 21272 53116 21324 53168
rect 49700 53116 49752 53168
rect 19616 53091 19668 53100
rect 19616 53057 19625 53091
rect 19625 53057 19659 53091
rect 19659 53057 19668 53091
rect 19616 53048 19668 53057
rect 46388 53091 46440 53100
rect 46388 53057 46397 53091
rect 46397 53057 46431 53091
rect 46431 53057 46440 53091
rect 46388 53048 46440 53057
rect 47676 53048 47728 53100
rect 2596 52980 2648 53032
rect 4896 52980 4948 53032
rect 7748 52980 7800 53032
rect 9956 52980 10008 53032
rect 12808 52980 12860 53032
rect 15108 52980 15160 53032
rect 17316 52980 17368 53032
rect 19524 52980 19576 53032
rect 1952 52912 2004 52964
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 32950 52742 33002 52794
rect 33014 52742 33066 52794
rect 33078 52742 33130 52794
rect 33142 52742 33194 52794
rect 33206 52742 33258 52794
rect 42950 52742 43002 52794
rect 43014 52742 43066 52794
rect 43078 52742 43130 52794
rect 43142 52742 43194 52794
rect 43206 52742 43258 52794
rect 1124 52504 1176 52556
rect 5816 52572 5868 52624
rect 4068 52504 4120 52556
rect 9220 52504 9272 52556
rect 14372 52504 14424 52556
rect 9128 52436 9180 52488
rect 14464 52436 14516 52488
rect 19156 52436 19208 52488
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 27950 52198 28002 52250
rect 28014 52198 28066 52250
rect 28078 52198 28130 52250
rect 28142 52198 28194 52250
rect 28206 52198 28258 52250
rect 37950 52198 38002 52250
rect 38014 52198 38066 52250
rect 38078 52198 38130 52250
rect 38142 52198 38194 52250
rect 38206 52198 38258 52250
rect 47950 52198 48002 52250
rect 48014 52198 48066 52250
rect 48078 52198 48130 52250
rect 48142 52198 48194 52250
rect 48206 52198 48258 52250
rect 22744 52096 22796 52148
rect 2872 52028 2924 52080
rect 1584 52003 1636 52012
rect 1584 51969 1593 52003
rect 1593 51969 1627 52003
rect 1627 51969 1636 52003
rect 1584 51960 1636 51969
rect 23756 52003 23808 52012
rect 23756 51969 23765 52003
rect 23765 51969 23799 52003
rect 23799 51969 23808 52003
rect 23756 51960 23808 51969
rect 49056 52003 49108 52012
rect 49056 51969 49065 52003
rect 49065 51969 49099 52003
rect 49099 51969 49108 52003
rect 49056 51960 49108 51969
rect 49240 51799 49292 51808
rect 49240 51765 49249 51799
rect 49249 51765 49283 51799
rect 49283 51765 49292 51799
rect 49240 51756 49292 51765
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 32950 51654 33002 51706
rect 33014 51654 33066 51706
rect 33078 51654 33130 51706
rect 33142 51654 33194 51706
rect 33206 51654 33258 51706
rect 42950 51654 43002 51706
rect 43014 51654 43066 51706
rect 43078 51654 43130 51706
rect 43142 51654 43194 51706
rect 43206 51654 43258 51706
rect 10048 51552 10100 51604
rect 14464 51595 14516 51604
rect 14464 51561 14473 51595
rect 14473 51561 14507 51595
rect 14507 51561 14516 51595
rect 14464 51552 14516 51561
rect 22836 51552 22888 51604
rect 26700 51348 26752 51400
rect 49056 51391 49108 51400
rect 49056 51357 49065 51391
rect 49065 51357 49099 51391
rect 49099 51357 49108 51391
rect 49056 51348 49108 51357
rect 14280 51280 14332 51332
rect 15936 51280 15988 51332
rect 49148 51212 49200 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 27950 51110 28002 51162
rect 28014 51110 28066 51162
rect 28078 51110 28130 51162
rect 28142 51110 28194 51162
rect 28206 51110 28258 51162
rect 37950 51110 38002 51162
rect 38014 51110 38066 51162
rect 38078 51110 38130 51162
rect 38142 51110 38194 51162
rect 38206 51110 38258 51162
rect 47950 51110 48002 51162
rect 48014 51110 48066 51162
rect 48078 51110 48130 51162
rect 48142 51110 48194 51162
rect 48206 51110 48258 51162
rect 22192 51051 22244 51060
rect 22192 51017 22201 51051
rect 22201 51017 22235 51051
rect 22235 51017 22244 51051
rect 22192 51008 22244 51017
rect 20352 50940 20404 50992
rect 940 50872 992 50924
rect 22744 50872 22796 50924
rect 24124 50872 24176 50924
rect 48964 50915 49016 50924
rect 48964 50881 48973 50915
rect 48973 50881 49007 50915
rect 49007 50881 49016 50915
rect 48964 50872 49016 50881
rect 1676 50668 1728 50720
rect 49424 50668 49476 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 32950 50566 33002 50618
rect 33014 50566 33066 50618
rect 33078 50566 33130 50618
rect 33142 50566 33194 50618
rect 33206 50566 33258 50618
rect 42950 50566 43002 50618
rect 43014 50566 43066 50618
rect 43078 50566 43130 50618
rect 43142 50566 43194 50618
rect 43206 50566 43258 50618
rect 17684 50464 17736 50516
rect 49056 50303 49108 50312
rect 49056 50269 49065 50303
rect 49065 50269 49099 50303
rect 49099 50269 49108 50303
rect 49056 50260 49108 50269
rect 21824 50192 21876 50244
rect 48412 50124 48464 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 27950 50022 28002 50074
rect 28014 50022 28066 50074
rect 28078 50022 28130 50074
rect 28142 50022 28194 50074
rect 28206 50022 28258 50074
rect 37950 50022 38002 50074
rect 38014 50022 38066 50074
rect 38078 50022 38130 50074
rect 38142 50022 38194 50074
rect 38206 50022 38258 50074
rect 47950 50022 48002 50074
rect 48014 50022 48066 50074
rect 48078 50022 48130 50074
rect 48142 50022 48194 50074
rect 48206 50022 48258 50074
rect 12348 49963 12400 49972
rect 12348 49929 12357 49963
rect 12357 49929 12391 49963
rect 12391 49929 12400 49963
rect 12348 49920 12400 49929
rect 14740 49963 14792 49972
rect 14740 49929 14749 49963
rect 14749 49929 14783 49963
rect 14783 49929 14792 49963
rect 14740 49920 14792 49929
rect 20904 49852 20956 49904
rect 16856 49784 16908 49836
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 32950 49478 33002 49530
rect 33014 49478 33066 49530
rect 33078 49478 33130 49530
rect 33142 49478 33194 49530
rect 33206 49478 33258 49530
rect 42950 49478 43002 49530
rect 43014 49478 43066 49530
rect 43078 49478 43130 49530
rect 43142 49478 43194 49530
rect 43206 49478 43258 49530
rect 15200 49376 15252 49428
rect 18420 49376 18472 49428
rect 20720 49172 20772 49224
rect 49056 49215 49108 49224
rect 49056 49181 49065 49215
rect 49065 49181 49099 49215
rect 49099 49181 49108 49215
rect 49056 49172 49108 49181
rect 22100 49104 22152 49156
rect 48872 49036 48924 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 27950 48934 28002 48986
rect 28014 48934 28066 48986
rect 28078 48934 28130 48986
rect 28142 48934 28194 48986
rect 28206 48934 28258 48986
rect 37950 48934 38002 48986
rect 38014 48934 38066 48986
rect 38078 48934 38130 48986
rect 38142 48934 38194 48986
rect 38206 48934 38258 48986
rect 47950 48934 48002 48986
rect 48014 48934 48066 48986
rect 48078 48934 48130 48986
rect 48142 48934 48194 48986
rect 48206 48934 48258 48986
rect 49056 48739 49108 48748
rect 49056 48705 49065 48739
rect 49065 48705 49099 48739
rect 49099 48705 49108 48739
rect 49056 48696 49108 48705
rect 48964 48492 49016 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 32950 48390 33002 48442
rect 33014 48390 33066 48442
rect 33078 48390 33130 48442
rect 33142 48390 33194 48442
rect 33206 48390 33258 48442
rect 42950 48390 43002 48442
rect 43014 48390 43066 48442
rect 43078 48390 43130 48442
rect 43142 48390 43194 48442
rect 43206 48390 43258 48442
rect 21088 48152 21140 48204
rect 49056 48127 49108 48136
rect 49056 48093 49065 48127
rect 49065 48093 49099 48127
rect 49099 48093 49108 48127
rect 49056 48084 49108 48093
rect 940 48016 992 48068
rect 1860 48059 1912 48068
rect 1860 48025 1869 48059
rect 1869 48025 1903 48059
rect 1903 48025 1912 48059
rect 1860 48016 1912 48025
rect 3976 48016 4028 48068
rect 21916 48016 21968 48068
rect 20536 47948 20588 48000
rect 40132 47948 40184 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 27950 47846 28002 47898
rect 28014 47846 28066 47898
rect 28078 47846 28130 47898
rect 28142 47846 28194 47898
rect 28206 47846 28258 47898
rect 37950 47846 38002 47898
rect 38014 47846 38066 47898
rect 38078 47846 38130 47898
rect 38142 47846 38194 47898
rect 38206 47846 38258 47898
rect 47950 47846 48002 47898
rect 48014 47846 48066 47898
rect 48078 47846 48130 47898
rect 48142 47846 48194 47898
rect 48206 47846 48258 47898
rect 23756 47744 23808 47796
rect 25872 47608 25924 47660
rect 49056 47651 49108 47660
rect 49056 47617 49065 47651
rect 49065 47617 49099 47651
rect 49099 47617 49108 47651
rect 49056 47608 49108 47617
rect 48688 47404 48740 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 32950 47302 33002 47354
rect 33014 47302 33066 47354
rect 33078 47302 33130 47354
rect 33142 47302 33194 47354
rect 33206 47302 33258 47354
rect 42950 47302 43002 47354
rect 43014 47302 43066 47354
rect 43078 47302 43130 47354
rect 43142 47302 43194 47354
rect 43206 47302 43258 47354
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 27950 46758 28002 46810
rect 28014 46758 28066 46810
rect 28078 46758 28130 46810
rect 28142 46758 28194 46810
rect 28206 46758 28258 46810
rect 37950 46758 38002 46810
rect 38014 46758 38066 46810
rect 38078 46758 38130 46810
rect 38142 46758 38194 46810
rect 38206 46758 38258 46810
rect 47950 46758 48002 46810
rect 48014 46758 48066 46810
rect 48078 46758 48130 46810
rect 48142 46758 48194 46810
rect 48206 46758 48258 46810
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 32950 46214 33002 46266
rect 33014 46214 33066 46266
rect 33078 46214 33130 46266
rect 33142 46214 33194 46266
rect 33206 46214 33258 46266
rect 42950 46214 43002 46266
rect 43014 46214 43066 46266
rect 43078 46214 43130 46266
rect 43142 46214 43194 46266
rect 43206 46214 43258 46266
rect 15936 46112 15988 46164
rect 26700 46155 26752 46164
rect 26700 46121 26709 46155
rect 26709 46121 26743 46155
rect 26743 46121 26752 46155
rect 26700 46112 26752 46121
rect 940 45840 992 45892
rect 14280 45840 14332 45892
rect 22008 45908 22060 45960
rect 27804 45908 27856 45960
rect 48596 45908 48648 45960
rect 1768 45815 1820 45824
rect 1768 45781 1777 45815
rect 1777 45781 1811 45815
rect 1811 45781 1820 45815
rect 1768 45772 1820 45781
rect 20628 45840 20680 45892
rect 49148 45883 49200 45892
rect 49148 45849 49157 45883
rect 49157 45849 49191 45883
rect 49191 45849 49200 45883
rect 49148 45840 49200 45849
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 27950 45670 28002 45722
rect 28014 45670 28066 45722
rect 28078 45670 28130 45722
rect 28142 45670 28194 45722
rect 28206 45670 28258 45722
rect 37950 45670 38002 45722
rect 38014 45670 38066 45722
rect 38078 45670 38130 45722
rect 38142 45670 38194 45722
rect 38206 45670 38258 45722
rect 47950 45670 48002 45722
rect 48014 45670 48066 45722
rect 48078 45670 48130 45722
rect 48142 45670 48194 45722
rect 48206 45670 48258 45722
rect 1768 45568 1820 45620
rect 22468 45568 22520 45620
rect 48596 45611 48648 45620
rect 48596 45577 48605 45611
rect 48605 45577 48639 45611
rect 48639 45577 48648 45611
rect 48596 45568 48648 45577
rect 10416 45500 10468 45552
rect 32128 45500 32180 45552
rect 46388 45500 46440 45552
rect 21548 45432 21600 45484
rect 29736 45432 29788 45484
rect 33416 45432 33468 45484
rect 48320 45432 48372 45484
rect 32864 45407 32916 45416
rect 32864 45373 32873 45407
rect 32873 45373 32907 45407
rect 32907 45373 32916 45407
rect 32864 45364 32916 45373
rect 33968 45407 34020 45416
rect 33968 45373 33977 45407
rect 33977 45373 34011 45407
rect 34011 45373 34020 45407
rect 33968 45364 34020 45373
rect 34152 45407 34204 45416
rect 34152 45373 34161 45407
rect 34161 45373 34195 45407
rect 34195 45373 34204 45407
rect 34152 45364 34204 45373
rect 32680 45228 32732 45280
rect 33508 45271 33560 45280
rect 33508 45237 33517 45271
rect 33517 45237 33551 45271
rect 33551 45237 33560 45271
rect 33508 45228 33560 45237
rect 46940 45228 46992 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 32950 45126 33002 45178
rect 33014 45126 33066 45178
rect 33078 45126 33130 45178
rect 33142 45126 33194 45178
rect 33206 45126 33258 45178
rect 42950 45126 43002 45178
rect 43014 45126 43066 45178
rect 43078 45126 43130 45178
rect 43142 45126 43194 45178
rect 43206 45126 43258 45178
rect 22744 45024 22796 45076
rect 24124 45024 24176 45076
rect 35992 44956 36044 45008
rect 35348 44931 35400 44940
rect 35348 44897 35357 44931
rect 35357 44897 35391 44931
rect 35391 44897 35400 44931
rect 35348 44888 35400 44897
rect 35532 44931 35584 44940
rect 35532 44897 35541 44931
rect 35541 44897 35575 44931
rect 35575 44897 35584 44931
rect 35532 44888 35584 44897
rect 24492 44820 24544 44872
rect 27160 44820 27212 44872
rect 38384 44820 38436 44872
rect 48504 44863 48556 44872
rect 48504 44829 48513 44863
rect 48513 44829 48547 44863
rect 48547 44829 48556 44863
rect 48504 44820 48556 44829
rect 35256 44727 35308 44736
rect 35256 44693 35265 44727
rect 35265 44693 35299 44727
rect 35299 44693 35308 44727
rect 35256 44684 35308 44693
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 27950 44582 28002 44634
rect 28014 44582 28066 44634
rect 28078 44582 28130 44634
rect 28142 44582 28194 44634
rect 28206 44582 28258 44634
rect 37950 44582 38002 44634
rect 38014 44582 38066 44634
rect 38078 44582 38130 44634
rect 38142 44582 38194 44634
rect 38206 44582 38258 44634
rect 47950 44582 48002 44634
rect 48014 44582 48066 44634
rect 48078 44582 48130 44634
rect 48142 44582 48194 44634
rect 48206 44582 48258 44634
rect 9772 44480 9824 44532
rect 37832 44480 37884 44532
rect 40684 44480 40736 44532
rect 14464 44344 14516 44396
rect 36544 44387 36596 44396
rect 36544 44353 36553 44387
rect 36553 44353 36587 44387
rect 36587 44353 36596 44387
rect 36544 44344 36596 44353
rect 37648 44344 37700 44396
rect 36912 44276 36964 44328
rect 38660 44276 38712 44328
rect 36176 44183 36228 44192
rect 36176 44149 36185 44183
rect 36185 44149 36219 44183
rect 36219 44149 36228 44183
rect 36176 44140 36228 44149
rect 38752 44183 38804 44192
rect 38752 44149 38761 44183
rect 38761 44149 38795 44183
rect 38795 44149 38804 44183
rect 38752 44140 38804 44149
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 32950 44038 33002 44090
rect 33014 44038 33066 44090
rect 33078 44038 33130 44090
rect 33142 44038 33194 44090
rect 33206 44038 33258 44090
rect 42950 44038 43002 44090
rect 43014 44038 43066 44090
rect 43078 44038 43130 44090
rect 43142 44038 43194 44090
rect 43206 44038 43258 44090
rect 11704 43936 11756 43988
rect 14648 43936 14700 43988
rect 16948 43979 17000 43988
rect 16948 43945 16957 43979
rect 16957 43945 16991 43979
rect 16991 43945 17000 43979
rect 16948 43936 17000 43945
rect 20444 43979 20496 43988
rect 20444 43945 20453 43979
rect 20453 43945 20487 43979
rect 20487 43945 20496 43979
rect 20444 43936 20496 43945
rect 21272 43979 21324 43988
rect 21272 43945 21281 43979
rect 21281 43945 21315 43979
rect 21315 43945 21324 43979
rect 21272 43936 21324 43945
rect 21824 43979 21876 43988
rect 21824 43945 21833 43979
rect 21833 43945 21867 43979
rect 21867 43945 21876 43979
rect 21824 43936 21876 43945
rect 32588 43936 32640 43988
rect 9036 43868 9088 43920
rect 19616 43868 19668 43920
rect 22284 43732 22336 43784
rect 12164 43707 12216 43716
rect 12164 43673 12173 43707
rect 12173 43673 12207 43707
rect 12207 43673 12216 43707
rect 12164 43664 12216 43673
rect 13452 43707 13504 43716
rect 13452 43673 13461 43707
rect 13461 43673 13495 43707
rect 13495 43673 13504 43707
rect 13452 43664 13504 43673
rect 16120 43707 16172 43716
rect 16120 43673 16129 43707
rect 16129 43673 16163 43707
rect 16163 43673 16172 43707
rect 16120 43664 16172 43673
rect 17040 43664 17092 43716
rect 21180 43707 21232 43716
rect 21180 43673 21189 43707
rect 21189 43673 21223 43707
rect 21223 43673 21232 43707
rect 21180 43664 21232 43673
rect 22744 43707 22796 43716
rect 22744 43673 22753 43707
rect 22753 43673 22787 43707
rect 22787 43673 22796 43707
rect 22744 43664 22796 43673
rect 28448 43800 28500 43852
rect 32864 43800 32916 43852
rect 37740 43843 37792 43852
rect 37740 43809 37749 43843
rect 37749 43809 37783 43843
rect 37783 43809 37792 43843
rect 37740 43800 37792 43809
rect 38292 43800 38344 43852
rect 26240 43732 26292 43784
rect 28724 43732 28776 43784
rect 32220 43775 32272 43784
rect 32220 43741 32229 43775
rect 32229 43741 32263 43775
rect 32263 43741 32272 43775
rect 32220 43732 32272 43741
rect 40776 43732 40828 43784
rect 48504 43775 48556 43784
rect 48504 43741 48513 43775
rect 48513 43741 48547 43775
rect 48547 43741 48556 43775
rect 48504 43732 48556 43741
rect 31300 43664 31352 43716
rect 27620 43596 27672 43648
rect 28908 43639 28960 43648
rect 28908 43605 28917 43639
rect 28917 43605 28951 43639
rect 28951 43605 28960 43639
rect 28908 43596 28960 43605
rect 31760 43639 31812 43648
rect 31760 43605 31769 43639
rect 31769 43605 31803 43639
rect 31803 43605 31812 43639
rect 31760 43596 31812 43605
rect 33232 43664 33284 43716
rect 37188 43664 37240 43716
rect 33324 43596 33376 43648
rect 37280 43639 37332 43648
rect 37280 43605 37289 43639
rect 37289 43605 37323 43639
rect 37323 43605 37332 43639
rect 37280 43596 37332 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 27950 43494 28002 43546
rect 28014 43494 28066 43546
rect 28078 43494 28130 43546
rect 28142 43494 28194 43546
rect 28206 43494 28258 43546
rect 37950 43494 38002 43546
rect 38014 43494 38066 43546
rect 38078 43494 38130 43546
rect 38142 43494 38194 43546
rect 38206 43494 38258 43546
rect 47950 43494 48002 43546
rect 48014 43494 48066 43546
rect 48078 43494 48130 43546
rect 48142 43494 48194 43546
rect 48206 43494 48258 43546
rect 16856 43435 16908 43444
rect 16856 43401 16865 43435
rect 16865 43401 16899 43435
rect 16899 43401 16908 43435
rect 16856 43392 16908 43401
rect 19156 43435 19208 43444
rect 19156 43401 19165 43435
rect 19165 43401 19199 43435
rect 19199 43401 19208 43435
rect 19156 43392 19208 43401
rect 20352 43435 20404 43444
rect 20352 43401 20361 43435
rect 20361 43401 20395 43435
rect 20395 43401 20404 43435
rect 20352 43392 20404 43401
rect 20904 43435 20956 43444
rect 20904 43401 20913 43435
rect 20913 43401 20947 43435
rect 20947 43401 20956 43435
rect 20904 43392 20956 43401
rect 25872 43435 25924 43444
rect 25872 43401 25881 43435
rect 25881 43401 25915 43435
rect 25915 43401 25924 43435
rect 25872 43392 25924 43401
rect 12164 43324 12216 43376
rect 21916 43324 21968 43376
rect 12072 43299 12124 43308
rect 12072 43265 12081 43299
rect 12081 43265 12115 43299
rect 12115 43265 12124 43299
rect 12072 43256 12124 43265
rect 8944 43188 8996 43240
rect 19064 43299 19116 43308
rect 19064 43265 19073 43299
rect 19073 43265 19107 43299
rect 19107 43265 19116 43299
rect 19064 43256 19116 43265
rect 20260 43299 20312 43308
rect 20260 43265 20269 43299
rect 20269 43265 20303 43299
rect 20303 43265 20312 43299
rect 20260 43256 20312 43265
rect 19432 43188 19484 43240
rect 25964 43256 26016 43308
rect 26332 43231 26384 43240
rect 26332 43197 26341 43231
rect 26341 43197 26375 43231
rect 26375 43197 26384 43231
rect 26332 43188 26384 43197
rect 27344 43188 27396 43240
rect 29184 43324 29236 43376
rect 30380 43324 30432 43376
rect 31300 43324 31352 43376
rect 32220 43256 32272 43308
rect 33232 43324 33284 43376
rect 40316 43435 40368 43444
rect 40316 43401 40325 43435
rect 40325 43401 40359 43435
rect 40359 43401 40368 43435
rect 40316 43392 40368 43401
rect 34796 43367 34848 43376
rect 34796 43333 34805 43367
rect 34805 43333 34839 43367
rect 34839 43333 34848 43367
rect 34796 43324 34848 43333
rect 34520 43299 34572 43308
rect 34520 43265 34529 43299
rect 34529 43265 34563 43299
rect 34563 43265 34572 43299
rect 34520 43256 34572 43265
rect 28724 43188 28776 43240
rect 31944 43188 31996 43240
rect 33232 43188 33284 43240
rect 38936 43256 38988 43308
rect 39764 43256 39816 43308
rect 28448 43052 28500 43104
rect 34152 43120 34204 43172
rect 40500 43231 40552 43240
rect 40500 43197 40509 43231
rect 40509 43197 40543 43231
rect 40543 43197 40552 43231
rect 40500 43188 40552 43197
rect 41604 43188 41656 43240
rect 48504 43231 48556 43240
rect 48504 43197 48513 43231
rect 48513 43197 48547 43231
rect 48547 43197 48556 43231
rect 48504 43188 48556 43197
rect 35900 43120 35952 43172
rect 34060 43095 34112 43104
rect 34060 43061 34069 43095
rect 34069 43061 34103 43095
rect 34103 43061 34112 43095
rect 34060 43052 34112 43061
rect 41236 43052 41288 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 32950 42950 33002 43002
rect 33014 42950 33066 43002
rect 33078 42950 33130 43002
rect 33142 42950 33194 43002
rect 33206 42950 33258 43002
rect 42950 42950 43002 43002
rect 43014 42950 43066 43002
rect 43078 42950 43130 43002
rect 43142 42950 43194 43002
rect 43206 42950 43258 43002
rect 27344 42891 27396 42900
rect 27344 42857 27353 42891
rect 27353 42857 27387 42891
rect 27387 42857 27396 42891
rect 27344 42848 27396 42857
rect 9128 42712 9180 42764
rect 14556 42712 14608 42764
rect 36912 42712 36964 42764
rect 40684 42755 40736 42764
rect 40684 42721 40693 42755
rect 40693 42721 40727 42755
rect 40727 42721 40736 42755
rect 40684 42712 40736 42721
rect 24676 42644 24728 42696
rect 34520 42644 34572 42696
rect 37004 42644 37056 42696
rect 43444 42644 43496 42696
rect 48504 42687 48556 42696
rect 48504 42653 48513 42687
rect 48513 42653 48547 42687
rect 48547 42653 48556 42687
rect 48504 42644 48556 42653
rect 9220 42619 9272 42628
rect 9220 42585 9229 42619
rect 9229 42585 9263 42619
rect 9263 42585 9272 42619
rect 9220 42576 9272 42585
rect 17408 42576 17460 42628
rect 25872 42619 25924 42628
rect 25872 42585 25881 42619
rect 25881 42585 25915 42619
rect 25915 42585 25924 42619
rect 25872 42576 25924 42585
rect 24860 42508 24912 42560
rect 37188 42508 37240 42560
rect 40040 42551 40092 42560
rect 40040 42517 40049 42551
rect 40049 42517 40083 42551
rect 40083 42517 40092 42551
rect 40040 42508 40092 42517
rect 40408 42551 40460 42560
rect 40408 42517 40417 42551
rect 40417 42517 40451 42551
rect 40451 42517 40460 42551
rect 40408 42508 40460 42517
rect 40592 42508 40644 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 27950 42406 28002 42458
rect 28014 42406 28066 42458
rect 28078 42406 28130 42458
rect 28142 42406 28194 42458
rect 28206 42406 28258 42458
rect 37950 42406 38002 42458
rect 38014 42406 38066 42458
rect 38078 42406 38130 42458
rect 38142 42406 38194 42458
rect 38206 42406 38258 42458
rect 47950 42406 48002 42458
rect 48014 42406 48066 42458
rect 48078 42406 48130 42458
rect 48142 42406 48194 42458
rect 48206 42406 48258 42458
rect 6276 42304 6328 42356
rect 20720 42347 20772 42356
rect 20720 42313 20729 42347
rect 20729 42313 20763 42347
rect 20763 42313 20772 42347
rect 20720 42304 20772 42313
rect 22100 42347 22152 42356
rect 22100 42313 22109 42347
rect 22109 42313 22143 42347
rect 22143 42313 22152 42347
rect 22100 42304 22152 42313
rect 6368 42236 6420 42288
rect 7104 42211 7156 42220
rect 7104 42177 7113 42211
rect 7113 42177 7147 42211
rect 7147 42177 7156 42211
rect 7104 42168 7156 42177
rect 7840 42211 7892 42220
rect 7840 42177 7849 42211
rect 7849 42177 7883 42211
rect 7883 42177 7892 42211
rect 7840 42168 7892 42177
rect 20996 42168 21048 42220
rect 22560 42168 22612 42220
rect 24676 42236 24728 42288
rect 24860 42236 24912 42288
rect 27344 42236 27396 42288
rect 30196 42304 30248 42356
rect 29368 42236 29420 42288
rect 31760 42304 31812 42356
rect 32772 42304 32824 42356
rect 34520 42304 34572 42356
rect 38292 42304 38344 42356
rect 45192 42304 45244 42356
rect 31300 42236 31352 42288
rect 35900 42236 35952 42288
rect 37004 42236 37056 42288
rect 39580 42236 39632 42288
rect 41052 42168 41104 42220
rect 41328 42168 41380 42220
rect 24400 42143 24452 42152
rect 24400 42109 24409 42143
rect 24409 42109 24443 42143
rect 24443 42109 24452 42143
rect 24400 42100 24452 42109
rect 27252 42100 27304 42152
rect 28724 42100 28776 42152
rect 29736 42032 29788 42084
rect 35532 42100 35584 42152
rect 37832 42100 37884 42152
rect 39304 42100 39356 42152
rect 41880 42143 41932 42152
rect 41880 42109 41889 42143
rect 41889 42109 41923 42143
rect 41923 42109 41932 42143
rect 41880 42100 41932 42109
rect 48504 42143 48556 42152
rect 48504 42109 48513 42143
rect 48513 42109 48547 42143
rect 48547 42109 48556 42143
rect 48504 42100 48556 42109
rect 39856 42032 39908 42084
rect 20536 41964 20588 42016
rect 22376 41964 22428 42016
rect 24860 41964 24912 42016
rect 25872 42007 25924 42016
rect 25872 41973 25881 42007
rect 25881 41973 25915 42007
rect 25915 41973 25924 42007
rect 25872 41964 25924 41973
rect 29460 42007 29512 42016
rect 29460 41973 29469 42007
rect 29469 41973 29503 42007
rect 29503 41973 29512 42007
rect 29460 41964 29512 41973
rect 31944 41964 31996 42016
rect 34888 41964 34940 42016
rect 42340 41964 42392 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 32950 41862 33002 41914
rect 33014 41862 33066 41914
rect 33078 41862 33130 41914
rect 33142 41862 33194 41914
rect 33206 41862 33258 41914
rect 42950 41862 43002 41914
rect 43014 41862 43066 41914
rect 43078 41862 43130 41914
rect 43142 41862 43194 41914
rect 43206 41862 43258 41914
rect 1584 41760 1636 41812
rect 23664 41760 23716 41812
rect 26332 41760 26384 41812
rect 22928 41692 22980 41744
rect 22652 41624 22704 41676
rect 23664 41667 23716 41676
rect 23664 41633 23673 41667
rect 23673 41633 23707 41667
rect 23707 41633 23716 41667
rect 23664 41624 23716 41633
rect 25872 41692 25924 41744
rect 26424 41556 26476 41608
rect 1676 41531 1728 41540
rect 1676 41497 1685 41531
rect 1685 41497 1719 41531
rect 1719 41497 1728 41531
rect 1676 41488 1728 41497
rect 10600 41420 10652 41472
rect 22376 41488 22428 41540
rect 32864 41760 32916 41812
rect 35532 41760 35584 41812
rect 36912 41760 36964 41812
rect 31668 41624 31720 41676
rect 34152 41624 34204 41676
rect 34520 41624 34572 41676
rect 34704 41624 34756 41676
rect 37832 41624 37884 41676
rect 29736 41556 29788 41608
rect 31208 41488 31260 41540
rect 31668 41531 31720 41540
rect 31668 41497 31677 41531
rect 31677 41497 31711 41531
rect 31711 41497 31720 41531
rect 31668 41488 31720 41497
rect 32956 41488 33008 41540
rect 24676 41420 24728 41472
rect 27252 41420 27304 41472
rect 34428 41488 34480 41540
rect 33324 41420 33376 41472
rect 34244 41420 34296 41472
rect 35808 41420 35860 41472
rect 36636 41488 36688 41540
rect 37004 41420 37056 41472
rect 39580 41488 39632 41540
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 27950 41318 28002 41370
rect 28014 41318 28066 41370
rect 28078 41318 28130 41370
rect 28142 41318 28194 41370
rect 28206 41318 28258 41370
rect 37950 41318 38002 41370
rect 38014 41318 38066 41370
rect 38078 41318 38130 41370
rect 38142 41318 38194 41370
rect 38206 41318 38258 41370
rect 47950 41318 48002 41370
rect 48014 41318 48066 41370
rect 48078 41318 48130 41370
rect 48142 41318 48194 41370
rect 48206 41318 48258 41370
rect 5816 41259 5868 41268
rect 5816 41225 5825 41259
rect 5825 41225 5859 41259
rect 5859 41225 5868 41259
rect 5816 41216 5868 41225
rect 9864 41259 9916 41268
rect 9864 41225 9873 41259
rect 9873 41225 9907 41259
rect 9907 41225 9916 41259
rect 9864 41216 9916 41225
rect 10784 41259 10836 41268
rect 10784 41225 10793 41259
rect 10793 41225 10827 41259
rect 10827 41225 10836 41259
rect 10784 41216 10836 41225
rect 22928 41216 22980 41268
rect 24860 41216 24912 41268
rect 1952 41148 2004 41200
rect 22468 41148 22520 41200
rect 25320 41148 25372 41200
rect 27804 41216 27856 41268
rect 30748 41148 30800 41200
rect 32864 41148 32916 41200
rect 34888 41216 34940 41268
rect 9772 41123 9824 41132
rect 9772 41089 9781 41123
rect 9781 41089 9815 41123
rect 9815 41089 9824 41123
rect 9772 41080 9824 41089
rect 10692 41123 10744 41132
rect 10692 41089 10701 41123
rect 10701 41089 10735 41123
rect 10735 41089 10744 41123
rect 10692 41080 10744 41089
rect 17684 41012 17736 41064
rect 21824 41012 21876 41064
rect 22376 41012 22428 41064
rect 27252 41123 27304 41132
rect 27252 41089 27261 41123
rect 27261 41089 27295 41123
rect 27295 41089 27304 41123
rect 27252 41080 27304 41089
rect 30840 41080 30892 41132
rect 24308 41012 24360 41064
rect 24584 41012 24636 41064
rect 25044 41055 25096 41064
rect 25044 41021 25053 41055
rect 25053 41021 25087 41055
rect 25087 41021 25096 41055
rect 25044 41012 25096 41021
rect 30012 41055 30064 41064
rect 30012 41021 30021 41055
rect 30021 41021 30055 41055
rect 30055 41021 30064 41055
rect 30012 41012 30064 41021
rect 32312 41012 32364 41064
rect 27252 40944 27304 40996
rect 31300 40944 31352 40996
rect 33048 40944 33100 40996
rect 33876 41012 33928 41064
rect 37004 41080 37056 41132
rect 37832 41080 37884 41132
rect 39580 41080 39632 41132
rect 38476 41055 38528 41064
rect 38476 41021 38485 41055
rect 38485 41021 38519 41055
rect 38519 41021 38528 41055
rect 38476 41012 38528 41021
rect 48504 41055 48556 41064
rect 48504 41021 48513 41055
rect 48513 41021 48547 41055
rect 48547 41021 48556 41055
rect 48504 41012 48556 41021
rect 48596 41012 48648 41064
rect 23388 40876 23440 40928
rect 26608 40876 26660 40928
rect 30380 40876 30432 40928
rect 32588 40876 32640 40928
rect 32956 40876 33008 40928
rect 34796 40876 34848 40928
rect 35716 40876 35768 40928
rect 39948 40919 40000 40928
rect 39948 40885 39957 40919
rect 39957 40885 39991 40919
rect 39991 40885 40000 40919
rect 39948 40876 40000 40885
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 32950 40774 33002 40826
rect 33014 40774 33066 40826
rect 33078 40774 33130 40826
rect 33142 40774 33194 40826
rect 33206 40774 33258 40826
rect 42950 40774 43002 40826
rect 43014 40774 43066 40826
rect 43078 40774 43130 40826
rect 43142 40774 43194 40826
rect 43206 40774 43258 40826
rect 22008 40672 22060 40724
rect 31024 40672 31076 40724
rect 20628 40604 20680 40656
rect 34428 40604 34480 40656
rect 25044 40536 25096 40588
rect 26608 40536 26660 40588
rect 27436 40536 27488 40588
rect 27712 40536 27764 40588
rect 28908 40536 28960 40588
rect 30012 40536 30064 40588
rect 32680 40579 32732 40588
rect 32680 40545 32689 40579
rect 32689 40545 32723 40579
rect 32723 40545 32732 40579
rect 32680 40536 32732 40545
rect 32772 40579 32824 40588
rect 32772 40545 32781 40579
rect 32781 40545 32815 40579
rect 32815 40545 32824 40579
rect 32772 40536 32824 40545
rect 33508 40536 33560 40588
rect 34152 40579 34204 40588
rect 34152 40545 34161 40579
rect 34161 40545 34195 40579
rect 34195 40545 34204 40579
rect 34152 40536 34204 40545
rect 38752 40536 38804 40588
rect 26976 40468 27028 40520
rect 27068 40511 27120 40520
rect 27068 40477 27077 40511
rect 27077 40477 27111 40511
rect 27111 40477 27120 40511
rect 27068 40468 27120 40477
rect 27528 40468 27580 40520
rect 29736 40511 29788 40520
rect 29736 40477 29745 40511
rect 29745 40477 29779 40511
rect 29779 40477 29788 40511
rect 29736 40468 29788 40477
rect 23480 40400 23532 40452
rect 28908 40400 28960 40452
rect 22192 40332 22244 40384
rect 26884 40332 26936 40384
rect 30472 40400 30524 40452
rect 31484 40332 31536 40384
rect 34152 40400 34204 40452
rect 37648 40400 37700 40452
rect 38844 40468 38896 40520
rect 39948 40536 40000 40588
rect 48412 40536 48464 40588
rect 48504 40511 48556 40520
rect 48504 40477 48513 40511
rect 48513 40477 48547 40511
rect 48547 40477 48556 40511
rect 48504 40468 48556 40477
rect 39212 40400 39264 40452
rect 33600 40375 33652 40384
rect 33600 40341 33609 40375
rect 33609 40341 33643 40375
rect 33643 40341 33652 40375
rect 33600 40332 33652 40341
rect 33692 40332 33744 40384
rect 37372 40332 37424 40384
rect 38384 40332 38436 40384
rect 38752 40375 38804 40384
rect 38752 40341 38761 40375
rect 38761 40341 38795 40375
rect 38795 40341 38804 40375
rect 38752 40332 38804 40341
rect 39120 40375 39172 40384
rect 39120 40341 39129 40375
rect 39129 40341 39163 40375
rect 39163 40341 39172 40375
rect 39120 40332 39172 40341
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 27950 40230 28002 40282
rect 28014 40230 28066 40282
rect 28078 40230 28130 40282
rect 28142 40230 28194 40282
rect 28206 40230 28258 40282
rect 37950 40230 38002 40282
rect 38014 40230 38066 40282
rect 38078 40230 38130 40282
rect 38142 40230 38194 40282
rect 38206 40230 38258 40282
rect 47950 40230 48002 40282
rect 48014 40230 48066 40282
rect 48078 40230 48130 40282
rect 48142 40230 48194 40282
rect 48206 40230 48258 40282
rect 25044 40128 25096 40180
rect 25320 40060 25372 40112
rect 30472 40128 30524 40180
rect 31300 40128 31352 40180
rect 35072 40128 35124 40180
rect 35900 40128 35952 40180
rect 36820 40128 36872 40180
rect 39488 40128 39540 40180
rect 42708 40128 42760 40180
rect 33876 40060 33928 40112
rect 38844 40103 38896 40112
rect 38844 40069 38853 40103
rect 38853 40069 38887 40103
rect 38887 40069 38896 40103
rect 38844 40060 38896 40069
rect 39580 40060 39632 40112
rect 41144 40103 41196 40112
rect 41144 40069 41153 40103
rect 41153 40069 41187 40103
rect 41187 40069 41196 40103
rect 41144 40060 41196 40069
rect 22652 39992 22704 40044
rect 34704 40035 34756 40044
rect 34704 40001 34713 40035
rect 34713 40001 34747 40035
rect 34747 40001 34756 40035
rect 34704 39992 34756 40001
rect 37832 39992 37884 40044
rect 38568 40035 38620 40044
rect 38568 40001 38577 40035
rect 38577 40001 38611 40035
rect 38611 40001 38620 40035
rect 38568 39992 38620 40001
rect 41236 40035 41288 40044
rect 41236 40001 41245 40035
rect 41245 40001 41279 40035
rect 41279 40001 41288 40035
rect 41236 39992 41288 40001
rect 23572 39924 23624 39976
rect 23664 39788 23716 39840
rect 27804 39788 27856 39840
rect 28448 39967 28500 39976
rect 28448 39933 28457 39967
rect 28457 39933 28491 39967
rect 28491 39933 28500 39967
rect 28448 39924 28500 39933
rect 32312 39967 32364 39976
rect 32312 39933 32321 39967
rect 32321 39933 32355 39967
rect 32355 39933 32364 39967
rect 32312 39924 32364 39933
rect 30380 39856 30432 39908
rect 33784 39924 33836 39976
rect 35624 39924 35676 39976
rect 40132 39924 40184 39976
rect 41788 39924 41840 39976
rect 48504 39967 48556 39976
rect 48504 39933 48513 39967
rect 48513 39933 48547 39967
rect 48547 39933 48556 39967
rect 48504 39924 48556 39933
rect 29736 39788 29788 39840
rect 29828 39788 29880 39840
rect 30104 39788 30156 39840
rect 34060 39788 34112 39840
rect 34336 39788 34388 39840
rect 41604 39856 41656 39908
rect 39948 39788 40000 39840
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 32950 39686 33002 39738
rect 33014 39686 33066 39738
rect 33078 39686 33130 39738
rect 33142 39686 33194 39738
rect 33206 39686 33258 39738
rect 42950 39686 43002 39738
rect 43014 39686 43066 39738
rect 43078 39686 43130 39738
rect 43142 39686 43194 39738
rect 43206 39686 43258 39738
rect 24400 39516 24452 39568
rect 22284 39448 22336 39500
rect 22468 39380 22520 39432
rect 28724 39584 28776 39636
rect 30840 39584 30892 39636
rect 31484 39516 31536 39568
rect 24584 39491 24636 39500
rect 24584 39457 24593 39491
rect 24593 39457 24627 39491
rect 24627 39457 24636 39491
rect 24584 39448 24636 39457
rect 24952 39448 25004 39500
rect 28356 39448 28408 39500
rect 32588 39448 32640 39500
rect 34060 39516 34112 39568
rect 35900 39516 35952 39568
rect 33508 39448 33560 39500
rect 38660 39584 38712 39636
rect 43812 39584 43864 39636
rect 43904 39584 43956 39636
rect 48320 39584 48372 39636
rect 38384 39516 38436 39568
rect 39948 39516 40000 39568
rect 37556 39448 37608 39500
rect 38292 39448 38344 39500
rect 38752 39448 38804 39500
rect 39304 39491 39356 39500
rect 39304 39457 39313 39491
rect 39313 39457 39347 39491
rect 39347 39457 39356 39491
rect 39304 39448 39356 39457
rect 42800 39448 42852 39500
rect 48780 39491 48832 39500
rect 48780 39457 48789 39491
rect 48789 39457 48823 39491
rect 48823 39457 48832 39491
rect 48780 39448 48832 39457
rect 28448 39380 28500 39432
rect 28816 39380 28868 39432
rect 34520 39380 34572 39432
rect 34704 39380 34756 39432
rect 40316 39380 40368 39432
rect 48504 39423 48556 39432
rect 48504 39389 48513 39423
rect 48513 39389 48547 39423
rect 48547 39389 48556 39423
rect 48504 39380 48556 39389
rect 1860 39244 1912 39296
rect 25136 39312 25188 39364
rect 25320 39312 25372 39364
rect 26148 39312 26200 39364
rect 23572 39244 23624 39296
rect 28632 39244 28684 39296
rect 29000 39312 29052 39364
rect 29460 39312 29512 39364
rect 30472 39355 30524 39364
rect 30472 39321 30481 39355
rect 30481 39321 30515 39355
rect 30515 39321 30524 39355
rect 30472 39312 30524 39321
rect 30564 39312 30616 39364
rect 31116 39244 31168 39296
rect 37004 39312 37056 39364
rect 39396 39312 39448 39364
rect 41236 39312 41288 39364
rect 43444 39312 43496 39364
rect 46388 39312 46440 39364
rect 34980 39244 35032 39296
rect 35256 39244 35308 39296
rect 37740 39287 37792 39296
rect 37740 39253 37749 39287
rect 37749 39253 37783 39287
rect 37783 39253 37792 39287
rect 37740 39244 37792 39253
rect 38844 39244 38896 39296
rect 39948 39244 40000 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 27950 39142 28002 39194
rect 28014 39142 28066 39194
rect 28078 39142 28130 39194
rect 28142 39142 28194 39194
rect 28206 39142 28258 39194
rect 37950 39142 38002 39194
rect 38014 39142 38066 39194
rect 38078 39142 38130 39194
rect 38142 39142 38194 39194
rect 38206 39142 38258 39194
rect 47950 39142 48002 39194
rect 48014 39142 48066 39194
rect 48078 39142 48130 39194
rect 48142 39142 48194 39194
rect 48206 39142 48258 39194
rect 940 38904 992 38956
rect 1860 38904 1912 38956
rect 23664 39040 23716 39092
rect 24492 39083 24544 39092
rect 24492 39049 24501 39083
rect 24501 39049 24535 39083
rect 24535 39049 24544 39083
rect 24492 39040 24544 39049
rect 25964 39040 26016 39092
rect 26240 39040 26292 39092
rect 27160 39040 27212 39092
rect 23388 38972 23440 39024
rect 24860 38947 24912 38956
rect 24860 38913 24869 38947
rect 24869 38913 24903 38947
rect 24903 38913 24912 38947
rect 24860 38904 24912 38913
rect 25136 38904 25188 38956
rect 26148 38904 26200 38956
rect 26240 38947 26292 38956
rect 26240 38913 26249 38947
rect 26249 38913 26283 38947
rect 26283 38913 26292 38947
rect 26240 38904 26292 38913
rect 28448 38972 28500 39024
rect 30104 39040 30156 39092
rect 30472 39040 30524 39092
rect 33508 39040 33560 39092
rect 33600 39040 33652 39092
rect 34428 39040 34480 39092
rect 35348 39040 35400 39092
rect 35624 39040 35676 39092
rect 35992 39083 36044 39092
rect 35992 39049 36001 39083
rect 36001 39049 36035 39083
rect 36035 39049 36044 39083
rect 35992 39040 36044 39049
rect 29920 38972 29972 39024
rect 34336 38972 34388 39024
rect 35440 38972 35492 39024
rect 24768 38836 24820 38888
rect 24952 38836 25004 38888
rect 25872 38836 25924 38888
rect 27896 38879 27948 38888
rect 27896 38845 27905 38879
rect 27905 38845 27939 38879
rect 27939 38845 27948 38879
rect 27896 38836 27948 38845
rect 25964 38768 26016 38820
rect 7380 38700 7432 38752
rect 27528 38700 27580 38752
rect 28356 38904 28408 38956
rect 28724 38836 28776 38888
rect 33324 38904 33376 38956
rect 36084 38972 36136 39024
rect 37280 39040 37332 39092
rect 38844 39040 38896 39092
rect 39120 39040 39172 39092
rect 40132 39040 40184 39092
rect 40408 39040 40460 39092
rect 36452 38972 36504 39024
rect 38292 38972 38344 39024
rect 38568 38972 38620 39024
rect 36176 38904 36228 38956
rect 37280 38904 37332 38956
rect 38844 38947 38896 38956
rect 38844 38913 38853 38947
rect 38853 38913 38887 38947
rect 38887 38913 38896 38947
rect 38844 38904 38896 38913
rect 39396 38904 39448 38956
rect 28080 38768 28132 38820
rect 28356 38768 28408 38820
rect 31944 38768 31996 38820
rect 34244 38879 34296 38888
rect 34244 38845 34253 38879
rect 34253 38845 34287 38879
rect 34287 38845 34296 38879
rect 34244 38836 34296 38845
rect 34888 38836 34940 38888
rect 33784 38768 33836 38820
rect 37188 38836 37240 38888
rect 37740 38836 37792 38888
rect 38936 38879 38988 38888
rect 38936 38845 38945 38879
rect 38945 38845 38979 38879
rect 38979 38845 38988 38879
rect 38936 38836 38988 38845
rect 39028 38879 39080 38888
rect 39028 38845 39037 38879
rect 39037 38845 39071 38879
rect 39071 38845 39080 38879
rect 39028 38836 39080 38845
rect 28540 38743 28592 38752
rect 28540 38709 28549 38743
rect 28549 38709 28583 38743
rect 28583 38709 28592 38743
rect 28540 38700 28592 38709
rect 32404 38743 32456 38752
rect 32404 38709 32413 38743
rect 32413 38709 32447 38743
rect 32447 38709 32456 38743
rect 32404 38700 32456 38709
rect 34980 38743 35032 38752
rect 34980 38709 34989 38743
rect 34989 38709 35023 38743
rect 35023 38709 35032 38743
rect 34980 38700 35032 38709
rect 37464 38743 37516 38752
rect 37464 38709 37473 38743
rect 37473 38709 37507 38743
rect 37507 38709 37516 38743
rect 37464 38700 37516 38709
rect 37832 38768 37884 38820
rect 38476 38768 38528 38820
rect 39948 38836 40000 38888
rect 43444 38972 43496 39024
rect 40316 38879 40368 38888
rect 40316 38845 40325 38879
rect 40325 38845 40359 38879
rect 40359 38845 40368 38879
rect 40316 38836 40368 38845
rect 41052 38836 41104 38888
rect 41236 38836 41288 38888
rect 43904 38836 43956 38888
rect 40960 38700 41012 38752
rect 41788 38700 41840 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 32950 38598 33002 38650
rect 33014 38598 33066 38650
rect 33078 38598 33130 38650
rect 33142 38598 33194 38650
rect 33206 38598 33258 38650
rect 42950 38598 43002 38650
rect 43014 38598 43066 38650
rect 43078 38598 43130 38650
rect 43142 38598 43194 38650
rect 43206 38598 43258 38650
rect 22100 38496 22152 38548
rect 26332 38496 26384 38548
rect 27252 38496 27304 38548
rect 31576 38496 31628 38548
rect 25044 38428 25096 38480
rect 26976 38428 27028 38480
rect 28632 38428 28684 38480
rect 20720 38360 20772 38412
rect 21088 38403 21140 38412
rect 21088 38369 21097 38403
rect 21097 38369 21131 38403
rect 21131 38369 21140 38403
rect 21088 38360 21140 38369
rect 22376 38360 22428 38412
rect 27528 38403 27580 38412
rect 27528 38369 27537 38403
rect 27537 38369 27571 38403
rect 27571 38369 27580 38403
rect 27528 38360 27580 38369
rect 24768 38292 24820 38344
rect 25044 38292 25096 38344
rect 26700 38292 26752 38344
rect 28540 38360 28592 38412
rect 31024 38428 31076 38480
rect 34428 38496 34480 38548
rect 36636 38539 36688 38548
rect 36636 38505 36645 38539
rect 36645 38505 36679 38539
rect 36679 38505 36688 38539
rect 36636 38496 36688 38505
rect 39212 38539 39264 38548
rect 39212 38505 39221 38539
rect 39221 38505 39255 38539
rect 39255 38505 39264 38539
rect 39212 38496 39264 38505
rect 41144 38496 41196 38548
rect 41236 38496 41288 38548
rect 34796 38428 34848 38480
rect 39488 38428 39540 38480
rect 27712 38292 27764 38344
rect 29736 38335 29788 38344
rect 29736 38301 29745 38335
rect 29745 38301 29779 38335
rect 29779 38301 29788 38335
rect 29736 38292 29788 38301
rect 31668 38292 31720 38344
rect 32588 38403 32640 38412
rect 32588 38369 32597 38403
rect 32597 38369 32631 38403
rect 32631 38369 32640 38403
rect 32588 38360 32640 38369
rect 32772 38360 32824 38412
rect 34152 38403 34204 38412
rect 34152 38369 34161 38403
rect 34161 38369 34195 38403
rect 34195 38369 34204 38403
rect 34152 38360 34204 38369
rect 21364 38267 21416 38276
rect 21364 38233 21373 38267
rect 21373 38233 21407 38267
rect 21407 38233 21416 38267
rect 21364 38224 21416 38233
rect 22100 38224 22152 38276
rect 25136 38224 25188 38276
rect 28540 38224 28592 38276
rect 29092 38224 29144 38276
rect 30012 38267 30064 38276
rect 30012 38233 30021 38267
rect 30021 38233 30055 38267
rect 30055 38233 30064 38267
rect 30012 38224 30064 38233
rect 30472 38224 30524 38276
rect 31576 38224 31628 38276
rect 31944 38224 31996 38276
rect 32036 38224 32088 38276
rect 34704 38360 34756 38412
rect 35808 38360 35860 38412
rect 35256 38224 35308 38276
rect 38292 38360 38344 38412
rect 41328 38428 41380 38480
rect 42800 38428 42852 38480
rect 43352 38428 43404 38480
rect 40500 38360 40552 38412
rect 41052 38360 41104 38412
rect 37004 38224 37056 38276
rect 37096 38267 37148 38276
rect 37096 38233 37105 38267
rect 37105 38233 37139 38267
rect 37139 38233 37148 38267
rect 37096 38224 37148 38233
rect 38476 38224 38528 38276
rect 25504 38156 25556 38208
rect 32220 38156 32272 38208
rect 33968 38156 34020 38208
rect 34060 38199 34112 38208
rect 34060 38165 34069 38199
rect 34069 38165 34103 38199
rect 34103 38165 34112 38199
rect 34060 38156 34112 38165
rect 35072 38156 35124 38208
rect 40132 38224 40184 38276
rect 39028 38156 39080 38208
rect 39856 38156 39908 38208
rect 48688 38360 48740 38412
rect 41512 38335 41564 38344
rect 41512 38301 41521 38335
rect 41521 38301 41555 38335
rect 41555 38301 41564 38335
rect 41512 38292 41564 38301
rect 49332 38335 49384 38344
rect 49332 38301 49341 38335
rect 49341 38301 49375 38335
rect 49375 38301 49384 38335
rect 49332 38292 49384 38301
rect 41788 38267 41840 38276
rect 41788 38233 41797 38267
rect 41797 38233 41831 38267
rect 41831 38233 41840 38267
rect 41788 38224 41840 38233
rect 43444 38224 43496 38276
rect 41328 38156 41380 38208
rect 48872 38156 48924 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 27950 38054 28002 38106
rect 28014 38054 28066 38106
rect 28078 38054 28130 38106
rect 28142 38054 28194 38106
rect 28206 38054 28258 38106
rect 37950 38054 38002 38106
rect 38014 38054 38066 38106
rect 38078 38054 38130 38106
rect 38142 38054 38194 38106
rect 38206 38054 38258 38106
rect 47950 38054 48002 38106
rect 48014 38054 48066 38106
rect 48078 38054 48130 38106
rect 48142 38054 48194 38106
rect 48206 38054 48258 38106
rect 22100 37884 22152 37936
rect 24124 37952 24176 38004
rect 25044 37952 25096 38004
rect 28172 37884 28224 37936
rect 29736 37952 29788 38004
rect 30656 37927 30708 37936
rect 30656 37893 30665 37927
rect 30665 37893 30699 37927
rect 30699 37893 30708 37927
rect 30656 37884 30708 37893
rect 31024 37816 31076 37868
rect 33508 37995 33560 38004
rect 33508 37961 33517 37995
rect 33517 37961 33551 37995
rect 33551 37961 33560 37995
rect 33508 37952 33560 37961
rect 33968 37995 34020 38004
rect 33968 37961 33977 37995
rect 33977 37961 34011 37995
rect 34011 37961 34020 37995
rect 33968 37952 34020 37961
rect 41236 37952 41288 38004
rect 31668 37884 31720 37936
rect 37096 37884 37148 37936
rect 39580 37884 39632 37936
rect 40132 37884 40184 37936
rect 43168 37952 43220 38004
rect 41972 37884 42024 37936
rect 32312 37816 32364 37868
rect 32680 37816 32732 37868
rect 33876 37859 33928 37868
rect 33876 37825 33885 37859
rect 33885 37825 33919 37859
rect 33919 37825 33928 37859
rect 33876 37816 33928 37825
rect 22468 37612 22520 37664
rect 26700 37748 26752 37800
rect 26792 37748 26844 37800
rect 27804 37748 27856 37800
rect 28908 37748 28960 37800
rect 30840 37748 30892 37800
rect 33416 37748 33468 37800
rect 28540 37680 28592 37732
rect 24676 37612 24728 37664
rect 24952 37612 25004 37664
rect 31300 37612 31352 37664
rect 31760 37680 31812 37732
rect 34704 37816 34756 37868
rect 38476 37748 38528 37800
rect 39212 37748 39264 37800
rect 37648 37612 37700 37664
rect 41328 37791 41380 37800
rect 41328 37757 41337 37791
rect 41337 37757 41371 37791
rect 41371 37757 41380 37791
rect 41328 37748 41380 37757
rect 49332 37859 49384 37868
rect 49332 37825 49341 37859
rect 49341 37825 49375 37859
rect 49375 37825 49384 37859
rect 49332 37816 49384 37825
rect 40132 37680 40184 37732
rect 43168 37791 43220 37800
rect 43168 37757 43177 37791
rect 43177 37757 43211 37791
rect 43211 37757 43220 37791
rect 43168 37748 43220 37757
rect 46940 37680 46992 37732
rect 39948 37612 40000 37664
rect 40316 37655 40368 37664
rect 40316 37621 40325 37655
rect 40325 37621 40359 37655
rect 40359 37621 40368 37655
rect 40316 37612 40368 37621
rect 42156 37612 42208 37664
rect 42248 37612 42300 37664
rect 44364 37612 44416 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 32950 37510 33002 37562
rect 33014 37510 33066 37562
rect 33078 37510 33130 37562
rect 33142 37510 33194 37562
rect 33206 37510 33258 37562
rect 42950 37510 43002 37562
rect 43014 37510 43066 37562
rect 43078 37510 43130 37562
rect 43142 37510 43194 37562
rect 43206 37510 43258 37562
rect 21548 37451 21600 37460
rect 21548 37417 21557 37451
rect 21557 37417 21591 37451
rect 21591 37417 21600 37451
rect 21548 37408 21600 37417
rect 22468 37247 22520 37256
rect 22468 37213 22477 37247
rect 22477 37213 22511 37247
rect 22511 37213 22520 37247
rect 22468 37204 22520 37213
rect 23572 37272 23624 37324
rect 27252 37408 27304 37460
rect 27804 37408 27856 37460
rect 30656 37408 30708 37460
rect 31668 37408 31720 37460
rect 33876 37408 33928 37460
rect 42248 37408 42300 37460
rect 43536 37408 43588 37460
rect 24676 37340 24728 37392
rect 24584 37272 24636 37324
rect 23296 37204 23348 37256
rect 14464 37136 14516 37188
rect 22192 37068 22244 37120
rect 23480 37068 23532 37120
rect 24400 37136 24452 37188
rect 29276 37340 29328 37392
rect 29828 37340 29880 37392
rect 27068 37315 27120 37324
rect 27068 37281 27077 37315
rect 27077 37281 27111 37315
rect 27111 37281 27120 37315
rect 27068 37272 27120 37281
rect 27620 37272 27672 37324
rect 28540 37272 28592 37324
rect 31208 37272 31260 37324
rect 31484 37315 31536 37324
rect 31484 37281 31493 37315
rect 31493 37281 31527 37315
rect 31527 37281 31536 37315
rect 31484 37272 31536 37281
rect 38108 37340 38160 37392
rect 38568 37383 38620 37392
rect 38568 37349 38577 37383
rect 38577 37349 38611 37383
rect 38611 37349 38620 37383
rect 38568 37340 38620 37349
rect 39764 37340 39816 37392
rect 39948 37340 40000 37392
rect 40040 37383 40092 37392
rect 40040 37349 40049 37383
rect 40049 37349 40083 37383
rect 40083 37349 40092 37383
rect 40040 37340 40092 37349
rect 37556 37315 37608 37324
rect 37556 37281 37565 37315
rect 37565 37281 37599 37315
rect 37599 37281 37608 37315
rect 37556 37272 37608 37281
rect 39212 37315 39264 37324
rect 39212 37281 39221 37315
rect 39221 37281 39255 37315
rect 39255 37281 39264 37315
rect 39212 37272 39264 37281
rect 26792 37247 26844 37256
rect 26792 37213 26801 37247
rect 26801 37213 26835 37247
rect 26835 37213 26844 37247
rect 26792 37204 26844 37213
rect 28172 37204 28224 37256
rect 28632 37204 28684 37256
rect 31300 37247 31352 37256
rect 31300 37213 31309 37247
rect 31309 37213 31343 37247
rect 31343 37213 31352 37247
rect 31300 37204 31352 37213
rect 32496 37204 32548 37256
rect 37096 37204 37148 37256
rect 39120 37204 39172 37256
rect 40684 37340 40736 37392
rect 40316 37272 40368 37324
rect 41512 37272 41564 37324
rect 42524 37272 42576 37324
rect 48504 37315 48556 37324
rect 48504 37281 48513 37315
rect 48513 37281 48547 37315
rect 48547 37281 48556 37315
rect 48504 37272 48556 37281
rect 40224 37204 40276 37256
rect 41420 37247 41472 37256
rect 41420 37213 41429 37247
rect 41429 37213 41463 37247
rect 41463 37213 41472 37247
rect 41420 37204 41472 37213
rect 48780 37247 48832 37256
rect 48780 37213 48789 37247
rect 48789 37213 48823 37247
rect 48823 37213 48832 37247
rect 48780 37204 48832 37213
rect 26976 37136 27028 37188
rect 25412 37068 25464 37120
rect 25504 37111 25556 37120
rect 25504 37077 25513 37111
rect 25513 37077 25547 37111
rect 25547 37077 25556 37111
rect 25504 37068 25556 37077
rect 33324 37136 33376 37188
rect 37556 37136 37608 37188
rect 38568 37136 38620 37188
rect 40684 37136 40736 37188
rect 29828 37068 29880 37120
rect 30748 37068 30800 37120
rect 31116 37068 31168 37120
rect 32128 37111 32180 37120
rect 32128 37077 32137 37111
rect 32137 37077 32171 37111
rect 32171 37077 32180 37111
rect 32128 37068 32180 37077
rect 32496 37111 32548 37120
rect 32496 37077 32505 37111
rect 32505 37077 32539 37111
rect 32539 37077 32548 37111
rect 32496 37068 32548 37077
rect 34244 37068 34296 37120
rect 34428 37068 34480 37120
rect 36912 37068 36964 37120
rect 37280 37068 37332 37120
rect 38108 37068 38160 37120
rect 41604 37068 41656 37120
rect 43444 37136 43496 37188
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 27950 36966 28002 37018
rect 28014 36966 28066 37018
rect 28078 36966 28130 37018
rect 28142 36966 28194 37018
rect 28206 36966 28258 37018
rect 37950 36966 38002 37018
rect 38014 36966 38066 37018
rect 38078 36966 38130 37018
rect 38142 36966 38194 37018
rect 38206 36966 38258 37018
rect 47950 36966 48002 37018
rect 48014 36966 48066 37018
rect 48078 36966 48130 37018
rect 48142 36966 48194 37018
rect 48206 36966 48258 37018
rect 19432 36907 19484 36916
rect 19432 36873 19441 36907
rect 19441 36873 19475 36907
rect 19475 36873 19484 36907
rect 19432 36864 19484 36873
rect 32036 36864 32088 36916
rect 21824 36796 21876 36848
rect 22100 36796 22152 36848
rect 24124 36796 24176 36848
rect 940 36728 992 36780
rect 17224 36728 17276 36780
rect 22008 36728 22060 36780
rect 22652 36728 22704 36780
rect 25504 36728 25556 36780
rect 21364 36660 21416 36712
rect 24952 36660 25004 36712
rect 25596 36660 25648 36712
rect 26424 36703 26476 36712
rect 26424 36669 26433 36703
rect 26433 36669 26467 36703
rect 26467 36669 26476 36703
rect 26424 36660 26476 36669
rect 27528 36771 27580 36780
rect 27528 36737 27537 36771
rect 27537 36737 27571 36771
rect 27571 36737 27580 36771
rect 27528 36728 27580 36737
rect 28724 36728 28776 36780
rect 30472 36796 30524 36848
rect 32404 36864 32456 36916
rect 34888 36864 34940 36916
rect 37372 36864 37424 36916
rect 39120 36796 39172 36848
rect 39672 36796 39724 36848
rect 32220 36728 32272 36780
rect 35808 36728 35860 36780
rect 38844 36728 38896 36780
rect 29368 36660 29420 36712
rect 29184 36592 29236 36644
rect 7564 36524 7616 36576
rect 23664 36524 23716 36576
rect 25872 36567 25924 36576
rect 25872 36533 25881 36567
rect 25881 36533 25915 36567
rect 25915 36533 25924 36567
rect 25872 36524 25924 36533
rect 29460 36524 29512 36576
rect 31668 36660 31720 36712
rect 32312 36660 32364 36712
rect 33968 36660 34020 36712
rect 35072 36660 35124 36712
rect 37372 36660 37424 36712
rect 33876 36592 33928 36644
rect 35072 36524 35124 36576
rect 35164 36524 35216 36576
rect 38476 36660 38528 36712
rect 41512 36864 41564 36916
rect 41604 36864 41656 36916
rect 48964 36864 49016 36916
rect 39948 36796 40000 36848
rect 42708 36796 42760 36848
rect 41328 36728 41380 36780
rect 49332 36771 49384 36780
rect 49332 36737 49341 36771
rect 49341 36737 49375 36771
rect 49375 36737 49384 36771
rect 49332 36728 49384 36737
rect 38568 36592 38620 36644
rect 39672 36592 39724 36644
rect 43352 36660 43404 36712
rect 43444 36592 43496 36644
rect 36728 36524 36780 36576
rect 36912 36524 36964 36576
rect 38016 36524 38068 36576
rect 41052 36524 41104 36576
rect 42524 36524 42576 36576
rect 46940 36524 46992 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 32950 36422 33002 36474
rect 33014 36422 33066 36474
rect 33078 36422 33130 36474
rect 33142 36422 33194 36474
rect 33206 36422 33258 36474
rect 42950 36422 43002 36474
rect 43014 36422 43066 36474
rect 43078 36422 43130 36474
rect 43142 36422 43194 36474
rect 43206 36422 43258 36474
rect 22376 36320 22428 36372
rect 26240 36320 26292 36372
rect 27528 36320 27580 36372
rect 29460 36320 29512 36372
rect 21916 36252 21968 36304
rect 23572 36252 23624 36304
rect 20536 36227 20588 36236
rect 20536 36193 20545 36227
rect 20545 36193 20579 36227
rect 20579 36193 20588 36227
rect 20536 36184 20588 36193
rect 23388 36184 23440 36236
rect 23664 36159 23716 36168
rect 23664 36125 23673 36159
rect 23673 36125 23707 36159
rect 23707 36125 23716 36159
rect 23664 36116 23716 36125
rect 24308 36184 24360 36236
rect 26608 36116 26660 36168
rect 31852 36252 31904 36304
rect 32036 36363 32088 36372
rect 32036 36329 32045 36363
rect 32045 36329 32079 36363
rect 32079 36329 32088 36363
rect 32036 36320 32088 36329
rect 33508 36320 33560 36372
rect 34152 36320 34204 36372
rect 37372 36320 37424 36372
rect 37648 36320 37700 36372
rect 41328 36320 41380 36372
rect 34060 36252 34112 36304
rect 36544 36252 36596 36304
rect 28356 36227 28408 36236
rect 28356 36193 28365 36227
rect 28365 36193 28399 36227
rect 28399 36193 28408 36227
rect 28356 36184 28408 36193
rect 28816 36184 28868 36236
rect 30472 36184 30524 36236
rect 31760 36184 31812 36236
rect 28264 36159 28316 36168
rect 28264 36125 28273 36159
rect 28273 36125 28307 36159
rect 28307 36125 28316 36159
rect 28264 36116 28316 36125
rect 32772 36184 32824 36236
rect 35532 36227 35584 36236
rect 35532 36193 35541 36227
rect 35541 36193 35575 36227
rect 35575 36193 35584 36227
rect 35532 36184 35584 36193
rect 35716 36227 35768 36236
rect 35716 36193 35725 36227
rect 35725 36193 35759 36227
rect 35759 36193 35768 36227
rect 35716 36184 35768 36193
rect 36452 36184 36504 36236
rect 36820 36227 36872 36236
rect 36820 36193 36829 36227
rect 36829 36193 36863 36227
rect 36863 36193 36872 36227
rect 36820 36184 36872 36193
rect 40592 36252 40644 36304
rect 48780 36320 48832 36372
rect 38016 36227 38068 36236
rect 38016 36193 38025 36227
rect 38025 36193 38059 36227
rect 38059 36193 38068 36227
rect 38016 36184 38068 36193
rect 42800 36252 42852 36304
rect 32680 36116 32732 36168
rect 34612 36116 34664 36168
rect 37740 36116 37792 36168
rect 41788 36184 41840 36236
rect 42340 36227 42392 36236
rect 42340 36193 42349 36227
rect 42349 36193 42383 36227
rect 42383 36193 42392 36227
rect 42340 36184 42392 36193
rect 42708 36184 42760 36236
rect 41420 36116 41472 36168
rect 21824 36048 21876 36100
rect 24584 36048 24636 36100
rect 26976 36048 27028 36100
rect 33048 36048 33100 36100
rect 33140 36048 33192 36100
rect 23572 35980 23624 36032
rect 26240 35980 26292 36032
rect 34060 35980 34112 36032
rect 37096 36048 37148 36100
rect 37556 36048 37608 36100
rect 40132 36048 40184 36100
rect 36452 35980 36504 36032
rect 40592 36023 40644 36032
rect 40592 35989 40601 36023
rect 40601 35989 40635 36023
rect 40635 35989 40644 36023
rect 40592 35980 40644 35989
rect 42248 36023 42300 36032
rect 42248 35989 42257 36023
rect 42257 35989 42291 36023
rect 42291 35989 42300 36023
rect 42248 35980 42300 35989
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 27950 35878 28002 35930
rect 28014 35878 28066 35930
rect 28078 35878 28130 35930
rect 28142 35878 28194 35930
rect 28206 35878 28258 35930
rect 37950 35878 38002 35930
rect 38014 35878 38066 35930
rect 38078 35878 38130 35930
rect 38142 35878 38194 35930
rect 38206 35878 38258 35930
rect 47950 35878 48002 35930
rect 48014 35878 48066 35930
rect 48078 35878 48130 35930
rect 48142 35878 48194 35930
rect 48206 35878 48258 35930
rect 16120 35776 16172 35828
rect 21180 35776 21232 35828
rect 21364 35776 21416 35828
rect 24768 35776 24820 35828
rect 21916 35708 21968 35760
rect 26424 35819 26476 35828
rect 26424 35785 26433 35819
rect 26433 35785 26467 35819
rect 26467 35785 26476 35819
rect 26424 35776 26476 35785
rect 26700 35776 26752 35828
rect 28632 35708 28684 35760
rect 24676 35683 24728 35692
rect 24676 35649 24685 35683
rect 24685 35649 24719 35683
rect 24719 35649 24728 35683
rect 24676 35640 24728 35649
rect 26792 35640 26844 35692
rect 32220 35776 32272 35828
rect 32588 35776 32640 35828
rect 33048 35776 33100 35828
rect 38752 35776 38804 35828
rect 39396 35776 39448 35828
rect 30380 35708 30432 35760
rect 30748 35708 30800 35760
rect 23296 35572 23348 35624
rect 25044 35572 25096 35624
rect 20536 35436 20588 35488
rect 21180 35436 21232 35488
rect 27712 35572 27764 35624
rect 29368 35615 29420 35624
rect 29368 35581 29377 35615
rect 29377 35581 29411 35615
rect 29411 35581 29420 35615
rect 31576 35640 31628 35692
rect 29368 35572 29420 35581
rect 27068 35504 27120 35556
rect 26884 35436 26936 35488
rect 32312 35572 32364 35624
rect 32772 35751 32824 35760
rect 32772 35717 32781 35751
rect 32781 35717 32815 35751
rect 32815 35717 32824 35751
rect 32772 35708 32824 35717
rect 35256 35640 35308 35692
rect 32864 35615 32916 35624
rect 32864 35581 32873 35615
rect 32873 35581 32907 35615
rect 32907 35581 32916 35615
rect 32864 35572 32916 35581
rect 34704 35572 34756 35624
rect 36820 35640 36872 35692
rect 37648 35640 37700 35692
rect 38476 35708 38528 35760
rect 39672 35708 39724 35760
rect 39948 35776 40000 35828
rect 40132 35776 40184 35828
rect 40776 35776 40828 35828
rect 49056 35776 49108 35828
rect 40224 35708 40276 35760
rect 41880 35708 41932 35760
rect 43168 35708 43220 35760
rect 43444 35708 43496 35760
rect 37832 35572 37884 35624
rect 38384 35615 38436 35624
rect 38384 35581 38393 35615
rect 38393 35581 38427 35615
rect 38427 35581 38436 35615
rect 38384 35572 38436 35581
rect 39764 35572 39816 35624
rect 40408 35572 40460 35624
rect 42616 35683 42668 35692
rect 42616 35649 42625 35683
rect 42625 35649 42659 35683
rect 42659 35649 42668 35683
rect 42616 35640 42668 35649
rect 49332 35683 49384 35692
rect 49332 35649 49341 35683
rect 49341 35649 49375 35683
rect 49375 35649 49384 35683
rect 49332 35640 49384 35649
rect 42340 35572 42392 35624
rect 42248 35504 42300 35556
rect 31760 35479 31812 35488
rect 31760 35445 31769 35479
rect 31769 35445 31803 35479
rect 31803 35445 31812 35479
rect 31760 35436 31812 35445
rect 33140 35436 33192 35488
rect 38936 35436 38988 35488
rect 42708 35436 42760 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 32950 35334 33002 35386
rect 33014 35334 33066 35386
rect 33078 35334 33130 35386
rect 33142 35334 33194 35386
rect 33206 35334 33258 35386
rect 42950 35334 43002 35386
rect 43014 35334 43066 35386
rect 43078 35334 43130 35386
rect 43142 35334 43194 35386
rect 43206 35334 43258 35386
rect 22008 35232 22060 35284
rect 25964 35232 26016 35284
rect 26884 35232 26936 35284
rect 27528 35232 27580 35284
rect 29184 35232 29236 35284
rect 30748 35232 30800 35284
rect 33876 35232 33928 35284
rect 35072 35232 35124 35284
rect 38752 35232 38804 35284
rect 49148 35232 49200 35284
rect 22100 35096 22152 35148
rect 20536 35028 20588 35080
rect 21732 35071 21784 35080
rect 21732 35037 21741 35071
rect 21741 35037 21775 35071
rect 21775 35037 21784 35071
rect 21732 35028 21784 35037
rect 23296 35096 23348 35148
rect 21916 34892 21968 34944
rect 24768 34960 24820 35012
rect 26240 35028 26292 35080
rect 27068 35164 27120 35216
rect 28908 35164 28960 35216
rect 26792 35096 26844 35148
rect 30012 35096 30064 35148
rect 30288 35139 30340 35148
rect 30288 35105 30297 35139
rect 30297 35105 30331 35139
rect 30331 35105 30340 35139
rect 30288 35096 30340 35105
rect 31208 35096 31260 35148
rect 31668 35139 31720 35148
rect 31668 35105 31677 35139
rect 31677 35105 31711 35139
rect 31711 35105 31720 35139
rect 31668 35096 31720 35105
rect 28632 35028 28684 35080
rect 28816 35028 28868 35080
rect 30104 35071 30156 35080
rect 30104 35037 30113 35071
rect 30113 35037 30147 35071
rect 30147 35037 30156 35071
rect 30104 35028 30156 35037
rect 31392 35071 31444 35080
rect 31392 35037 31401 35071
rect 31401 35037 31435 35071
rect 31435 35037 31444 35071
rect 31392 35028 31444 35037
rect 25596 34960 25648 35012
rect 26332 34960 26384 35012
rect 26608 34960 26660 35012
rect 24584 34892 24636 34944
rect 27804 34892 27856 34944
rect 30564 34960 30616 35012
rect 32220 35139 32272 35148
rect 32220 35105 32229 35139
rect 32229 35105 32263 35139
rect 32263 35105 32272 35139
rect 32220 35096 32272 35105
rect 36820 35164 36872 35216
rect 39028 35164 39080 35216
rect 36636 35139 36688 35148
rect 36636 35105 36645 35139
rect 36645 35105 36679 35139
rect 36679 35105 36688 35139
rect 36636 35096 36688 35105
rect 36728 35096 36780 35148
rect 38660 35096 38712 35148
rect 42616 35096 42668 35148
rect 43536 35096 43588 35148
rect 31024 34935 31076 34944
rect 31024 34901 31033 34935
rect 31033 34901 31067 34935
rect 31067 34901 31076 34935
rect 31024 34892 31076 34901
rect 31208 34892 31260 34944
rect 32772 34892 32824 34944
rect 33416 34892 33468 34944
rect 34980 35028 35032 35080
rect 35808 35028 35860 35080
rect 37464 35028 37516 35080
rect 39856 35028 39908 35080
rect 41696 35028 41748 35080
rect 34520 34960 34572 35012
rect 36176 34892 36228 34944
rect 36360 34935 36412 34944
rect 36360 34901 36369 34935
rect 36369 34901 36403 34935
rect 36403 34901 36412 34935
rect 36360 34892 36412 34901
rect 42432 34960 42484 35012
rect 42708 34960 42760 35012
rect 43444 34960 43496 35012
rect 38936 34935 38988 34944
rect 38936 34901 38945 34935
rect 38945 34901 38979 34935
rect 38979 34901 38988 34935
rect 38936 34892 38988 34901
rect 40500 34892 40552 34944
rect 40868 34892 40920 34944
rect 48412 35028 48464 35080
rect 49332 35071 49384 35080
rect 49332 35037 49341 35071
rect 49341 35037 49375 35071
rect 49375 35037 49384 35071
rect 49332 35028 49384 35037
rect 44548 34892 44600 34944
rect 46940 34892 46992 34944
rect 49056 34892 49108 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 27950 34790 28002 34842
rect 28014 34790 28066 34842
rect 28078 34790 28130 34842
rect 28142 34790 28194 34842
rect 28206 34790 28258 34842
rect 37950 34790 38002 34842
rect 38014 34790 38066 34842
rect 38078 34790 38130 34842
rect 38142 34790 38194 34842
rect 38206 34790 38258 34842
rect 47950 34790 48002 34842
rect 48014 34790 48066 34842
rect 48078 34790 48130 34842
rect 48142 34790 48194 34842
rect 48206 34790 48258 34842
rect 7840 34688 7892 34740
rect 24860 34688 24912 34740
rect 25596 34688 25648 34740
rect 28264 34688 28316 34740
rect 29184 34688 29236 34740
rect 24768 34620 24820 34672
rect 28632 34620 28684 34672
rect 30380 34620 30432 34672
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 22652 34552 22704 34604
rect 25688 34595 25740 34604
rect 25688 34561 25697 34595
rect 25697 34561 25731 34595
rect 25731 34561 25740 34595
rect 25688 34552 25740 34561
rect 26792 34552 26844 34604
rect 29920 34552 29972 34604
rect 31300 34688 31352 34740
rect 31760 34688 31812 34740
rect 32772 34731 32824 34740
rect 32772 34697 32781 34731
rect 32781 34697 32815 34731
rect 32815 34697 32824 34731
rect 32772 34688 32824 34697
rect 32588 34552 32640 34604
rect 32680 34552 32732 34604
rect 34612 34620 34664 34672
rect 34980 34620 35032 34672
rect 24860 34484 24912 34536
rect 26424 34484 26476 34536
rect 24308 34416 24360 34468
rect 30932 34416 30984 34468
rect 33968 34484 34020 34536
rect 37648 34620 37700 34672
rect 40040 34688 40092 34740
rect 40500 34731 40552 34740
rect 40500 34697 40509 34731
rect 40509 34697 40543 34731
rect 40543 34697 40552 34731
rect 40500 34688 40552 34697
rect 40960 34688 41012 34740
rect 41236 34620 41288 34672
rect 41696 34731 41748 34740
rect 41696 34697 41705 34731
rect 41705 34697 41739 34731
rect 41739 34697 41748 34731
rect 41696 34688 41748 34697
rect 42800 34688 42852 34740
rect 49148 34731 49200 34740
rect 49148 34697 49157 34731
rect 49157 34697 49191 34731
rect 49191 34697 49200 34731
rect 49148 34688 49200 34697
rect 37280 34552 37332 34604
rect 37096 34484 37148 34536
rect 39948 34484 40000 34536
rect 33784 34416 33836 34468
rect 37740 34416 37792 34468
rect 38568 34416 38620 34468
rect 40500 34552 40552 34604
rect 44548 34552 44600 34604
rect 49332 34595 49384 34604
rect 49332 34561 49341 34595
rect 49341 34561 49375 34595
rect 49375 34561 49384 34595
rect 49332 34552 49384 34561
rect 40868 34484 40920 34536
rect 42708 34484 42760 34536
rect 43536 34527 43588 34536
rect 43536 34493 43545 34527
rect 43545 34493 43579 34527
rect 43579 34493 43588 34527
rect 43536 34484 43588 34493
rect 41604 34416 41656 34468
rect 44272 34484 44324 34536
rect 22376 34348 22428 34400
rect 27712 34348 27764 34400
rect 29276 34348 29328 34400
rect 30012 34391 30064 34400
rect 30012 34357 30021 34391
rect 30021 34357 30055 34391
rect 30055 34357 30064 34391
rect 30012 34348 30064 34357
rect 31484 34348 31536 34400
rect 39764 34348 39816 34400
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 32950 34246 33002 34298
rect 33014 34246 33066 34298
rect 33078 34246 33130 34298
rect 33142 34246 33194 34298
rect 33206 34246 33258 34298
rect 42950 34246 43002 34298
rect 43014 34246 43066 34298
rect 43078 34246 43130 34298
rect 43142 34246 43194 34298
rect 43206 34246 43258 34298
rect 20996 34144 21048 34196
rect 27528 34144 27580 34196
rect 29092 34144 29144 34196
rect 35992 34144 36044 34196
rect 40592 34144 40644 34196
rect 22560 34076 22612 34128
rect 36360 34076 36412 34128
rect 24032 34008 24084 34060
rect 25596 34008 25648 34060
rect 27528 34008 27580 34060
rect 30380 34008 30432 34060
rect 35348 34008 35400 34060
rect 37372 34076 37424 34128
rect 48964 34144 49016 34196
rect 42064 34076 42116 34128
rect 26056 33872 26108 33924
rect 29092 33940 29144 33992
rect 26792 33872 26844 33924
rect 28816 33872 28868 33924
rect 32588 33872 32640 33924
rect 38476 34008 38528 34060
rect 42156 34051 42208 34060
rect 42156 34017 42165 34051
rect 42165 34017 42199 34051
rect 42199 34017 42208 34051
rect 42156 34008 42208 34017
rect 37464 33940 37516 33992
rect 38568 33983 38620 33992
rect 38568 33949 38577 33983
rect 38577 33949 38611 33983
rect 38611 33949 38620 33983
rect 38568 33940 38620 33949
rect 38660 33983 38712 33992
rect 38660 33949 38669 33983
rect 38669 33949 38703 33983
rect 38703 33949 38712 33983
rect 38660 33940 38712 33949
rect 41052 33940 41104 33992
rect 41972 33940 42024 33992
rect 49332 33983 49384 33992
rect 49332 33949 49341 33983
rect 49341 33949 49375 33983
rect 49375 33949 49384 33983
rect 49332 33940 49384 33949
rect 22744 33804 22796 33856
rect 24676 33804 24728 33856
rect 27528 33804 27580 33856
rect 31208 33847 31260 33856
rect 31208 33813 31217 33847
rect 31217 33813 31251 33847
rect 31251 33813 31260 33847
rect 31208 33804 31260 33813
rect 33692 33804 33744 33856
rect 37464 33804 37516 33856
rect 37740 33804 37792 33856
rect 38844 33804 38896 33856
rect 49240 33872 49292 33924
rect 41420 33804 41472 33856
rect 41880 33804 41932 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 27950 33702 28002 33754
rect 28014 33702 28066 33754
rect 28078 33702 28130 33754
rect 28142 33702 28194 33754
rect 28206 33702 28258 33754
rect 37950 33702 38002 33754
rect 38014 33702 38066 33754
rect 38078 33702 38130 33754
rect 38142 33702 38194 33754
rect 38206 33702 38258 33754
rect 47950 33702 48002 33754
rect 48014 33702 48066 33754
rect 48078 33702 48130 33754
rect 48142 33702 48194 33754
rect 48206 33702 48258 33754
rect 24032 33600 24084 33652
rect 25136 33600 25188 33652
rect 28724 33643 28776 33652
rect 28724 33609 28733 33643
rect 28733 33609 28767 33643
rect 28767 33609 28776 33643
rect 28724 33600 28776 33609
rect 29092 33643 29144 33652
rect 29092 33609 29101 33643
rect 29101 33609 29135 33643
rect 29135 33609 29144 33643
rect 29092 33600 29144 33609
rect 24768 33532 24820 33584
rect 25136 33464 25188 33516
rect 27436 33464 27488 33516
rect 21088 33396 21140 33448
rect 21732 33396 21784 33448
rect 24584 33396 24636 33448
rect 27068 33396 27120 33448
rect 29184 33439 29236 33448
rect 29184 33405 29193 33439
rect 29193 33405 29227 33439
rect 29227 33405 29236 33439
rect 29184 33396 29236 33405
rect 29644 33464 29696 33516
rect 34060 33600 34112 33652
rect 34888 33600 34940 33652
rect 42340 33600 42392 33652
rect 30380 33532 30432 33584
rect 33876 33532 33928 33584
rect 34980 33532 35032 33584
rect 37464 33532 37516 33584
rect 40868 33532 40920 33584
rect 42616 33532 42668 33584
rect 43444 33532 43496 33584
rect 33968 33507 34020 33516
rect 33968 33473 33977 33507
rect 33977 33473 34011 33507
rect 34011 33473 34020 33507
rect 33968 33464 34020 33473
rect 34244 33396 34296 33448
rect 34704 33396 34756 33448
rect 36912 33396 36964 33448
rect 37832 33507 37884 33516
rect 37832 33473 37841 33507
rect 37841 33473 37875 33507
rect 37875 33473 37884 33507
rect 37832 33464 37884 33473
rect 39212 33507 39264 33516
rect 39212 33473 39221 33507
rect 39221 33473 39255 33507
rect 39255 33473 39264 33507
rect 39212 33464 39264 33473
rect 40224 33464 40276 33516
rect 30564 33328 30616 33380
rect 22376 33260 22428 33312
rect 28356 33260 28408 33312
rect 29920 33303 29972 33312
rect 29920 33269 29929 33303
rect 29929 33269 29963 33303
rect 29963 33269 29972 33303
rect 29920 33260 29972 33269
rect 31576 33260 31628 33312
rect 37004 33328 37056 33380
rect 37464 33371 37516 33380
rect 37464 33337 37473 33371
rect 37473 33337 37507 33371
rect 37507 33337 37516 33371
rect 37464 33328 37516 33337
rect 35900 33260 35952 33312
rect 38200 33328 38252 33380
rect 40316 33439 40368 33448
rect 40316 33405 40325 33439
rect 40325 33405 40359 33439
rect 40359 33405 40368 33439
rect 40316 33396 40368 33405
rect 40592 33439 40644 33448
rect 40592 33405 40601 33439
rect 40601 33405 40635 33439
rect 40635 33405 40644 33439
rect 40592 33396 40644 33405
rect 41144 33396 41196 33448
rect 38844 33260 38896 33312
rect 42064 33303 42116 33312
rect 42064 33269 42073 33303
rect 42073 33269 42107 33303
rect 42107 33269 42116 33303
rect 42064 33260 42116 33269
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 32950 33158 33002 33210
rect 33014 33158 33066 33210
rect 33078 33158 33130 33210
rect 33142 33158 33194 33210
rect 33206 33158 33258 33210
rect 42950 33158 43002 33210
rect 43014 33158 43066 33210
rect 43078 33158 43130 33210
rect 43142 33158 43194 33210
rect 43206 33158 43258 33210
rect 22836 33099 22888 33108
rect 22836 33065 22845 33099
rect 22845 33065 22879 33099
rect 22879 33065 22888 33099
rect 22836 33056 22888 33065
rect 23296 33056 23348 33108
rect 27528 33056 27580 33108
rect 28908 33056 28960 33108
rect 26056 32988 26108 33040
rect 22376 32920 22428 32972
rect 21088 32895 21140 32904
rect 21088 32861 21097 32895
rect 21097 32861 21131 32895
rect 21131 32861 21140 32895
rect 21088 32852 21140 32861
rect 23664 32920 23716 32972
rect 26792 32920 26844 32972
rect 12072 32716 12124 32768
rect 26884 32852 26936 32904
rect 23664 32716 23716 32768
rect 24768 32716 24820 32768
rect 26608 32759 26660 32768
rect 26608 32725 26617 32759
rect 26617 32725 26651 32759
rect 26651 32725 26660 32759
rect 26608 32716 26660 32725
rect 28356 32920 28408 32972
rect 28724 32920 28776 32972
rect 31852 33056 31904 33108
rect 32588 33056 32640 33108
rect 36912 33056 36964 33108
rect 29276 32920 29328 32972
rect 30380 32963 30432 32972
rect 30380 32929 30389 32963
rect 30389 32929 30423 32963
rect 30423 32929 30432 32963
rect 30380 32920 30432 32929
rect 31484 32963 31536 32972
rect 31484 32929 31493 32963
rect 31493 32929 31527 32963
rect 31527 32929 31536 32963
rect 31484 32920 31536 32929
rect 40592 32988 40644 33040
rect 31024 32852 31076 32904
rect 32128 32852 32180 32904
rect 29000 32716 29052 32768
rect 34612 32784 34664 32836
rect 37280 32920 37332 32972
rect 37556 32920 37608 32972
rect 40684 32920 40736 32972
rect 41236 32920 41288 32972
rect 36268 32895 36320 32904
rect 36268 32861 36277 32895
rect 36277 32861 36311 32895
rect 36311 32861 36320 32895
rect 36268 32852 36320 32861
rect 38752 32895 38804 32904
rect 38752 32861 38761 32895
rect 38761 32861 38795 32895
rect 38795 32861 38804 32895
rect 38752 32852 38804 32861
rect 39028 32852 39080 32904
rect 40776 32895 40828 32904
rect 40776 32861 40785 32895
rect 40785 32861 40819 32895
rect 40819 32861 40828 32895
rect 40776 32852 40828 32861
rect 30932 32716 30984 32768
rect 31300 32759 31352 32768
rect 31300 32725 31309 32759
rect 31309 32725 31343 32759
rect 31343 32725 31352 32759
rect 31300 32716 31352 32725
rect 34060 32716 34112 32768
rect 34980 32716 35032 32768
rect 35900 32716 35952 32768
rect 37280 32784 37332 32836
rect 37832 32784 37884 32836
rect 48780 32988 48832 33040
rect 41788 32920 41840 32972
rect 42248 32963 42300 32972
rect 42248 32929 42257 32963
rect 42257 32929 42291 32963
rect 42291 32929 42300 32963
rect 42248 32920 42300 32929
rect 42340 32852 42392 32904
rect 43812 32895 43864 32904
rect 43812 32861 43821 32895
rect 43821 32861 43855 32895
rect 43855 32861 43864 32895
rect 43812 32852 43864 32861
rect 49332 32895 49384 32904
rect 49332 32861 49341 32895
rect 49341 32861 49375 32895
rect 49375 32861 49384 32895
rect 49332 32852 49384 32861
rect 38292 32716 38344 32768
rect 38752 32716 38804 32768
rect 39304 32716 39356 32768
rect 40224 32716 40276 32768
rect 41052 32716 41104 32768
rect 47216 32716 47268 32768
rect 49148 32759 49200 32768
rect 49148 32725 49157 32759
rect 49157 32725 49191 32759
rect 49191 32725 49200 32759
rect 49148 32716 49200 32725
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 27950 32614 28002 32666
rect 28014 32614 28066 32666
rect 28078 32614 28130 32666
rect 28142 32614 28194 32666
rect 28206 32614 28258 32666
rect 37950 32614 38002 32666
rect 38014 32614 38066 32666
rect 38078 32614 38130 32666
rect 38142 32614 38194 32666
rect 38206 32614 38258 32666
rect 47950 32614 48002 32666
rect 48014 32614 48066 32666
rect 48078 32614 48130 32666
rect 48142 32614 48194 32666
rect 48206 32614 48258 32666
rect 17224 32555 17276 32564
rect 17224 32521 17233 32555
rect 17233 32521 17267 32555
rect 17267 32521 17276 32555
rect 17224 32512 17276 32521
rect 17684 32555 17736 32564
rect 17684 32521 17693 32555
rect 17693 32521 17727 32555
rect 17727 32521 17736 32555
rect 17684 32512 17736 32521
rect 13452 32444 13504 32496
rect 23756 32444 23808 32496
rect 24768 32444 24820 32496
rect 940 32376 992 32428
rect 22652 32376 22704 32428
rect 23480 32376 23532 32428
rect 22836 32308 22888 32360
rect 24124 32351 24176 32360
rect 24124 32317 24133 32351
rect 24133 32317 24167 32351
rect 24167 32317 24176 32351
rect 24124 32308 24176 32317
rect 24768 32308 24820 32360
rect 25596 32555 25648 32564
rect 25596 32521 25605 32555
rect 25605 32521 25639 32555
rect 25639 32521 25648 32555
rect 25596 32512 25648 32521
rect 26056 32512 26108 32564
rect 31300 32512 31352 32564
rect 31576 32512 31628 32564
rect 26608 32444 26660 32496
rect 31116 32444 31168 32496
rect 34060 32444 34112 32496
rect 37740 32512 37792 32564
rect 29092 32376 29144 32428
rect 30380 32376 30432 32428
rect 26424 32240 26476 32292
rect 7472 32172 7524 32224
rect 20260 32172 20312 32224
rect 25964 32172 26016 32224
rect 27160 32172 27212 32224
rect 27896 32351 27948 32360
rect 27896 32317 27905 32351
rect 27905 32317 27939 32351
rect 27939 32317 27948 32351
rect 27896 32308 27948 32317
rect 28264 32308 28316 32360
rect 28448 32308 28500 32360
rect 28356 32240 28408 32292
rect 29276 32308 29328 32360
rect 32128 32308 32180 32360
rect 35072 32376 35124 32428
rect 35164 32419 35216 32428
rect 35164 32385 35173 32419
rect 35173 32385 35207 32419
rect 35207 32385 35216 32419
rect 35164 32376 35216 32385
rect 37648 32444 37700 32496
rect 37924 32444 37976 32496
rect 36268 32376 36320 32428
rect 40316 32512 40368 32564
rect 41328 32512 41380 32564
rect 49148 32512 49200 32564
rect 39672 32444 39724 32496
rect 42524 32376 42576 32428
rect 48780 32419 48832 32428
rect 48780 32385 48789 32419
rect 48789 32385 48823 32419
rect 48823 32385 48832 32419
rect 48780 32376 48832 32385
rect 36084 32308 36136 32360
rect 42064 32308 42116 32360
rect 48504 32351 48556 32360
rect 48504 32317 48513 32351
rect 48513 32317 48547 32351
rect 48547 32317 48556 32351
rect 48504 32308 48556 32317
rect 29184 32240 29236 32292
rect 32220 32172 32272 32224
rect 34520 32172 34572 32224
rect 39304 32240 39356 32292
rect 37832 32172 37884 32224
rect 39672 32172 39724 32224
rect 45284 32240 45336 32292
rect 40960 32172 41012 32224
rect 42800 32215 42852 32224
rect 42800 32181 42809 32215
rect 42809 32181 42843 32215
rect 42843 32181 42852 32215
rect 42800 32172 42852 32181
rect 44824 32215 44876 32224
rect 44824 32181 44833 32215
rect 44833 32181 44867 32215
rect 44867 32181 44876 32215
rect 44824 32172 44876 32181
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 32950 32070 33002 32122
rect 33014 32070 33066 32122
rect 33078 32070 33130 32122
rect 33142 32070 33194 32122
rect 33206 32070 33258 32122
rect 42950 32070 43002 32122
rect 43014 32070 43066 32122
rect 43078 32070 43130 32122
rect 43142 32070 43194 32122
rect 43206 32070 43258 32122
rect 22652 31968 22704 32020
rect 24032 32011 24084 32020
rect 24032 31977 24041 32011
rect 24041 31977 24075 32011
rect 24075 31977 24084 32011
rect 24032 31968 24084 31977
rect 23756 31900 23808 31952
rect 23940 31832 23992 31884
rect 24032 31832 24084 31884
rect 27068 31968 27120 32020
rect 27528 32011 27580 32020
rect 27528 31977 27537 32011
rect 27537 31977 27571 32011
rect 27571 31977 27580 32011
rect 27528 31968 27580 31977
rect 27804 31968 27856 32020
rect 27160 31900 27212 31952
rect 35900 31968 35952 32020
rect 38476 31968 38528 32020
rect 39764 31968 39816 32020
rect 40960 31968 41012 32020
rect 26056 31875 26108 31884
rect 26056 31841 26065 31875
rect 26065 31841 26099 31875
rect 26099 31841 26108 31875
rect 26056 31832 26108 31841
rect 32220 31900 32272 31952
rect 29000 31875 29052 31884
rect 29000 31841 29009 31875
rect 29009 31841 29043 31875
rect 29043 31841 29052 31875
rect 29000 31832 29052 31841
rect 32772 31875 32824 31884
rect 32772 31841 32781 31875
rect 32781 31841 32815 31875
rect 32815 31841 32824 31875
rect 32772 31832 32824 31841
rect 35072 31900 35124 31952
rect 36360 31900 36412 31952
rect 40500 31900 40552 31952
rect 40592 31900 40644 31952
rect 43352 31900 43404 31952
rect 23664 31764 23716 31816
rect 23848 31764 23900 31816
rect 27528 31764 27580 31816
rect 31668 31764 31720 31816
rect 36084 31875 36136 31884
rect 36084 31841 36093 31875
rect 36093 31841 36127 31875
rect 36127 31841 36136 31875
rect 36084 31832 36136 31841
rect 34704 31764 34756 31816
rect 34980 31764 35032 31816
rect 35716 31764 35768 31816
rect 37280 31832 37332 31884
rect 37464 31832 37516 31884
rect 38476 31875 38528 31884
rect 38476 31841 38485 31875
rect 38485 31841 38519 31875
rect 38519 31841 38528 31875
rect 38476 31832 38528 31841
rect 24860 31696 24912 31748
rect 23204 31628 23256 31680
rect 25688 31628 25740 31680
rect 26516 31696 26568 31748
rect 30288 31696 30340 31748
rect 30380 31696 30432 31748
rect 35624 31696 35676 31748
rect 39304 31764 39356 31816
rect 38660 31696 38712 31748
rect 27712 31628 27764 31680
rect 28724 31628 28776 31680
rect 35440 31671 35492 31680
rect 35440 31637 35449 31671
rect 35449 31637 35483 31671
rect 35483 31637 35492 31671
rect 35440 31628 35492 31637
rect 37096 31628 37148 31680
rect 37372 31628 37424 31680
rect 37924 31628 37976 31680
rect 39672 31628 39724 31680
rect 40316 31832 40368 31884
rect 42708 31832 42760 31884
rect 48504 31807 48556 31816
rect 48504 31773 48513 31807
rect 48513 31773 48547 31807
rect 48547 31773 48556 31807
rect 48504 31764 48556 31773
rect 42616 31696 42668 31748
rect 41788 31628 41840 31680
rect 42248 31628 42300 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 27950 31526 28002 31578
rect 28014 31526 28066 31578
rect 28078 31526 28130 31578
rect 28142 31526 28194 31578
rect 28206 31526 28258 31578
rect 37950 31526 38002 31578
rect 38014 31526 38066 31578
rect 38078 31526 38130 31578
rect 38142 31526 38194 31578
rect 38206 31526 38258 31578
rect 47950 31526 48002 31578
rect 48014 31526 48066 31578
rect 48078 31526 48130 31578
rect 48142 31526 48194 31578
rect 48206 31526 48258 31578
rect 23848 31467 23900 31476
rect 23848 31433 23857 31467
rect 23857 31433 23891 31467
rect 23891 31433 23900 31467
rect 23848 31424 23900 31433
rect 23940 31424 23992 31476
rect 28908 31424 28960 31476
rect 23480 31356 23532 31408
rect 24768 31356 24820 31408
rect 22836 31288 22888 31340
rect 23296 31288 23348 31340
rect 26240 31288 26292 31340
rect 26516 31288 26568 31340
rect 27160 31288 27212 31340
rect 33876 31288 33928 31340
rect 36268 31424 36320 31476
rect 35808 31356 35860 31408
rect 36544 31356 36596 31408
rect 38200 31356 38252 31408
rect 39304 31424 39356 31476
rect 39488 31424 39540 31476
rect 42800 31424 42852 31476
rect 47860 31424 47912 31476
rect 42432 31356 42484 31408
rect 45744 31356 45796 31408
rect 37740 31331 37792 31340
rect 37740 31297 37749 31331
rect 37749 31297 37783 31331
rect 37783 31297 37792 31331
rect 37740 31288 37792 31297
rect 38384 31288 38436 31340
rect 22468 31263 22520 31272
rect 22468 31229 22477 31263
rect 22477 31229 22511 31263
rect 22511 31229 22520 31263
rect 22468 31220 22520 31229
rect 21824 31084 21876 31136
rect 23204 31084 23256 31136
rect 24124 31263 24176 31272
rect 24124 31229 24133 31263
rect 24133 31229 24167 31263
rect 24167 31229 24176 31263
rect 24124 31220 24176 31229
rect 24584 31220 24636 31272
rect 27528 31220 27580 31272
rect 31668 31220 31720 31272
rect 24676 31152 24728 31204
rect 24952 31084 25004 31136
rect 25780 31084 25832 31136
rect 30380 31084 30432 31136
rect 32864 31084 32916 31136
rect 34060 31220 34112 31272
rect 35532 31220 35584 31272
rect 36360 31220 36412 31272
rect 36452 31220 36504 31272
rect 39028 31288 39080 31340
rect 42064 31288 42116 31340
rect 33416 31152 33468 31204
rect 38476 31152 38528 31204
rect 42156 31220 42208 31272
rect 44272 31288 44324 31340
rect 47400 31288 47452 31340
rect 44364 31220 44416 31272
rect 48504 31263 48556 31272
rect 48504 31229 48513 31263
rect 48513 31229 48547 31263
rect 48547 31229 48556 31263
rect 48504 31220 48556 31229
rect 46020 31152 46072 31204
rect 37004 31084 37056 31136
rect 37556 31127 37608 31136
rect 37556 31093 37565 31127
rect 37565 31093 37599 31127
rect 37599 31093 37608 31127
rect 37556 31084 37608 31093
rect 40408 31084 40460 31136
rect 40776 31084 40828 31136
rect 46940 31084 46992 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 32950 30982 33002 31034
rect 33014 30982 33066 31034
rect 33078 30982 33130 31034
rect 33142 30982 33194 31034
rect 33206 30982 33258 31034
rect 42950 30982 43002 31034
rect 43014 30982 43066 31034
rect 43078 30982 43130 31034
rect 43142 30982 43194 31034
rect 43206 30982 43258 31034
rect 22744 30880 22796 30932
rect 22100 30787 22152 30796
rect 22100 30753 22109 30787
rect 22109 30753 22143 30787
rect 22143 30753 22152 30787
rect 22100 30744 22152 30753
rect 22836 30855 22888 30864
rect 22836 30821 22845 30855
rect 22845 30821 22879 30855
rect 22879 30821 22888 30855
rect 22836 30812 22888 30821
rect 25136 30880 25188 30932
rect 24124 30812 24176 30864
rect 23940 30787 23992 30796
rect 23940 30753 23949 30787
rect 23949 30753 23983 30787
rect 23983 30753 23992 30787
rect 23940 30744 23992 30753
rect 24768 30744 24820 30796
rect 28356 30880 28408 30932
rect 21824 30719 21876 30728
rect 21824 30685 21833 30719
rect 21833 30685 21867 30719
rect 21867 30685 21876 30719
rect 21824 30676 21876 30685
rect 23388 30676 23440 30728
rect 24584 30676 24636 30728
rect 26240 30676 26292 30728
rect 27068 30787 27120 30796
rect 27068 30753 27077 30787
rect 27077 30753 27111 30787
rect 27111 30753 27120 30787
rect 27068 30744 27120 30753
rect 30288 30787 30340 30796
rect 30288 30753 30297 30787
rect 30297 30753 30331 30787
rect 30331 30753 30340 30787
rect 30288 30744 30340 30753
rect 32128 30744 32180 30796
rect 32312 30744 32364 30796
rect 36176 30880 36228 30932
rect 22192 30608 22244 30660
rect 24860 30608 24912 30660
rect 25136 30651 25188 30660
rect 25136 30617 25145 30651
rect 25145 30617 25179 30651
rect 25179 30617 25188 30651
rect 25136 30608 25188 30617
rect 27344 30651 27396 30660
rect 27344 30617 27353 30651
rect 27353 30617 27387 30651
rect 27387 30617 27396 30651
rect 27344 30608 27396 30617
rect 9220 30540 9272 30592
rect 21824 30540 21876 30592
rect 23572 30540 23624 30592
rect 25412 30540 25464 30592
rect 30380 30676 30432 30728
rect 31300 30719 31352 30728
rect 31300 30685 31309 30719
rect 31309 30685 31343 30719
rect 31343 30685 31352 30719
rect 31300 30676 31352 30685
rect 34796 30676 34848 30728
rect 34980 30676 35032 30728
rect 35900 30812 35952 30864
rect 35992 30812 36044 30864
rect 36544 30812 36596 30864
rect 38936 30812 38988 30864
rect 39488 30880 39540 30932
rect 41880 30880 41932 30932
rect 47676 30880 47728 30932
rect 35716 30744 35768 30796
rect 36912 30787 36964 30796
rect 36912 30753 36921 30787
rect 36921 30753 36955 30787
rect 36955 30753 36964 30787
rect 36912 30744 36964 30753
rect 37004 30744 37056 30796
rect 38752 30744 38804 30796
rect 39396 30744 39448 30796
rect 40500 30787 40552 30796
rect 40500 30753 40509 30787
rect 40509 30753 40543 30787
rect 40543 30753 40552 30787
rect 40500 30744 40552 30753
rect 40592 30787 40644 30796
rect 40592 30753 40601 30787
rect 40601 30753 40635 30787
rect 40635 30753 40644 30787
rect 40592 30744 40644 30753
rect 39488 30676 39540 30728
rect 40408 30719 40460 30728
rect 40408 30685 40417 30719
rect 40417 30685 40451 30719
rect 40451 30685 40460 30719
rect 40408 30676 40460 30685
rect 41512 30812 41564 30864
rect 42156 30719 42208 30728
rect 42156 30685 42165 30719
rect 42165 30685 42199 30719
rect 42199 30685 42208 30719
rect 42156 30676 42208 30685
rect 31576 30651 31628 30660
rect 28816 30583 28868 30592
rect 28816 30549 28825 30583
rect 28825 30549 28859 30583
rect 28859 30549 28868 30583
rect 28816 30540 28868 30549
rect 28908 30540 28960 30592
rect 31576 30617 31585 30651
rect 31585 30617 31619 30651
rect 31619 30617 31628 30651
rect 31576 30608 31628 30617
rect 32404 30540 32456 30592
rect 32588 30540 32640 30592
rect 34612 30608 34664 30660
rect 34796 30540 34848 30592
rect 36544 30540 36596 30592
rect 37096 30540 37148 30592
rect 41236 30608 41288 30660
rect 37740 30583 37792 30592
rect 37740 30549 37749 30583
rect 37749 30549 37783 30583
rect 37783 30549 37792 30583
rect 37740 30540 37792 30549
rect 38752 30540 38804 30592
rect 40040 30583 40092 30592
rect 40040 30549 40049 30583
rect 40049 30549 40083 30583
rect 40083 30549 40092 30583
rect 40040 30540 40092 30549
rect 46112 30608 46164 30660
rect 48688 30651 48740 30660
rect 48688 30617 48697 30651
rect 48697 30617 48731 30651
rect 48731 30617 48740 30651
rect 48688 30608 48740 30617
rect 41972 30583 42024 30592
rect 41972 30549 41981 30583
rect 41981 30549 42015 30583
rect 42015 30549 42024 30583
rect 41972 30540 42024 30549
rect 47032 30540 47084 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 27950 30438 28002 30490
rect 28014 30438 28066 30490
rect 28078 30438 28130 30490
rect 28142 30438 28194 30490
rect 28206 30438 28258 30490
rect 37950 30438 38002 30490
rect 38014 30438 38066 30490
rect 38078 30438 38130 30490
rect 38142 30438 38194 30490
rect 38206 30438 38258 30490
rect 47950 30438 48002 30490
rect 48014 30438 48066 30490
rect 48078 30438 48130 30490
rect 48142 30438 48194 30490
rect 48206 30438 48258 30490
rect 24768 30268 24820 30320
rect 26056 30311 26108 30320
rect 26056 30277 26065 30311
rect 26065 30277 26099 30311
rect 26099 30277 26108 30311
rect 26056 30268 26108 30277
rect 7380 30243 7432 30252
rect 7380 30209 7389 30243
rect 7389 30209 7423 30243
rect 7423 30209 7432 30243
rect 7380 30200 7432 30209
rect 21180 30200 21232 30252
rect 25504 30200 25556 30252
rect 25596 30200 25648 30252
rect 7656 30132 7708 30184
rect 9128 30175 9180 30184
rect 9128 30141 9137 30175
rect 9137 30141 9171 30175
rect 9171 30141 9180 30175
rect 9128 30132 9180 30141
rect 23572 30175 23624 30184
rect 23572 30141 23581 30175
rect 23581 30141 23615 30175
rect 23615 30141 23624 30175
rect 23572 30132 23624 30141
rect 27528 30132 27580 30184
rect 28724 30200 28776 30252
rect 30472 30336 30524 30388
rect 36912 30336 36964 30388
rect 37464 30336 37516 30388
rect 38384 30336 38436 30388
rect 41236 30336 41288 30388
rect 30012 30268 30064 30320
rect 31300 30268 31352 30320
rect 30472 30200 30524 30252
rect 33692 30268 33744 30320
rect 18696 30064 18748 30116
rect 26332 30064 26384 30116
rect 27436 30064 27488 30116
rect 29460 30132 29512 30184
rect 32128 30200 32180 30252
rect 34152 30243 34204 30252
rect 34152 30209 34161 30243
rect 34161 30209 34195 30243
rect 34195 30209 34204 30243
rect 34152 30200 34204 30209
rect 33968 30132 34020 30184
rect 35808 30268 35860 30320
rect 36084 30268 36136 30320
rect 37832 30311 37884 30320
rect 37832 30277 37841 30311
rect 37841 30277 37875 30311
rect 37875 30277 37884 30311
rect 37832 30268 37884 30277
rect 38292 30268 38344 30320
rect 38476 30268 38528 30320
rect 34428 30200 34480 30252
rect 37188 30200 37240 30252
rect 41696 30200 41748 30252
rect 42616 30200 42668 30252
rect 49332 30243 49384 30252
rect 49332 30209 49341 30243
rect 49341 30209 49375 30243
rect 49375 30209 49384 30243
rect 49332 30200 49384 30209
rect 28632 29996 28684 30048
rect 33876 30064 33928 30116
rect 34060 30064 34112 30116
rect 34612 30064 34664 30116
rect 36268 30064 36320 30116
rect 40684 30132 40736 30184
rect 40868 30132 40920 30184
rect 40132 30064 40184 30116
rect 41328 30064 41380 30116
rect 32772 29996 32824 30048
rect 35164 29996 35216 30048
rect 36176 29996 36228 30048
rect 40500 30039 40552 30048
rect 40500 30005 40509 30039
rect 40509 30005 40543 30039
rect 40543 30005 40552 30039
rect 40500 29996 40552 30005
rect 45744 29996 45796 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 32950 29894 33002 29946
rect 33014 29894 33066 29946
rect 33078 29894 33130 29946
rect 33142 29894 33194 29946
rect 33206 29894 33258 29946
rect 42950 29894 43002 29946
rect 43014 29894 43066 29946
rect 43078 29894 43130 29946
rect 43142 29894 43194 29946
rect 43206 29894 43258 29946
rect 10692 29792 10744 29844
rect 25596 29792 25648 29844
rect 28816 29792 28868 29844
rect 1308 29656 1360 29708
rect 21088 29656 21140 29708
rect 27344 29656 27396 29708
rect 27528 29656 27580 29708
rect 29368 29656 29420 29708
rect 30472 29792 30524 29844
rect 32220 29792 32272 29844
rect 34428 29792 34480 29844
rect 34704 29792 34756 29844
rect 35256 29724 35308 29776
rect 36452 29792 36504 29844
rect 42708 29835 42760 29844
rect 42708 29801 42717 29835
rect 42717 29801 42751 29835
rect 42751 29801 42760 29835
rect 42708 29792 42760 29801
rect 4804 29588 4856 29640
rect 27068 29588 27120 29640
rect 30012 29588 30064 29640
rect 30472 29656 30524 29708
rect 33876 29656 33928 29708
rect 34704 29656 34756 29708
rect 36268 29656 36320 29708
rect 38568 29724 38620 29776
rect 37464 29656 37516 29708
rect 39764 29656 39816 29708
rect 40316 29656 40368 29708
rect 40684 29656 40736 29708
rect 34244 29588 34296 29640
rect 40776 29588 40828 29640
rect 48504 29631 48556 29640
rect 48504 29597 48513 29631
rect 48513 29597 48547 29631
rect 48547 29597 48556 29631
rect 48504 29588 48556 29597
rect 21180 29563 21232 29572
rect 21180 29529 21189 29563
rect 21189 29529 21223 29563
rect 21223 29529 21232 29563
rect 21180 29520 21232 29529
rect 28540 29520 28592 29572
rect 28724 29520 28776 29572
rect 29460 29520 29512 29572
rect 22744 29452 22796 29504
rect 23664 29452 23716 29504
rect 36636 29520 36688 29572
rect 37280 29520 37332 29572
rect 40500 29520 40552 29572
rect 41696 29520 41748 29572
rect 29920 29452 29972 29504
rect 31944 29495 31996 29504
rect 31944 29461 31953 29495
rect 31953 29461 31987 29495
rect 31987 29461 31996 29495
rect 31944 29452 31996 29461
rect 32404 29495 32456 29504
rect 32404 29461 32413 29495
rect 32413 29461 32447 29495
rect 32447 29461 32456 29495
rect 32404 29452 32456 29461
rect 35900 29452 35952 29504
rect 36268 29452 36320 29504
rect 41420 29452 41472 29504
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 27950 29350 28002 29402
rect 28014 29350 28066 29402
rect 28078 29350 28130 29402
rect 28142 29350 28194 29402
rect 28206 29350 28258 29402
rect 37950 29350 38002 29402
rect 38014 29350 38066 29402
rect 38078 29350 38130 29402
rect 38142 29350 38194 29402
rect 38206 29350 38258 29402
rect 47950 29350 48002 29402
rect 48014 29350 48066 29402
rect 48078 29350 48130 29402
rect 48142 29350 48194 29402
rect 48206 29350 48258 29402
rect 23296 29248 23348 29300
rect 17224 29180 17276 29232
rect 28816 29248 28868 29300
rect 30104 29248 30156 29300
rect 30472 29248 30524 29300
rect 34152 29248 34204 29300
rect 34428 29248 34480 29300
rect 35532 29248 35584 29300
rect 40040 29248 40092 29300
rect 22376 29155 22428 29164
rect 22376 29121 22385 29155
rect 22385 29121 22419 29155
rect 22419 29121 22428 29155
rect 22376 29112 22428 29121
rect 29736 29180 29788 29232
rect 33508 29180 33560 29232
rect 33784 29180 33836 29232
rect 34796 29180 34848 29232
rect 37648 29180 37700 29232
rect 41328 29180 41380 29232
rect 23296 29155 23348 29164
rect 23296 29121 23305 29155
rect 23305 29121 23339 29155
rect 23339 29121 23348 29155
rect 23296 29112 23348 29121
rect 27068 29112 27120 29164
rect 29276 29112 29328 29164
rect 29552 29112 29604 29164
rect 32404 29112 32456 29164
rect 41144 29155 41196 29164
rect 41144 29121 41153 29155
rect 41153 29121 41187 29155
rect 41187 29121 41196 29155
rect 41144 29112 41196 29121
rect 25136 29044 25188 29096
rect 7748 28976 7800 29028
rect 22376 28976 22428 29028
rect 25688 28976 25740 29028
rect 26148 28976 26200 29028
rect 29000 28976 29052 29028
rect 30472 29087 30524 29096
rect 30472 29053 30481 29087
rect 30481 29053 30515 29087
rect 30515 29053 30524 29087
rect 30472 29044 30524 29053
rect 33968 29087 34020 29096
rect 33968 29053 33977 29087
rect 33977 29053 34011 29087
rect 34011 29053 34020 29087
rect 33968 29044 34020 29053
rect 37280 29044 37332 29096
rect 37832 29044 37884 29096
rect 38660 29044 38712 29096
rect 39028 29044 39080 29096
rect 42708 29044 42760 29096
rect 28540 28908 28592 28960
rect 29460 28951 29512 28960
rect 29460 28917 29469 28951
rect 29469 28917 29503 28951
rect 29503 28917 29512 28951
rect 29460 28908 29512 28917
rect 32128 28976 32180 29028
rect 35808 28976 35860 29028
rect 39396 28976 39448 29028
rect 44180 28976 44232 29028
rect 49332 29155 49384 29164
rect 49332 29121 49341 29155
rect 49341 29121 49375 29155
rect 49375 29121 49384 29155
rect 49332 29112 49384 29121
rect 32036 28908 32088 28960
rect 32588 28908 32640 28960
rect 36268 28908 36320 28960
rect 36360 28951 36412 28960
rect 36360 28917 36369 28951
rect 36369 28917 36403 28951
rect 36403 28917 36412 28951
rect 36360 28908 36412 28917
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 32950 28806 33002 28858
rect 33014 28806 33066 28858
rect 33078 28806 33130 28858
rect 33142 28806 33194 28858
rect 33206 28806 33258 28858
rect 42950 28806 43002 28858
rect 43014 28806 43066 28858
rect 43078 28806 43130 28858
rect 43142 28806 43194 28858
rect 43206 28806 43258 28858
rect 22192 28747 22244 28756
rect 22192 28713 22201 28747
rect 22201 28713 22235 28747
rect 22235 28713 22244 28747
rect 22192 28704 22244 28713
rect 35440 28704 35492 28756
rect 39120 28704 39172 28756
rect 27620 28636 27672 28688
rect 28816 28636 28868 28688
rect 22560 28568 22612 28620
rect 23388 28568 23440 28620
rect 29460 28568 29512 28620
rect 32864 28568 32916 28620
rect 34152 28611 34204 28620
rect 34152 28577 34161 28611
rect 34161 28577 34195 28611
rect 34195 28577 34204 28611
rect 34152 28568 34204 28577
rect 24952 28500 25004 28552
rect 27620 28500 27672 28552
rect 29920 28543 29972 28552
rect 29920 28509 29929 28543
rect 29929 28509 29963 28543
rect 29963 28509 29972 28543
rect 29920 28500 29972 28509
rect 33324 28500 33376 28552
rect 33784 28500 33836 28552
rect 36820 28636 36872 28688
rect 39212 28636 39264 28688
rect 39488 28636 39540 28688
rect 35808 28568 35860 28620
rect 36268 28568 36320 28620
rect 38292 28568 38344 28620
rect 36360 28500 36412 28552
rect 40224 28568 40276 28620
rect 40684 28611 40736 28620
rect 40684 28577 40693 28611
rect 40693 28577 40727 28611
rect 40727 28577 40736 28611
rect 40684 28568 40736 28577
rect 39028 28500 39080 28552
rect 41052 28500 41104 28552
rect 49332 28543 49384 28552
rect 49332 28509 49341 28543
rect 49341 28509 49375 28543
rect 49375 28509 49384 28543
rect 49332 28500 49384 28509
rect 7104 28364 7156 28416
rect 19340 28364 19392 28416
rect 25504 28475 25556 28484
rect 25504 28441 25513 28475
rect 25513 28441 25547 28475
rect 25547 28441 25556 28475
rect 25504 28432 25556 28441
rect 27068 28475 27120 28484
rect 27068 28441 27077 28475
rect 27077 28441 27111 28475
rect 27111 28441 27120 28475
rect 27068 28432 27120 28441
rect 30196 28432 30248 28484
rect 22560 28407 22612 28416
rect 22560 28373 22569 28407
rect 22569 28373 22603 28407
rect 22603 28373 22612 28407
rect 22560 28364 22612 28373
rect 28356 28407 28408 28416
rect 28356 28373 28365 28407
rect 28365 28373 28399 28407
rect 28399 28373 28408 28407
rect 28356 28364 28408 28373
rect 31116 28364 31168 28416
rect 35164 28432 35216 28484
rect 38936 28432 38988 28484
rect 31300 28364 31352 28416
rect 32864 28364 32916 28416
rect 35072 28364 35124 28416
rect 35256 28407 35308 28416
rect 35256 28373 35265 28407
rect 35265 28373 35299 28407
rect 35299 28373 35308 28407
rect 35256 28364 35308 28373
rect 35440 28364 35492 28416
rect 36084 28407 36136 28416
rect 36084 28373 36093 28407
rect 36093 28373 36127 28407
rect 36127 28373 36136 28407
rect 36084 28364 36136 28373
rect 36544 28407 36596 28416
rect 36544 28373 36553 28407
rect 36553 28373 36587 28407
rect 36587 28373 36596 28407
rect 36544 28364 36596 28373
rect 37280 28407 37332 28416
rect 37280 28373 37289 28407
rect 37289 28373 37323 28407
rect 37323 28373 37332 28407
rect 37280 28364 37332 28373
rect 40224 28364 40276 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 27950 28262 28002 28314
rect 28014 28262 28066 28314
rect 28078 28262 28130 28314
rect 28142 28262 28194 28314
rect 28206 28262 28258 28314
rect 37950 28262 38002 28314
rect 38014 28262 38066 28314
rect 38078 28262 38130 28314
rect 38142 28262 38194 28314
rect 38206 28262 38258 28314
rect 47950 28262 48002 28314
rect 48014 28262 48066 28314
rect 48078 28262 48130 28314
rect 48142 28262 48194 28314
rect 48206 28262 48258 28314
rect 4804 28203 4856 28212
rect 4804 28169 4813 28203
rect 4813 28169 4847 28203
rect 4847 28169 4856 28203
rect 4804 28160 4856 28169
rect 21180 28092 21232 28144
rect 7564 28067 7616 28076
rect 7564 28033 7573 28067
rect 7573 28033 7607 28067
rect 7607 28033 7616 28067
rect 7564 28024 7616 28033
rect 22100 28024 22152 28076
rect 23848 28024 23900 28076
rect 24952 28092 25004 28144
rect 26240 28092 26292 28144
rect 7748 27999 7800 28008
rect 7748 27965 7757 27999
rect 7757 27965 7791 27999
rect 7791 27965 7800 27999
rect 7748 27956 7800 27965
rect 9496 27956 9548 28008
rect 21456 27956 21508 28008
rect 23388 27956 23440 28008
rect 9680 27888 9732 27940
rect 24216 27863 24268 27872
rect 24216 27829 24225 27863
rect 24225 27829 24259 27863
rect 24259 27829 24268 27863
rect 24216 27820 24268 27829
rect 26700 27956 26752 28008
rect 30288 28160 30340 28212
rect 32128 28160 32180 28212
rect 27804 28092 27856 28144
rect 28540 28092 28592 28144
rect 29736 28092 29788 28144
rect 30196 28092 30248 28144
rect 29552 28024 29604 28076
rect 27620 27956 27672 28008
rect 29736 27956 29788 28008
rect 30748 27956 30800 28008
rect 32036 28092 32088 28144
rect 33416 28160 33468 28212
rect 35900 28160 35952 28212
rect 36544 28160 36596 28212
rect 38660 28160 38712 28212
rect 39028 28203 39080 28212
rect 39028 28169 39037 28203
rect 39037 28169 39071 28203
rect 39071 28169 39080 28203
rect 39028 28160 39080 28169
rect 33876 28092 33928 28144
rect 34796 28092 34848 28144
rect 36820 28092 36872 28144
rect 37464 28024 37516 28076
rect 28448 27820 28500 27872
rect 28632 27820 28684 27872
rect 29828 27820 29880 27872
rect 32312 27999 32364 28008
rect 32312 27965 32321 27999
rect 32321 27965 32355 27999
rect 32355 27965 32364 27999
rect 32312 27956 32364 27965
rect 34520 27956 34572 28008
rect 37648 27956 37700 28008
rect 38476 28024 38528 28076
rect 38660 28024 38712 28076
rect 39488 28024 39540 28076
rect 46940 28092 46992 28144
rect 41604 28024 41656 28076
rect 39120 27999 39172 28008
rect 39120 27965 39129 27999
rect 39129 27965 39163 27999
rect 39163 27965 39172 27999
rect 39120 27956 39172 27965
rect 40500 27956 40552 28008
rect 33784 27888 33836 27940
rect 38384 27888 38436 27940
rect 41144 27888 41196 27940
rect 32588 27820 32640 27872
rect 34152 27820 34204 27872
rect 35164 27820 35216 27872
rect 35440 27820 35492 27872
rect 35992 27863 36044 27872
rect 35992 27829 36001 27863
rect 36001 27829 36035 27863
rect 36035 27829 36044 27863
rect 35992 27820 36044 27829
rect 37188 27820 37240 27872
rect 41236 27820 41288 27872
rect 47768 27820 47820 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 32950 27718 33002 27770
rect 33014 27718 33066 27770
rect 33078 27718 33130 27770
rect 33142 27718 33194 27770
rect 33206 27718 33258 27770
rect 42950 27718 43002 27770
rect 43014 27718 43066 27770
rect 43078 27718 43130 27770
rect 43142 27718 43194 27770
rect 43206 27718 43258 27770
rect 28356 27616 28408 27668
rect 30656 27616 30708 27668
rect 30748 27616 30800 27668
rect 39120 27616 39172 27668
rect 40776 27616 40828 27668
rect 7656 27548 7708 27600
rect 29552 27548 29604 27600
rect 1308 27480 1360 27532
rect 24952 27523 25004 27532
rect 24952 27489 24961 27523
rect 24961 27489 24995 27523
rect 24995 27489 25004 27523
rect 24952 27480 25004 27489
rect 30288 27480 30340 27532
rect 4988 27412 5040 27464
rect 4896 27344 4948 27396
rect 9772 27412 9824 27464
rect 23112 27412 23164 27464
rect 29920 27412 29972 27464
rect 25228 27387 25280 27396
rect 25228 27353 25237 27387
rect 25237 27353 25271 27387
rect 25271 27353 25280 27387
rect 25228 27344 25280 27353
rect 26240 27344 26292 27396
rect 27620 27344 27672 27396
rect 32772 27548 32824 27600
rect 32036 27480 32088 27532
rect 32220 27480 32272 27532
rect 35348 27523 35400 27532
rect 35348 27489 35357 27523
rect 35357 27489 35391 27523
rect 35391 27489 35400 27523
rect 35348 27480 35400 27489
rect 35532 27523 35584 27532
rect 35532 27489 35541 27523
rect 35541 27489 35575 27523
rect 35575 27489 35584 27523
rect 35532 27480 35584 27489
rect 41604 27548 41656 27600
rect 34888 27412 34940 27464
rect 36084 27412 36136 27464
rect 40316 27480 40368 27532
rect 31484 27344 31536 27396
rect 26700 27319 26752 27328
rect 26700 27285 26709 27319
rect 26709 27285 26743 27319
rect 26743 27285 26752 27319
rect 26700 27276 26752 27285
rect 27252 27276 27304 27328
rect 28540 27276 28592 27328
rect 30196 27319 30248 27328
rect 30196 27285 30205 27319
rect 30205 27285 30239 27319
rect 30239 27285 30248 27319
rect 30196 27276 30248 27285
rect 30656 27319 30708 27328
rect 30656 27285 30665 27319
rect 30665 27285 30699 27319
rect 30699 27285 30708 27319
rect 30656 27276 30708 27285
rect 30748 27276 30800 27328
rect 32312 27344 32364 27396
rect 33968 27344 34020 27396
rect 37188 27344 37240 27396
rect 37924 27344 37976 27396
rect 41420 27412 41472 27464
rect 31760 27319 31812 27328
rect 31760 27285 31769 27319
rect 31769 27285 31803 27319
rect 31803 27285 31812 27319
rect 31760 27276 31812 27285
rect 32588 27276 32640 27328
rect 34796 27276 34848 27328
rect 35900 27276 35952 27328
rect 36084 27276 36136 27328
rect 38292 27276 38344 27328
rect 47124 27480 47176 27532
rect 44180 27455 44232 27464
rect 44180 27421 44189 27455
rect 44189 27421 44223 27455
rect 44223 27421 44232 27455
rect 44180 27412 44232 27421
rect 47216 27455 47268 27464
rect 47216 27421 47225 27455
rect 47225 27421 47259 27455
rect 47259 27421 47268 27455
rect 47216 27412 47268 27421
rect 48504 27455 48556 27464
rect 48504 27421 48513 27455
rect 48513 27421 48547 27455
rect 48547 27421 48556 27455
rect 48504 27412 48556 27421
rect 47584 27344 47636 27396
rect 47676 27344 47728 27396
rect 43996 27319 44048 27328
rect 43996 27285 44005 27319
rect 44005 27285 44039 27319
rect 44039 27285 44048 27319
rect 43996 27276 44048 27285
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 27950 27174 28002 27226
rect 28014 27174 28066 27226
rect 28078 27174 28130 27226
rect 28142 27174 28194 27226
rect 28206 27174 28258 27226
rect 37950 27174 38002 27226
rect 38014 27174 38066 27226
rect 38078 27174 38130 27226
rect 38142 27174 38194 27226
rect 38206 27174 38258 27226
rect 47950 27174 48002 27226
rect 48014 27174 48066 27226
rect 48078 27174 48130 27226
rect 48142 27174 48194 27226
rect 48206 27174 48258 27226
rect 23112 27115 23164 27124
rect 23112 27081 23121 27115
rect 23121 27081 23155 27115
rect 23155 27081 23164 27115
rect 23112 27072 23164 27081
rect 26700 27072 26752 27124
rect 27160 27072 27212 27124
rect 30656 27072 30708 27124
rect 30840 27072 30892 27124
rect 31208 27072 31260 27124
rect 31852 27072 31904 27124
rect 22560 27004 22612 27056
rect 25872 27004 25924 27056
rect 33876 27004 33928 27056
rect 34980 27004 35032 27056
rect 7840 26979 7892 26988
rect 7840 26945 7849 26979
rect 7849 26945 7883 26979
rect 7883 26945 7892 26979
rect 7840 26936 7892 26945
rect 30288 26936 30340 26988
rect 31300 26936 31352 26988
rect 37096 27072 37148 27124
rect 40592 27072 40644 27124
rect 40684 27072 40736 27124
rect 42156 27072 42208 27124
rect 48780 27072 48832 27124
rect 41604 27004 41656 27056
rect 44824 27004 44876 27056
rect 37740 26979 37792 26988
rect 37740 26945 37749 26979
rect 37749 26945 37783 26979
rect 37783 26945 37792 26979
rect 37740 26936 37792 26945
rect 39856 26936 39908 26988
rect 40316 26979 40368 26988
rect 40316 26945 40332 26979
rect 40332 26945 40366 26979
rect 40366 26945 40368 26979
rect 40316 26936 40368 26945
rect 47032 26979 47084 26988
rect 47032 26945 47041 26979
rect 47041 26945 47075 26979
rect 47075 26945 47084 26979
rect 47032 26936 47084 26945
rect 47124 26936 47176 26988
rect 8300 26868 8352 26920
rect 9588 26911 9640 26920
rect 9588 26877 9597 26911
rect 9597 26877 9631 26911
rect 9631 26877 9640 26911
rect 9588 26868 9640 26877
rect 23388 26911 23440 26920
rect 23388 26877 23397 26911
rect 23397 26877 23431 26911
rect 23431 26877 23440 26911
rect 23388 26868 23440 26877
rect 28448 26868 28500 26920
rect 29828 26868 29880 26920
rect 28172 26800 28224 26852
rect 31024 26868 31076 26920
rect 31392 26911 31444 26920
rect 31392 26877 31401 26911
rect 31401 26877 31435 26911
rect 31435 26877 31444 26911
rect 31392 26868 31444 26877
rect 33232 26868 33284 26920
rect 34060 26868 34112 26920
rect 31484 26800 31536 26852
rect 34152 26800 34204 26852
rect 24032 26732 24084 26784
rect 26976 26732 27028 26784
rect 30104 26732 30156 26784
rect 30380 26732 30432 26784
rect 31300 26732 31352 26784
rect 33968 26732 34020 26784
rect 40132 26868 40184 26920
rect 35808 26800 35860 26852
rect 34980 26732 35032 26784
rect 36084 26732 36136 26784
rect 39028 26732 39080 26784
rect 47676 26868 47728 26920
rect 48504 26911 48556 26920
rect 48504 26877 48513 26911
rect 48513 26877 48547 26911
rect 48547 26877 48556 26911
rect 48504 26868 48556 26877
rect 46756 26732 46808 26784
rect 47676 26732 47728 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 32950 26630 33002 26682
rect 33014 26630 33066 26682
rect 33078 26630 33130 26682
rect 33142 26630 33194 26682
rect 33206 26630 33258 26682
rect 42950 26630 43002 26682
rect 43014 26630 43066 26682
rect 43078 26630 43130 26682
rect 43142 26630 43194 26682
rect 43206 26630 43258 26682
rect 7748 26528 7800 26580
rect 9680 26571 9732 26580
rect 9680 26537 9689 26571
rect 9689 26537 9723 26571
rect 9723 26537 9732 26571
rect 9680 26528 9732 26537
rect 25044 26528 25096 26580
rect 25320 26528 25372 26580
rect 25780 26528 25832 26580
rect 27160 26528 27212 26580
rect 27804 26528 27856 26580
rect 35532 26528 35584 26580
rect 40132 26528 40184 26580
rect 41788 26571 41840 26580
rect 41788 26537 41797 26571
rect 41797 26537 41831 26571
rect 41831 26537 41840 26571
rect 41788 26528 41840 26537
rect 23756 26460 23808 26512
rect 24216 26460 24268 26512
rect 10876 26392 10928 26444
rect 22100 26435 22152 26444
rect 22100 26401 22109 26435
rect 22109 26401 22143 26435
rect 22143 26401 22152 26435
rect 22100 26392 22152 26401
rect 25044 26435 25096 26444
rect 25044 26401 25053 26435
rect 25053 26401 25087 26435
rect 25087 26401 25096 26435
rect 25044 26392 25096 26401
rect 7748 26367 7800 26376
rect 7748 26333 7792 26367
rect 7792 26333 7800 26367
rect 7748 26324 7800 26333
rect 9772 26324 9824 26376
rect 10968 26324 11020 26376
rect 23756 26324 23808 26376
rect 26976 26367 27028 26376
rect 26976 26333 26985 26367
rect 26985 26333 27019 26367
rect 27019 26333 27028 26367
rect 26976 26324 27028 26333
rect 27160 26435 27212 26444
rect 27160 26401 27169 26435
rect 27169 26401 27203 26435
rect 27203 26401 27212 26435
rect 27160 26392 27212 26401
rect 29368 26392 29420 26444
rect 30748 26392 30800 26444
rect 28172 26367 28224 26376
rect 28172 26333 28181 26367
rect 28181 26333 28215 26367
rect 28215 26333 28224 26367
rect 28172 26324 28224 26333
rect 28908 26324 28960 26376
rect 29092 26324 29144 26376
rect 31024 26324 31076 26376
rect 38384 26460 38436 26512
rect 39028 26460 39080 26512
rect 31208 26435 31260 26444
rect 31208 26401 31217 26435
rect 31217 26401 31251 26435
rect 31251 26401 31260 26435
rect 31208 26392 31260 26401
rect 31300 26435 31352 26444
rect 31300 26401 31309 26435
rect 31309 26401 31343 26435
rect 31343 26401 31352 26435
rect 31300 26392 31352 26401
rect 31852 26392 31904 26444
rect 32036 26392 32088 26444
rect 32220 26435 32272 26444
rect 32220 26401 32229 26435
rect 32229 26401 32263 26435
rect 32263 26401 32272 26435
rect 32220 26392 32272 26401
rect 33876 26392 33928 26444
rect 35992 26392 36044 26444
rect 39396 26435 39448 26444
rect 39396 26401 39405 26435
rect 39405 26401 39439 26435
rect 39439 26401 39448 26435
rect 39396 26392 39448 26401
rect 39856 26392 39908 26444
rect 34888 26367 34940 26376
rect 34888 26333 34897 26367
rect 34897 26333 34931 26367
rect 34931 26333 34940 26367
rect 34888 26324 34940 26333
rect 37740 26324 37792 26376
rect 39948 26324 40000 26376
rect 41420 26324 41472 26376
rect 48780 26435 48832 26444
rect 48780 26401 48789 26435
rect 48789 26401 48823 26435
rect 48823 26401 48832 26435
rect 48780 26392 48832 26401
rect 42800 26324 42852 26376
rect 43996 26324 44048 26376
rect 48228 26324 48280 26376
rect 23664 26256 23716 26308
rect 23848 26256 23900 26308
rect 32036 26256 32088 26308
rect 32404 26256 32456 26308
rect 32496 26299 32548 26308
rect 32496 26265 32505 26299
rect 32505 26265 32539 26299
rect 32539 26265 32548 26299
rect 32496 26256 32548 26265
rect 32588 26256 32640 26308
rect 33784 26256 33836 26308
rect 24584 26231 24636 26240
rect 24584 26197 24593 26231
rect 24593 26197 24627 26231
rect 24627 26197 24636 26231
rect 24584 26188 24636 26197
rect 26884 26188 26936 26240
rect 27804 26231 27856 26240
rect 27804 26197 27813 26231
rect 27813 26197 27847 26231
rect 27847 26197 27856 26231
rect 27804 26188 27856 26197
rect 32128 26188 32180 26240
rect 34980 26256 35032 26308
rect 38568 26256 38620 26308
rect 39488 26256 39540 26308
rect 34888 26188 34940 26240
rect 47216 26231 47268 26240
rect 47216 26197 47225 26231
rect 47225 26197 47259 26231
rect 47259 26197 47268 26231
rect 47216 26188 47268 26197
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 27950 26086 28002 26138
rect 28014 26086 28066 26138
rect 28078 26086 28130 26138
rect 28142 26086 28194 26138
rect 28206 26086 28258 26138
rect 37950 26086 38002 26138
rect 38014 26086 38066 26138
rect 38078 26086 38130 26138
rect 38142 26086 38194 26138
rect 38206 26086 38258 26138
rect 47950 26086 48002 26138
rect 48014 26086 48066 26138
rect 48078 26086 48130 26138
rect 48142 26086 48194 26138
rect 48206 26086 48258 26138
rect 26976 25984 27028 26036
rect 29092 25984 29144 26036
rect 32680 26027 32732 26036
rect 32680 25993 32689 26027
rect 32689 25993 32723 26027
rect 32723 25993 32732 26027
rect 32680 25984 32732 25993
rect 38660 25984 38712 26036
rect 38844 25984 38896 26036
rect 39304 25984 39356 26036
rect 40776 25984 40828 26036
rect 30288 25916 30340 25968
rect 32772 25959 32824 25968
rect 32772 25925 32781 25959
rect 32781 25925 32815 25959
rect 32815 25925 32824 25959
rect 32772 25916 32824 25925
rect 34704 25916 34756 25968
rect 35808 25916 35860 25968
rect 38568 25916 38620 25968
rect 7472 25848 7524 25900
rect 30564 25848 30616 25900
rect 34520 25848 34572 25900
rect 9036 25780 9088 25832
rect 9404 25823 9456 25832
rect 9404 25789 9413 25823
rect 9413 25789 9447 25823
rect 9447 25789 9456 25823
rect 9404 25780 9456 25789
rect 22376 25780 22428 25832
rect 25228 25780 25280 25832
rect 28448 25823 28500 25832
rect 28448 25789 28457 25823
rect 28457 25789 28491 25823
rect 28491 25789 28500 25823
rect 28448 25780 28500 25789
rect 26240 25712 26292 25764
rect 30104 25780 30156 25832
rect 32496 25780 32548 25832
rect 32220 25712 32272 25764
rect 34704 25780 34756 25832
rect 36084 25780 36136 25832
rect 37464 25780 37516 25832
rect 37648 25780 37700 25832
rect 40132 25848 40184 25900
rect 40684 25916 40736 25968
rect 46112 25959 46164 25968
rect 46112 25925 46121 25959
rect 46121 25925 46155 25959
rect 46155 25925 46164 25959
rect 46112 25916 46164 25925
rect 41604 25848 41656 25900
rect 39212 25823 39264 25832
rect 39212 25789 39221 25823
rect 39221 25789 39255 25823
rect 39255 25789 39264 25823
rect 39212 25780 39264 25789
rect 37832 25712 37884 25764
rect 39672 25712 39724 25764
rect 25780 25644 25832 25696
rect 25872 25644 25924 25696
rect 27436 25644 27488 25696
rect 28540 25644 28592 25696
rect 29920 25644 29972 25696
rect 31024 25687 31076 25696
rect 31024 25653 31033 25687
rect 31033 25653 31067 25687
rect 31067 25653 31076 25687
rect 31024 25644 31076 25653
rect 36820 25644 36872 25696
rect 36912 25687 36964 25696
rect 36912 25653 36921 25687
rect 36921 25653 36955 25687
rect 36955 25653 36964 25687
rect 36912 25644 36964 25653
rect 37464 25687 37516 25696
rect 37464 25653 37473 25687
rect 37473 25653 37507 25687
rect 37507 25653 37516 25687
rect 37464 25644 37516 25653
rect 38660 25687 38712 25696
rect 38660 25653 38669 25687
rect 38669 25653 38703 25687
rect 38703 25653 38712 25687
rect 38660 25644 38712 25653
rect 39580 25644 39632 25696
rect 41972 25848 42024 25900
rect 49332 25891 49384 25900
rect 49332 25857 49341 25891
rect 49341 25857 49375 25891
rect 49375 25857 49384 25891
rect 49332 25848 49384 25857
rect 46296 25755 46348 25764
rect 46296 25721 46305 25755
rect 46305 25721 46339 25755
rect 46339 25721 46348 25755
rect 46296 25712 46348 25721
rect 47032 25755 47084 25764
rect 47032 25721 47041 25755
rect 47041 25721 47075 25755
rect 47075 25721 47084 25755
rect 47032 25712 47084 25721
rect 49148 25687 49200 25696
rect 49148 25653 49157 25687
rect 49157 25653 49191 25687
rect 49191 25653 49200 25687
rect 49148 25644 49200 25653
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 32950 25542 33002 25594
rect 33014 25542 33066 25594
rect 33078 25542 33130 25594
rect 33142 25542 33194 25594
rect 33206 25542 33258 25594
rect 42950 25542 43002 25594
rect 43014 25542 43066 25594
rect 43078 25542 43130 25594
rect 43142 25542 43194 25594
rect 43206 25542 43258 25594
rect 4988 25483 5040 25492
rect 4988 25449 4997 25483
rect 4997 25449 5031 25483
rect 5031 25449 5040 25483
rect 4988 25440 5040 25449
rect 1308 25304 1360 25356
rect 10968 25440 11020 25492
rect 25228 25440 25280 25492
rect 30012 25440 30064 25492
rect 37556 25440 37608 25492
rect 10876 25372 10928 25424
rect 27252 25372 27304 25424
rect 11060 25304 11112 25356
rect 24216 25304 24268 25356
rect 25136 25347 25188 25356
rect 25136 25313 25145 25347
rect 25145 25313 25179 25347
rect 25179 25313 25188 25347
rect 25136 25304 25188 25313
rect 25780 25304 25832 25356
rect 4160 25236 4212 25288
rect 6000 25236 6052 25288
rect 10600 25279 10652 25288
rect 10600 25245 10609 25279
rect 10609 25245 10643 25279
rect 10643 25245 10652 25279
rect 10600 25236 10652 25245
rect 16488 25236 16540 25288
rect 25964 25279 26016 25288
rect 25964 25245 25973 25279
rect 25973 25245 26007 25279
rect 26007 25245 26016 25279
rect 25964 25236 26016 25245
rect 30012 25304 30064 25356
rect 31760 25304 31812 25356
rect 32588 25347 32640 25356
rect 32588 25313 32597 25347
rect 32597 25313 32631 25347
rect 32631 25313 32640 25347
rect 32588 25304 32640 25313
rect 33968 25347 34020 25356
rect 33968 25313 33977 25347
rect 33977 25313 34011 25347
rect 34011 25313 34020 25347
rect 33968 25304 34020 25313
rect 34060 25347 34112 25356
rect 34060 25313 34069 25347
rect 34069 25313 34103 25347
rect 34103 25313 34112 25347
rect 34060 25304 34112 25313
rect 29000 25236 29052 25288
rect 29092 25236 29144 25288
rect 31944 25236 31996 25288
rect 34612 25236 34664 25288
rect 25504 25168 25556 25220
rect 25688 25168 25740 25220
rect 22284 25143 22336 25152
rect 22284 25109 22293 25143
rect 22293 25109 22327 25143
rect 22327 25109 22336 25143
rect 22284 25100 22336 25109
rect 22652 25143 22704 25152
rect 22652 25109 22661 25143
rect 22661 25109 22695 25143
rect 22695 25109 22704 25143
rect 22652 25100 22704 25109
rect 23296 25100 23348 25152
rect 26148 25100 26200 25152
rect 26332 25168 26384 25220
rect 29184 25168 29236 25220
rect 36176 25372 36228 25424
rect 39488 25483 39540 25492
rect 39488 25449 39497 25483
rect 39497 25449 39531 25483
rect 39531 25449 39540 25483
rect 39488 25440 39540 25449
rect 39672 25440 39724 25492
rect 49148 25440 49200 25492
rect 35624 25304 35676 25356
rect 36820 25304 36872 25356
rect 37372 25304 37424 25356
rect 37464 25304 37516 25356
rect 40684 25347 40736 25356
rect 40684 25313 40693 25347
rect 40693 25313 40727 25347
rect 40727 25313 40736 25347
rect 40684 25304 40736 25313
rect 34980 25236 35032 25288
rect 35072 25168 35124 25220
rect 27620 25100 27672 25152
rect 30656 25100 30708 25152
rect 31116 25100 31168 25152
rect 31392 25100 31444 25152
rect 32772 25100 32824 25152
rect 34152 25100 34204 25152
rect 36544 25143 36596 25152
rect 36544 25109 36553 25143
rect 36553 25109 36587 25143
rect 36587 25109 36596 25143
rect 36544 25100 36596 25109
rect 36912 25211 36964 25220
rect 36912 25177 36921 25211
rect 36921 25177 36955 25211
rect 36955 25177 36964 25211
rect 36912 25168 36964 25177
rect 37372 25168 37424 25220
rect 38292 25168 38344 25220
rect 39580 25168 39632 25220
rect 45284 25279 45336 25288
rect 45284 25245 45293 25279
rect 45293 25245 45327 25279
rect 45327 25245 45336 25279
rect 45284 25236 45336 25245
rect 46020 25279 46072 25288
rect 46020 25245 46029 25279
rect 46029 25245 46063 25279
rect 46063 25245 46072 25279
rect 46020 25236 46072 25245
rect 44640 25211 44692 25220
rect 44640 25177 44649 25211
rect 44649 25177 44683 25211
rect 44683 25177 44692 25211
rect 44640 25168 44692 25177
rect 45468 25211 45520 25220
rect 45468 25177 45477 25211
rect 45477 25177 45511 25211
rect 45511 25177 45520 25211
rect 45468 25168 45520 25177
rect 47860 25168 47912 25220
rect 38752 25100 38804 25152
rect 40040 25143 40092 25152
rect 40040 25109 40049 25143
rect 40049 25109 40083 25143
rect 40083 25109 40092 25143
rect 40040 25100 40092 25109
rect 40408 25143 40460 25152
rect 40408 25109 40417 25143
rect 40417 25109 40451 25143
rect 40451 25109 40460 25143
rect 40408 25100 40460 25109
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 27950 24998 28002 25050
rect 28014 24998 28066 25050
rect 28078 24998 28130 25050
rect 28142 24998 28194 25050
rect 28206 24998 28258 25050
rect 37950 24998 38002 25050
rect 38014 24998 38066 25050
rect 38078 24998 38130 25050
rect 38142 24998 38194 25050
rect 38206 24998 38258 25050
rect 47950 24998 48002 25050
rect 48014 24998 48066 25050
rect 48078 24998 48130 25050
rect 48142 24998 48194 25050
rect 48206 24998 48258 25050
rect 9404 24896 9456 24948
rect 27436 24896 27488 24948
rect 21364 24828 21416 24880
rect 23664 24828 23716 24880
rect 25872 24871 25924 24880
rect 25872 24837 25881 24871
rect 25881 24837 25915 24871
rect 25915 24837 25924 24871
rect 25872 24828 25924 24837
rect 25964 24828 26016 24880
rect 26148 24828 26200 24880
rect 26976 24828 27028 24880
rect 28448 24896 28500 24948
rect 9312 24760 9364 24812
rect 22652 24760 22704 24812
rect 27896 24828 27948 24880
rect 30288 24896 30340 24948
rect 29920 24828 29972 24880
rect 31024 24896 31076 24948
rect 36544 24896 36596 24948
rect 31668 24828 31720 24880
rect 34888 24828 34940 24880
rect 36176 24828 36228 24880
rect 36728 24828 36780 24880
rect 32864 24760 32916 24812
rect 8300 24692 8352 24744
rect 19708 24735 19760 24744
rect 19708 24701 19717 24735
rect 19717 24701 19751 24735
rect 19751 24701 19760 24735
rect 19708 24692 19760 24701
rect 21272 24692 21324 24744
rect 25596 24692 25648 24744
rect 25964 24735 26016 24744
rect 25964 24701 25973 24735
rect 25973 24701 26007 24735
rect 26007 24701 26016 24735
rect 25964 24692 26016 24701
rect 26240 24692 26292 24744
rect 21088 24624 21140 24676
rect 25136 24624 25188 24676
rect 29184 24692 29236 24744
rect 31300 24692 31352 24744
rect 32680 24692 32732 24744
rect 33692 24760 33744 24812
rect 36636 24760 36688 24812
rect 37280 24760 37332 24812
rect 40408 24760 40460 24812
rect 47216 24760 47268 24812
rect 33876 24692 33928 24744
rect 32312 24624 32364 24676
rect 34244 24735 34296 24744
rect 34244 24701 34253 24735
rect 34253 24701 34287 24735
rect 34287 24701 34296 24735
rect 34244 24692 34296 24701
rect 34704 24692 34756 24744
rect 39488 24692 39540 24744
rect 49148 24735 49200 24744
rect 49148 24701 49157 24735
rect 49157 24701 49191 24735
rect 49191 24701 49200 24735
rect 49148 24692 49200 24701
rect 21548 24556 21600 24608
rect 27528 24556 27580 24608
rect 27620 24556 27672 24608
rect 30288 24556 30340 24608
rect 31208 24556 31260 24608
rect 32220 24556 32272 24608
rect 32404 24556 32456 24608
rect 34980 24556 35032 24608
rect 35440 24556 35492 24608
rect 43812 24556 43864 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 14096 24352 14148 24404
rect 21824 24352 21876 24404
rect 19708 24216 19760 24268
rect 21456 24216 21508 24268
rect 25504 24259 25556 24268
rect 25504 24225 25513 24259
rect 25513 24225 25547 24259
rect 25547 24225 25556 24259
rect 25504 24216 25556 24225
rect 26792 24352 26844 24404
rect 34428 24352 34480 24404
rect 34612 24352 34664 24404
rect 27436 24284 27488 24336
rect 10600 24148 10652 24200
rect 12624 24148 12676 24200
rect 22836 24148 22888 24200
rect 27528 24216 27580 24268
rect 28080 24259 28132 24268
rect 28080 24225 28089 24259
rect 28089 24225 28123 24259
rect 28123 24225 28132 24259
rect 28080 24216 28132 24225
rect 31208 24284 31260 24336
rect 30196 24259 30248 24268
rect 30196 24225 30205 24259
rect 30205 24225 30239 24259
rect 30239 24225 30248 24259
rect 30196 24216 30248 24225
rect 30288 24259 30340 24268
rect 30288 24225 30297 24259
rect 30297 24225 30331 24259
rect 30331 24225 30340 24259
rect 30288 24216 30340 24225
rect 32864 24216 32916 24268
rect 34980 24259 35032 24268
rect 34980 24225 34989 24259
rect 34989 24225 35023 24259
rect 35023 24225 35032 24259
rect 34980 24216 35032 24225
rect 35716 24216 35768 24268
rect 39488 24284 39540 24336
rect 37740 24259 37792 24268
rect 37740 24225 37749 24259
rect 37749 24225 37783 24259
rect 37783 24225 37792 24259
rect 37740 24216 37792 24225
rect 40224 24216 40276 24268
rect 40776 24216 40828 24268
rect 21088 24123 21140 24132
rect 21088 24089 21097 24123
rect 21097 24089 21131 24123
rect 21131 24089 21140 24123
rect 21088 24080 21140 24089
rect 23664 24080 23716 24132
rect 11152 24055 11204 24064
rect 11152 24021 11161 24055
rect 11161 24021 11195 24055
rect 11195 24021 11204 24055
rect 11152 24012 11204 24021
rect 21272 24012 21324 24064
rect 22560 24055 22612 24064
rect 22560 24021 22569 24055
rect 22569 24021 22603 24055
rect 22603 24021 22612 24055
rect 22560 24012 22612 24021
rect 23848 24012 23900 24064
rect 26148 24012 26200 24064
rect 30472 24148 30524 24200
rect 32680 24148 32732 24200
rect 33416 24148 33468 24200
rect 34428 24148 34480 24200
rect 37832 24148 37884 24200
rect 40040 24148 40092 24200
rect 47768 24148 47820 24200
rect 29092 24080 29144 24132
rect 26608 24055 26660 24064
rect 26608 24021 26617 24055
rect 26617 24021 26651 24055
rect 26651 24021 26660 24055
rect 26608 24012 26660 24021
rect 27620 24055 27672 24064
rect 27620 24021 27629 24055
rect 27629 24021 27663 24055
rect 27663 24021 27672 24055
rect 27620 24012 27672 24021
rect 28080 24012 28132 24064
rect 28448 24012 28500 24064
rect 34704 24080 34756 24132
rect 30196 24012 30248 24064
rect 33416 24012 33468 24064
rect 33876 24012 33928 24064
rect 34428 24012 34480 24064
rect 34520 24012 34572 24064
rect 35716 24080 35768 24132
rect 37372 24080 37424 24132
rect 38476 24080 38528 24132
rect 49148 24123 49200 24132
rect 49148 24089 49157 24123
rect 49157 24089 49191 24123
rect 49191 24089 49200 24123
rect 49148 24080 49200 24089
rect 35164 24012 35216 24064
rect 35624 24012 35676 24064
rect 37464 24012 37516 24064
rect 37648 24012 37700 24064
rect 37832 24012 37884 24064
rect 40040 24055 40092 24064
rect 40040 24021 40049 24055
rect 40049 24021 40083 24055
rect 40083 24021 40092 24055
rect 40040 24012 40092 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 6000 23808 6052 23860
rect 11060 23808 11112 23860
rect 16488 23808 16540 23860
rect 23296 23808 23348 23860
rect 26792 23808 26844 23860
rect 30472 23808 30524 23860
rect 34060 23851 34112 23860
rect 34060 23817 34069 23851
rect 34069 23817 34103 23851
rect 34103 23817 34112 23851
rect 34060 23808 34112 23817
rect 34428 23808 34480 23860
rect 37096 23808 37148 23860
rect 39396 23808 39448 23860
rect 15292 23740 15344 23792
rect 20996 23740 21048 23792
rect 21824 23740 21876 23792
rect 23664 23740 23716 23792
rect 12164 23672 12216 23724
rect 7840 23604 7892 23656
rect 11152 23604 11204 23656
rect 21456 23672 21508 23724
rect 26608 23740 26660 23792
rect 27620 23740 27672 23792
rect 30564 23740 30616 23792
rect 14096 23579 14148 23588
rect 14096 23545 14105 23579
rect 14105 23545 14139 23579
rect 14139 23545 14148 23579
rect 14096 23536 14148 23545
rect 16488 23604 16540 23656
rect 16212 23468 16264 23520
rect 20904 23604 20956 23656
rect 21272 23647 21324 23656
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 21548 23536 21600 23588
rect 22100 23468 22152 23520
rect 22468 23468 22520 23520
rect 26148 23672 26200 23724
rect 31576 23672 31628 23724
rect 32496 23740 32548 23792
rect 33876 23740 33928 23792
rect 37740 23740 37792 23792
rect 39580 23740 39632 23792
rect 32312 23715 32364 23724
rect 32312 23681 32321 23715
rect 32321 23681 32355 23715
rect 32355 23681 32364 23715
rect 32312 23672 32364 23681
rect 33692 23672 33744 23724
rect 34520 23672 34572 23724
rect 23664 23536 23716 23588
rect 26424 23647 26476 23656
rect 26424 23613 26433 23647
rect 26433 23613 26467 23647
rect 26467 23613 26476 23647
rect 26424 23604 26476 23613
rect 26516 23604 26568 23656
rect 24676 23536 24728 23588
rect 32680 23604 32732 23656
rect 38568 23672 38620 23724
rect 46756 23672 46808 23724
rect 35164 23647 35216 23656
rect 35164 23613 35173 23647
rect 35173 23613 35207 23647
rect 35207 23613 35216 23647
rect 35164 23604 35216 23613
rect 49148 23647 49200 23656
rect 49148 23613 49157 23647
rect 49157 23613 49191 23647
rect 49191 23613 49200 23647
rect 49148 23604 49200 23613
rect 24952 23468 25004 23520
rect 25872 23511 25924 23520
rect 25872 23477 25881 23511
rect 25881 23477 25915 23511
rect 25915 23477 25924 23511
rect 25872 23468 25924 23477
rect 26148 23468 26200 23520
rect 34336 23468 34388 23520
rect 34520 23511 34572 23520
rect 34520 23477 34529 23511
rect 34529 23477 34563 23511
rect 34563 23477 34572 23511
rect 34520 23468 34572 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 4160 23264 4212 23316
rect 26976 23264 27028 23316
rect 27528 23264 27580 23316
rect 27620 23264 27672 23316
rect 31852 23307 31904 23316
rect 31852 23273 31861 23307
rect 31861 23273 31895 23307
rect 31895 23273 31904 23307
rect 31852 23264 31904 23273
rect 32588 23264 32640 23316
rect 34244 23264 34296 23316
rect 34336 23196 34388 23248
rect 44088 23196 44140 23248
rect 1308 23128 1360 23180
rect 5540 23128 5592 23180
rect 9036 23128 9088 23180
rect 16212 23128 16264 23180
rect 19708 23128 19760 23180
rect 21364 23128 21416 23180
rect 23664 23171 23716 23180
rect 23664 23137 23673 23171
rect 23673 23137 23707 23171
rect 23707 23137 23716 23171
rect 23664 23128 23716 23137
rect 25228 23171 25280 23180
rect 25228 23137 25237 23171
rect 25237 23137 25271 23171
rect 25271 23137 25280 23171
rect 25228 23128 25280 23137
rect 27160 23171 27212 23180
rect 27160 23137 27169 23171
rect 27169 23137 27203 23171
rect 27203 23137 27212 23171
rect 27160 23128 27212 23137
rect 29828 23128 29880 23180
rect 4896 23060 4948 23112
rect 9772 23060 9824 23112
rect 20812 23060 20864 23112
rect 24860 23060 24912 23112
rect 24952 23103 25004 23112
rect 24952 23069 24961 23103
rect 24961 23069 24995 23103
rect 24995 23069 25004 23103
rect 24952 23060 25004 23069
rect 28540 23060 28592 23112
rect 28816 23060 28868 23112
rect 37556 23128 37608 23180
rect 38752 23128 38804 23180
rect 39396 23128 39448 23180
rect 9680 22992 9732 23044
rect 15292 22992 15344 23044
rect 16212 22992 16264 23044
rect 17408 23035 17460 23044
rect 17408 23001 17417 23035
rect 17417 23001 17451 23035
rect 17451 23001 17460 23035
rect 17408 22992 17460 23001
rect 2780 22924 2832 22976
rect 18880 22967 18932 22976
rect 18880 22933 18889 22967
rect 18889 22933 18923 22967
rect 18923 22933 18932 22967
rect 18880 22924 18932 22933
rect 19708 23035 19760 23044
rect 19708 23001 19717 23035
rect 19717 23001 19751 23035
rect 19751 23001 19760 23035
rect 19708 22992 19760 23001
rect 22192 22992 22244 23044
rect 22744 22992 22796 23044
rect 24768 22992 24820 23044
rect 21180 22967 21232 22976
rect 21180 22933 21189 22967
rect 21189 22933 21223 22967
rect 21223 22933 21232 22967
rect 21180 22924 21232 22933
rect 22652 22924 22704 22976
rect 24952 22924 25004 22976
rect 25044 22967 25096 22976
rect 25044 22933 25053 22967
rect 25053 22933 25087 22967
rect 25087 22933 25096 22967
rect 25044 22924 25096 22933
rect 27528 22992 27580 23044
rect 29276 22924 29328 22976
rect 31668 22992 31720 23044
rect 33692 23060 33744 23112
rect 31760 22924 31812 22976
rect 32496 22992 32548 23044
rect 32588 23035 32640 23044
rect 32588 23001 32597 23035
rect 32597 23001 32631 23035
rect 32631 23001 32640 23035
rect 32588 22992 32640 23001
rect 33600 22924 33652 22976
rect 35164 23035 35216 23044
rect 35164 23001 35173 23035
rect 35173 23001 35207 23035
rect 35207 23001 35216 23035
rect 35164 22992 35216 23001
rect 35900 22992 35952 23044
rect 35532 22924 35584 22976
rect 47676 23060 47728 23112
rect 37464 22992 37516 23044
rect 49148 23035 49200 23044
rect 49148 23001 49157 23035
rect 49157 23001 49191 23035
rect 49191 23001 49200 23035
rect 49148 22992 49200 23001
rect 38292 22924 38344 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 22284 22720 22336 22772
rect 23664 22720 23716 22772
rect 24952 22720 25004 22772
rect 30380 22720 30432 22772
rect 32680 22720 32732 22772
rect 34520 22720 34572 22772
rect 37556 22720 37608 22772
rect 38568 22720 38620 22772
rect 17408 22652 17460 22704
rect 16488 22584 16540 22636
rect 18880 22584 18932 22636
rect 19892 22559 19944 22568
rect 19892 22525 19901 22559
rect 19901 22525 19935 22559
rect 19935 22525 19944 22559
rect 19892 22516 19944 22525
rect 23388 22652 23440 22704
rect 26884 22652 26936 22704
rect 28816 22652 28868 22704
rect 30472 22652 30524 22704
rect 23296 22584 23348 22636
rect 24768 22584 24820 22636
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 28540 22584 28592 22636
rect 21180 22516 21232 22568
rect 21364 22448 21416 22500
rect 25504 22516 25556 22568
rect 27528 22516 27580 22568
rect 30380 22584 30432 22636
rect 34152 22695 34204 22704
rect 34152 22661 34161 22695
rect 34161 22661 34195 22695
rect 34195 22661 34204 22695
rect 34152 22652 34204 22661
rect 37372 22584 37424 22636
rect 39580 22652 39632 22704
rect 42800 22652 42852 22704
rect 32864 22516 32916 22568
rect 34244 22559 34296 22568
rect 34244 22525 34253 22559
rect 34253 22525 34287 22559
rect 34287 22525 34296 22559
rect 34244 22516 34296 22525
rect 37832 22559 37884 22568
rect 37832 22525 37841 22559
rect 37841 22525 37875 22559
rect 37875 22525 37884 22559
rect 37832 22516 37884 22525
rect 39028 22516 39080 22568
rect 39488 22516 39540 22568
rect 26516 22448 26568 22500
rect 36912 22448 36964 22500
rect 46756 22448 46808 22500
rect 13360 22380 13412 22432
rect 16580 22380 16632 22432
rect 17408 22423 17460 22432
rect 17408 22389 17417 22423
rect 17417 22389 17451 22423
rect 17451 22389 17460 22423
rect 17408 22380 17460 22389
rect 21180 22380 21232 22432
rect 25044 22380 25096 22432
rect 25228 22380 25280 22432
rect 31300 22380 31352 22432
rect 32312 22380 32364 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 13360 22176 13412 22228
rect 5540 22151 5592 22160
rect 5540 22117 5549 22151
rect 5549 22117 5583 22151
rect 5583 22117 5592 22151
rect 5540 22108 5592 22117
rect 14096 22108 14148 22160
rect 23296 22219 23348 22228
rect 23296 22185 23305 22219
rect 23305 22185 23339 22219
rect 23339 22185 23348 22219
rect 23296 22176 23348 22185
rect 16488 22108 16540 22160
rect 21088 22108 21140 22160
rect 22560 22108 22612 22160
rect 9128 21972 9180 22024
rect 10232 21904 10284 21956
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 14832 22015 14884 22024
rect 14832 21981 14841 22015
rect 14841 21981 14875 22015
rect 14875 21981 14884 22015
rect 14832 21972 14884 21981
rect 16212 21972 16264 22024
rect 25044 22176 25096 22228
rect 26608 22176 26660 22228
rect 24216 22040 24268 22092
rect 25228 22108 25280 22160
rect 25596 22108 25648 22160
rect 31760 22176 31812 22228
rect 32680 22176 32732 22228
rect 34244 22176 34296 22228
rect 25780 22040 25832 22092
rect 26884 22108 26936 22160
rect 27804 22040 27856 22092
rect 30380 22108 30432 22160
rect 31668 22108 31720 22160
rect 33508 22108 33560 22160
rect 34428 22108 34480 22160
rect 9312 21836 9364 21888
rect 13544 21879 13596 21888
rect 13544 21845 13553 21879
rect 13553 21845 13587 21879
rect 13587 21845 13596 21879
rect 13544 21836 13596 21845
rect 16488 21904 16540 21956
rect 17408 21904 17460 21956
rect 20720 21904 20772 21956
rect 20996 21904 21048 21956
rect 22284 21904 22336 21956
rect 23572 21904 23624 21956
rect 23848 21904 23900 21956
rect 28448 21972 28500 22024
rect 29920 22015 29972 22024
rect 29920 21981 29929 22015
rect 29929 21981 29963 22015
rect 29963 21981 29972 22015
rect 29920 21972 29972 21981
rect 31116 22040 31168 22092
rect 26792 21904 26844 21956
rect 32864 21972 32916 22024
rect 37464 22040 37516 22092
rect 47584 21972 47636 22024
rect 49148 22015 49200 22024
rect 49148 21981 49157 22015
rect 49157 21981 49191 22015
rect 49191 21981 49200 22015
rect 49148 21972 49200 21981
rect 16580 21879 16632 21888
rect 16580 21845 16589 21879
rect 16589 21845 16623 21879
rect 16623 21845 16632 21879
rect 16580 21836 16632 21845
rect 20904 21879 20956 21888
rect 20904 21845 20913 21879
rect 20913 21845 20947 21879
rect 20947 21845 20956 21879
rect 20904 21836 20956 21845
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 24952 21836 25004 21888
rect 25596 21879 25648 21888
rect 25596 21845 25605 21879
rect 25605 21845 25639 21879
rect 25639 21845 25648 21879
rect 25596 21836 25648 21845
rect 26424 21836 26476 21888
rect 28724 21836 28776 21888
rect 35256 21904 35308 21956
rect 36084 21904 36136 21956
rect 32128 21836 32180 21888
rect 44180 21836 44232 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 10232 21675 10284 21684
rect 10232 21641 10241 21675
rect 10241 21641 10275 21675
rect 10275 21641 10284 21675
rect 10232 21632 10284 21641
rect 12164 21632 12216 21684
rect 23572 21632 23624 21684
rect 25872 21632 25924 21684
rect 29920 21632 29972 21684
rect 30472 21632 30524 21684
rect 13544 21496 13596 21548
rect 9772 21471 9824 21480
rect 9772 21437 9781 21471
rect 9781 21437 9815 21471
rect 9815 21437 9824 21471
rect 9772 21428 9824 21437
rect 14832 21496 14884 21548
rect 19616 21564 19668 21616
rect 20812 21564 20864 21616
rect 23480 21564 23532 21616
rect 25596 21564 25648 21616
rect 25136 21496 25188 21548
rect 16028 21428 16080 21480
rect 19524 21292 19576 21344
rect 22468 21471 22520 21480
rect 22468 21437 22477 21471
rect 22477 21437 22511 21471
rect 22511 21437 22520 21471
rect 22468 21428 22520 21437
rect 22836 21428 22888 21480
rect 25596 21471 25648 21480
rect 25596 21437 25605 21471
rect 25605 21437 25639 21471
rect 25639 21437 25648 21471
rect 25596 21428 25648 21437
rect 28632 21496 28684 21548
rect 30196 21564 30248 21616
rect 31760 21632 31812 21684
rect 32588 21632 32640 21684
rect 33508 21564 33560 21616
rect 25780 21428 25832 21480
rect 31668 21496 31720 21548
rect 32496 21539 32548 21548
rect 32496 21505 32505 21539
rect 32505 21505 32539 21539
rect 32539 21505 32548 21539
rect 32496 21496 32548 21505
rect 35256 21539 35308 21548
rect 35256 21505 35265 21539
rect 35265 21505 35299 21539
rect 35299 21505 35308 21539
rect 35256 21496 35308 21505
rect 38752 21607 38804 21616
rect 38752 21573 38761 21607
rect 38761 21573 38795 21607
rect 38795 21573 38804 21607
rect 38752 21564 38804 21573
rect 38844 21564 38896 21616
rect 39028 21564 39080 21616
rect 38476 21539 38528 21548
rect 38476 21505 38485 21539
rect 38485 21505 38519 21539
rect 38519 21505 38528 21539
rect 38476 21496 38528 21505
rect 46296 21496 46348 21548
rect 29828 21471 29880 21480
rect 29828 21437 29837 21471
rect 29837 21437 29871 21471
rect 29871 21437 29880 21471
rect 29828 21428 29880 21437
rect 31852 21428 31904 21480
rect 32220 21428 32272 21480
rect 34060 21428 34112 21480
rect 37832 21428 37884 21480
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 23940 21292 23992 21344
rect 24216 21335 24268 21344
rect 24216 21301 24225 21335
rect 24225 21301 24259 21335
rect 24259 21301 24268 21335
rect 24216 21292 24268 21301
rect 24768 21292 24820 21344
rect 27804 21292 27856 21344
rect 30656 21292 30708 21344
rect 32128 21292 32180 21344
rect 36820 21360 36872 21412
rect 34244 21335 34296 21344
rect 34244 21301 34253 21335
rect 34253 21301 34287 21335
rect 34287 21301 34296 21335
rect 34244 21292 34296 21301
rect 35072 21335 35124 21344
rect 35072 21301 35081 21335
rect 35081 21301 35115 21335
rect 35115 21301 35124 21335
rect 35072 21292 35124 21301
rect 43352 21292 43404 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 9680 21131 9732 21140
rect 9680 21097 9689 21131
rect 9689 21097 9723 21131
rect 9723 21097 9732 21131
rect 9680 21088 9732 21097
rect 19892 21088 19944 21140
rect 32496 21088 32548 21140
rect 32864 21088 32916 21140
rect 35072 21088 35124 21140
rect 42800 21088 42852 21140
rect 43720 21020 43772 21072
rect 10968 20952 11020 21004
rect 19708 20952 19760 21004
rect 24216 20952 24268 21004
rect 31760 20952 31812 21004
rect 7840 20884 7892 20936
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 19340 20884 19392 20936
rect 19524 20884 19576 20936
rect 30656 20927 30708 20936
rect 30656 20893 30665 20927
rect 30665 20893 30699 20927
rect 30699 20893 30708 20927
rect 30656 20884 30708 20893
rect 30748 20884 30800 20936
rect 34796 20952 34848 21004
rect 37832 20952 37884 21004
rect 34704 20884 34756 20936
rect 38292 20884 38344 20936
rect 43812 20927 43864 20936
rect 43812 20893 43821 20927
rect 43821 20893 43855 20927
rect 43855 20893 43864 20927
rect 43812 20884 43864 20893
rect 47032 20884 47084 20936
rect 45192 20816 45244 20868
rect 49148 20859 49200 20868
rect 49148 20825 49157 20859
rect 49157 20825 49191 20859
rect 49191 20825 49200 20859
rect 49148 20816 49200 20825
rect 2872 20748 2924 20800
rect 19892 20791 19944 20800
rect 19892 20757 19901 20791
rect 19901 20757 19935 20791
rect 19935 20757 19944 20791
rect 19892 20748 19944 20757
rect 30288 20791 30340 20800
rect 30288 20757 30297 20791
rect 30297 20757 30331 20791
rect 30331 20757 30340 20791
rect 30288 20748 30340 20757
rect 31392 20748 31444 20800
rect 32128 20791 32180 20800
rect 32128 20757 32137 20791
rect 32137 20757 32171 20791
rect 32171 20757 32180 20791
rect 32128 20748 32180 20757
rect 36452 20748 36504 20800
rect 38384 20748 38436 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 21180 20587 21232 20596
rect 21180 20553 21189 20587
rect 21189 20553 21223 20587
rect 21223 20553 21232 20587
rect 21180 20544 21232 20553
rect 25136 20544 25188 20596
rect 26148 20544 26200 20596
rect 23296 20476 23348 20528
rect 23480 20476 23532 20528
rect 2780 20408 2832 20460
rect 20812 20408 20864 20460
rect 22376 20408 22428 20460
rect 22468 20408 22520 20460
rect 26148 20451 26200 20460
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 30472 20587 30524 20596
rect 30472 20553 30481 20587
rect 30481 20553 30515 20587
rect 30515 20553 30524 20587
rect 30472 20544 30524 20553
rect 32864 20587 32916 20596
rect 32864 20553 32873 20587
rect 32873 20553 32907 20587
rect 32907 20553 32916 20587
rect 32864 20544 32916 20553
rect 30748 20476 30800 20528
rect 36912 20451 36964 20460
rect 36912 20417 36921 20451
rect 36921 20417 36955 20451
rect 36955 20417 36964 20451
rect 36912 20408 36964 20417
rect 47860 20408 47912 20460
rect 1308 20340 1360 20392
rect 21916 20340 21968 20392
rect 25504 20340 25556 20392
rect 26608 20340 26660 20392
rect 32220 20340 32272 20392
rect 34244 20340 34296 20392
rect 49148 20383 49200 20392
rect 49148 20349 49157 20383
rect 49157 20349 49191 20383
rect 49191 20349 49200 20383
rect 49148 20340 49200 20349
rect 18604 20272 18656 20324
rect 21180 20204 21232 20256
rect 27160 20272 27212 20324
rect 34980 20272 35032 20324
rect 37188 20272 37240 20324
rect 24584 20204 24636 20256
rect 24860 20204 24912 20256
rect 32588 20204 32640 20256
rect 44456 20204 44508 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 10968 20000 11020 20052
rect 19984 20000 20036 20052
rect 20536 20000 20588 20052
rect 24952 20000 25004 20052
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 31760 20000 31812 20052
rect 25504 19932 25556 19984
rect 27068 19932 27120 19984
rect 44916 19932 44968 19984
rect 18604 19907 18656 19916
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 19432 19864 19484 19916
rect 19616 19907 19668 19916
rect 19616 19873 19625 19907
rect 19625 19873 19659 19907
rect 19659 19873 19668 19907
rect 19616 19864 19668 19873
rect 22468 19864 22520 19916
rect 25136 19864 25188 19916
rect 15660 19796 15712 19848
rect 17316 19796 17368 19848
rect 17684 19796 17736 19848
rect 23940 19796 23992 19848
rect 27160 19839 27212 19848
rect 27160 19805 27169 19839
rect 27169 19805 27203 19839
rect 27203 19805 27212 19839
rect 27160 19796 27212 19805
rect 27528 19864 27580 19916
rect 32680 19864 32732 19916
rect 35348 19864 35400 19916
rect 27804 19796 27856 19848
rect 31944 19796 31996 19848
rect 32220 19796 32272 19848
rect 32312 19839 32364 19848
rect 32312 19805 32321 19839
rect 32321 19805 32355 19839
rect 32355 19805 32364 19839
rect 32312 19796 32364 19805
rect 33324 19796 33376 19848
rect 33968 19796 34020 19848
rect 35440 19796 35492 19848
rect 36360 19796 36412 19848
rect 44088 19796 44140 19848
rect 19800 19728 19852 19780
rect 20904 19728 20956 19780
rect 23480 19728 23532 19780
rect 24216 19728 24268 19780
rect 27344 19728 27396 19780
rect 34336 19728 34388 19780
rect 46204 19728 46256 19780
rect 21272 19660 21324 19712
rect 21456 19660 21508 19712
rect 23572 19703 23624 19712
rect 23572 19669 23581 19703
rect 23581 19669 23615 19703
rect 23615 19669 23624 19703
rect 23572 19660 23624 19669
rect 26516 19660 26568 19712
rect 27252 19703 27304 19712
rect 27252 19669 27261 19703
rect 27261 19669 27295 19703
rect 27295 19669 27304 19703
rect 27252 19660 27304 19669
rect 31944 19660 31996 19712
rect 33324 19660 33376 19712
rect 34980 19660 35032 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 16028 19456 16080 19508
rect 21364 19456 21416 19508
rect 20076 19388 20128 19440
rect 21732 19388 21784 19440
rect 22468 19388 22520 19440
rect 23296 19388 23348 19440
rect 20996 19320 21048 19372
rect 21456 19320 21508 19372
rect 22284 19320 22336 19372
rect 21272 19295 21324 19304
rect 21272 19261 21281 19295
rect 21281 19261 21315 19295
rect 21315 19261 21324 19295
rect 21272 19252 21324 19261
rect 21548 19252 21600 19304
rect 23296 19252 23348 19304
rect 23664 19388 23716 19440
rect 24124 19388 24176 19440
rect 24216 19388 24268 19440
rect 28356 19388 28408 19440
rect 23940 19320 23992 19372
rect 24400 19320 24452 19372
rect 26608 19363 26660 19372
rect 26608 19329 26617 19363
rect 26617 19329 26651 19363
rect 26651 19329 26660 19363
rect 26608 19320 26660 19329
rect 26792 19320 26844 19372
rect 28448 19320 28500 19372
rect 29736 19320 29788 19372
rect 36084 19388 36136 19440
rect 35348 19320 35400 19372
rect 23572 19116 23624 19168
rect 24584 19184 24636 19236
rect 27896 19252 27948 19304
rect 28816 19252 28868 19304
rect 29828 19252 29880 19304
rect 37280 19320 37332 19372
rect 38476 19456 38528 19508
rect 38568 19456 38620 19508
rect 38752 19388 38804 19440
rect 45468 19320 45520 19372
rect 49148 19363 49200 19372
rect 49148 19329 49157 19363
rect 49157 19329 49191 19363
rect 49191 19329 49200 19363
rect 49148 19320 49200 19329
rect 36636 19184 36688 19236
rect 37464 19184 37516 19236
rect 26332 19116 26384 19168
rect 27436 19116 27488 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 9772 18844 9824 18896
rect 19892 18912 19944 18964
rect 20996 18912 21048 18964
rect 23388 18912 23440 18964
rect 26148 18912 26200 18964
rect 24676 18844 24728 18896
rect 22376 18776 22428 18828
rect 22836 18776 22888 18828
rect 23572 18776 23624 18828
rect 24768 18776 24820 18828
rect 25596 18776 25648 18828
rect 9312 18708 9364 18760
rect 12624 18708 12676 18760
rect 21732 18751 21784 18760
rect 21732 18717 21741 18751
rect 21741 18717 21775 18751
rect 21775 18717 21784 18751
rect 21732 18708 21784 18717
rect 24860 18708 24912 18760
rect 22468 18640 22520 18692
rect 22560 18683 22612 18692
rect 22560 18649 22569 18683
rect 22569 18649 22603 18683
rect 22603 18649 22612 18683
rect 22560 18640 22612 18649
rect 26240 18708 26292 18760
rect 26424 18819 26476 18828
rect 26424 18785 26433 18819
rect 26433 18785 26467 18819
rect 26467 18785 26476 18819
rect 26424 18776 26476 18785
rect 26608 18819 26660 18828
rect 26608 18785 26617 18819
rect 26617 18785 26651 18819
rect 26651 18785 26660 18819
rect 26608 18776 26660 18785
rect 27896 18776 27948 18828
rect 28632 18776 28684 18828
rect 28724 18776 28776 18828
rect 28908 18819 28960 18828
rect 28908 18785 28917 18819
rect 28917 18785 28951 18819
rect 28951 18785 28960 18819
rect 28908 18776 28960 18785
rect 27160 18640 27212 18692
rect 2780 18572 2832 18624
rect 21364 18572 21416 18624
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 25964 18615 26016 18624
rect 25964 18581 25973 18615
rect 25973 18581 26007 18615
rect 26007 18581 26016 18615
rect 25964 18572 26016 18581
rect 26332 18615 26384 18624
rect 26332 18581 26341 18615
rect 26341 18581 26375 18615
rect 26375 18581 26384 18615
rect 26332 18572 26384 18581
rect 27252 18572 27304 18624
rect 34980 18912 35032 18964
rect 32864 18844 32916 18896
rect 31484 18819 31536 18828
rect 31484 18785 31493 18819
rect 31493 18785 31527 18819
rect 31527 18785 31536 18819
rect 31484 18776 31536 18785
rect 32496 18776 32548 18828
rect 37280 18776 37332 18828
rect 31300 18708 31352 18760
rect 34244 18708 34296 18760
rect 36084 18708 36136 18760
rect 36176 18708 36228 18760
rect 44180 18751 44232 18760
rect 44180 18717 44189 18751
rect 44189 18717 44223 18751
rect 44223 18717 44232 18751
rect 44180 18708 44232 18717
rect 44640 18708 44692 18760
rect 36728 18640 36780 18692
rect 34152 18572 34204 18624
rect 35164 18572 35216 18624
rect 38752 18640 38804 18692
rect 47860 18640 47912 18692
rect 49148 18683 49200 18692
rect 49148 18649 49157 18683
rect 49157 18649 49191 18683
rect 49191 18649 49200 18683
rect 49148 18640 49200 18649
rect 37372 18572 37424 18624
rect 37464 18572 37516 18624
rect 39212 18572 39264 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 21180 18411 21232 18420
rect 21180 18377 21189 18411
rect 21189 18377 21223 18411
rect 21223 18377 21232 18411
rect 21180 18368 21232 18377
rect 21272 18300 21324 18352
rect 21456 18300 21508 18352
rect 23572 18300 23624 18352
rect 24308 18368 24360 18420
rect 24952 18368 25004 18420
rect 28448 18368 28500 18420
rect 33600 18368 33652 18420
rect 34796 18368 34848 18420
rect 35072 18368 35124 18420
rect 38660 18368 38712 18420
rect 25044 18343 25096 18352
rect 25044 18309 25053 18343
rect 25053 18309 25087 18343
rect 25087 18309 25096 18343
rect 25044 18300 25096 18309
rect 27252 18300 27304 18352
rect 30840 18300 30892 18352
rect 32496 18300 32548 18352
rect 33876 18300 33928 18352
rect 34244 18300 34296 18352
rect 36084 18300 36136 18352
rect 36544 18300 36596 18352
rect 2872 18232 2924 18284
rect 22836 18232 22888 18284
rect 27620 18232 27672 18284
rect 1308 18164 1360 18216
rect 20996 18164 21048 18216
rect 20904 18096 20956 18148
rect 22560 18164 22612 18216
rect 27528 18164 27580 18216
rect 31944 18232 31996 18284
rect 46756 18232 46808 18284
rect 30380 18207 30432 18216
rect 30380 18173 30389 18207
rect 30389 18173 30423 18207
rect 30423 18173 30432 18207
rect 30380 18164 30432 18173
rect 30196 18096 30248 18148
rect 15660 18028 15712 18080
rect 22468 18028 22520 18080
rect 27896 18028 27948 18080
rect 34796 18207 34848 18216
rect 34796 18173 34805 18207
rect 34805 18173 34839 18207
rect 34839 18173 34848 18207
rect 34796 18164 34848 18173
rect 35348 18164 35400 18216
rect 38016 18164 38068 18216
rect 38568 18164 38620 18216
rect 49148 18207 49200 18216
rect 49148 18173 49157 18207
rect 49157 18173 49191 18207
rect 49191 18173 49200 18207
rect 49148 18164 49200 18173
rect 34888 18028 34940 18080
rect 35900 18028 35952 18080
rect 39764 18028 39816 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 20076 17824 20128 17876
rect 27344 17867 27396 17876
rect 27344 17833 27353 17867
rect 27353 17833 27387 17867
rect 27387 17833 27396 17867
rect 27344 17824 27396 17833
rect 32496 17824 32548 17876
rect 27436 17756 27488 17808
rect 20536 17731 20588 17740
rect 20536 17697 20545 17731
rect 20545 17697 20579 17731
rect 20579 17697 20588 17731
rect 20536 17688 20588 17697
rect 20996 17688 21048 17740
rect 21456 17688 21508 17740
rect 22376 17688 22428 17740
rect 27528 17688 27580 17740
rect 28908 17756 28960 17808
rect 29736 17688 29788 17740
rect 30196 17688 30248 17740
rect 31024 17688 31076 17740
rect 32220 17688 32272 17740
rect 37372 17824 37424 17876
rect 38200 17824 38252 17876
rect 33784 17731 33836 17740
rect 33784 17697 33793 17731
rect 33793 17697 33827 17731
rect 33827 17697 33836 17731
rect 33784 17688 33836 17697
rect 19248 17620 19300 17672
rect 23204 17620 23256 17672
rect 27620 17620 27672 17672
rect 28448 17620 28500 17672
rect 28632 17620 28684 17672
rect 23296 17552 23348 17604
rect 23572 17552 23624 17604
rect 30288 17552 30340 17604
rect 30932 17595 30984 17604
rect 30932 17561 30941 17595
rect 30941 17561 30975 17595
rect 30975 17561 30984 17595
rect 30932 17552 30984 17561
rect 19984 17484 20036 17536
rect 22744 17484 22796 17536
rect 29368 17484 29420 17536
rect 30564 17484 30616 17536
rect 33876 17620 33928 17672
rect 35808 17688 35860 17740
rect 37280 17688 37332 17740
rect 38016 17731 38068 17740
rect 38016 17697 38025 17731
rect 38025 17697 38059 17731
rect 38059 17697 38068 17731
rect 38016 17688 38068 17697
rect 42800 17620 42852 17672
rect 43352 17620 43404 17672
rect 33692 17527 33744 17536
rect 33692 17493 33701 17527
rect 33701 17493 33735 17527
rect 33735 17493 33744 17527
rect 33692 17484 33744 17493
rect 35900 17552 35952 17604
rect 36544 17552 36596 17604
rect 37096 17552 37148 17604
rect 37740 17484 37792 17536
rect 38660 17552 38712 17604
rect 44456 17595 44508 17604
rect 44456 17561 44465 17595
rect 44465 17561 44499 17595
rect 44499 17561 44508 17595
rect 44456 17552 44508 17561
rect 44548 17484 44600 17536
rect 45192 17620 45244 17672
rect 46848 17552 46900 17604
rect 49148 17595 49200 17604
rect 49148 17561 49157 17595
rect 49157 17561 49191 17595
rect 49191 17561 49200 17595
rect 49148 17552 49200 17561
rect 46664 17484 46716 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 20904 17280 20956 17332
rect 21456 17323 21508 17332
rect 21456 17289 21465 17323
rect 21465 17289 21499 17323
rect 21499 17289 21508 17323
rect 21456 17280 21508 17289
rect 22836 17323 22888 17332
rect 22836 17289 22845 17323
rect 22845 17289 22879 17323
rect 22879 17289 22888 17323
rect 22836 17280 22888 17289
rect 23204 17323 23256 17332
rect 23204 17289 23213 17323
rect 23213 17289 23247 17323
rect 23247 17289 23256 17323
rect 23204 17280 23256 17289
rect 25964 17280 26016 17332
rect 26332 17280 26384 17332
rect 31024 17280 31076 17332
rect 31116 17280 31168 17332
rect 34428 17280 34480 17332
rect 36544 17280 36596 17332
rect 38660 17280 38712 17332
rect 23388 17212 23440 17264
rect 21088 17144 21140 17196
rect 23204 17144 23256 17196
rect 24032 17144 24084 17196
rect 24308 17144 24360 17196
rect 19248 17076 19300 17128
rect 21916 17076 21968 17128
rect 25044 17212 25096 17264
rect 25872 17144 25924 17196
rect 21272 17008 21324 17060
rect 26608 17008 26660 17060
rect 27712 17119 27764 17128
rect 27712 17085 27721 17119
rect 27721 17085 27755 17119
rect 27755 17085 27764 17119
rect 27712 17076 27764 17085
rect 30564 17212 30616 17264
rect 28724 17144 28776 17196
rect 28172 17076 28224 17128
rect 28356 17076 28408 17128
rect 29552 17144 29604 17196
rect 32404 17144 32456 17196
rect 29736 17076 29788 17128
rect 30288 17119 30340 17128
rect 30288 17085 30297 17119
rect 30297 17085 30331 17119
rect 30331 17085 30340 17119
rect 30288 17076 30340 17085
rect 30932 17076 30984 17128
rect 33508 17076 33560 17128
rect 37556 17212 37608 17264
rect 43720 17255 43772 17264
rect 43720 17221 43729 17255
rect 43729 17221 43763 17255
rect 43763 17221 43772 17255
rect 43720 17212 43772 17221
rect 28448 16983 28500 16992
rect 28448 16949 28457 16983
rect 28457 16949 28491 16983
rect 28491 16949 28500 16983
rect 28448 16940 28500 16949
rect 32128 16940 32180 16992
rect 32312 16983 32364 16992
rect 32312 16949 32321 16983
rect 32321 16949 32355 16983
rect 32355 16949 32364 16983
rect 32312 16940 32364 16949
rect 32864 16940 32916 16992
rect 35348 17119 35400 17128
rect 35348 17085 35357 17119
rect 35357 17085 35391 17119
rect 35391 17085 35400 17119
rect 35348 17076 35400 17085
rect 35532 17008 35584 17060
rect 39948 17008 40000 17060
rect 46756 17008 46808 17060
rect 38108 16983 38160 16992
rect 38108 16949 38117 16983
rect 38117 16949 38151 16983
rect 38151 16949 38160 16983
rect 38108 16940 38160 16949
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 18604 16600 18656 16652
rect 19248 16600 19300 16652
rect 22468 16736 22520 16788
rect 23388 16779 23440 16788
rect 23388 16745 23397 16779
rect 23397 16745 23431 16779
rect 23431 16745 23440 16779
rect 23388 16736 23440 16745
rect 26608 16736 26660 16788
rect 27436 16736 27488 16788
rect 31116 16736 31168 16788
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 21916 16600 21968 16609
rect 24400 16600 24452 16652
rect 24768 16643 24820 16652
rect 24768 16609 24777 16643
rect 24777 16609 24811 16643
rect 24811 16609 24820 16643
rect 24768 16600 24820 16609
rect 25044 16643 25096 16652
rect 25044 16609 25053 16643
rect 25053 16609 25087 16643
rect 25087 16609 25096 16643
rect 25044 16600 25096 16609
rect 26792 16600 26844 16652
rect 28172 16600 28224 16652
rect 28908 16600 28960 16652
rect 32036 16600 32088 16652
rect 37096 16736 37148 16788
rect 34888 16643 34940 16652
rect 34888 16609 34897 16643
rect 34897 16609 34931 16643
rect 34931 16609 34940 16643
rect 34888 16600 34940 16609
rect 35532 16600 35584 16652
rect 37372 16600 37424 16652
rect 28448 16532 28500 16584
rect 30656 16532 30708 16584
rect 38108 16532 38160 16584
rect 46204 16532 46256 16584
rect 9772 16464 9824 16516
rect 19800 16464 19852 16516
rect 5632 16439 5684 16448
rect 5632 16405 5641 16439
rect 5641 16405 5675 16439
rect 5675 16405 5684 16439
rect 5632 16396 5684 16405
rect 19248 16396 19300 16448
rect 23296 16464 23348 16516
rect 24768 16464 24820 16516
rect 28724 16464 28776 16516
rect 21088 16396 21140 16448
rect 21180 16439 21232 16448
rect 21180 16405 21189 16439
rect 21189 16405 21223 16439
rect 21223 16405 21232 16439
rect 21180 16396 21232 16405
rect 26332 16396 26384 16448
rect 28264 16396 28316 16448
rect 28448 16396 28500 16448
rect 28816 16396 28868 16448
rect 29736 16396 29788 16448
rect 35440 16464 35492 16516
rect 36544 16464 36596 16516
rect 37740 16464 37792 16516
rect 49148 16507 49200 16516
rect 49148 16473 49157 16507
rect 49157 16473 49191 16507
rect 49191 16473 49200 16507
rect 49148 16464 49200 16473
rect 36636 16439 36688 16448
rect 36636 16405 36645 16439
rect 36645 16405 36679 16439
rect 36679 16405 36688 16439
rect 36636 16396 36688 16405
rect 39488 16396 39540 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 19984 16192 20036 16244
rect 27160 16235 27212 16244
rect 27160 16201 27169 16235
rect 27169 16201 27203 16235
rect 27203 16201 27212 16235
rect 27160 16192 27212 16201
rect 27436 16192 27488 16244
rect 28356 16192 28408 16244
rect 16580 16124 16632 16176
rect 24676 16124 24728 16176
rect 26884 16124 26936 16176
rect 29368 16124 29420 16176
rect 30472 16124 30524 16176
rect 2780 16056 2832 16108
rect 1308 15988 1360 16040
rect 22468 15988 22520 16040
rect 36452 16056 36504 16108
rect 40040 16056 40092 16108
rect 47860 16056 47912 16108
rect 24768 15988 24820 16040
rect 26148 15988 26200 16040
rect 27528 15988 27580 16040
rect 27804 15988 27856 16040
rect 28816 16031 28868 16040
rect 28816 15997 28825 16031
rect 28825 15997 28859 16031
rect 28859 15997 28868 16031
rect 28816 15988 28868 15997
rect 29460 15988 29512 16040
rect 28264 15852 28316 15904
rect 29644 15852 29696 15904
rect 32496 15988 32548 16040
rect 37464 15988 37516 16040
rect 49148 16031 49200 16040
rect 49148 15997 49157 16031
rect 49157 15997 49191 16031
rect 49191 15997 49200 16031
rect 49148 15988 49200 15997
rect 35072 15920 35124 15972
rect 30564 15895 30616 15904
rect 30564 15861 30573 15895
rect 30573 15861 30607 15895
rect 30607 15861 30616 15895
rect 30564 15852 30616 15861
rect 32864 15852 32916 15904
rect 33416 15852 33468 15904
rect 36452 15852 36504 15904
rect 37648 15895 37700 15904
rect 37648 15861 37657 15895
rect 37657 15861 37691 15895
rect 37691 15861 37700 15895
rect 37648 15852 37700 15861
rect 38476 15852 38528 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 26516 15691 26568 15700
rect 26516 15657 26525 15691
rect 26525 15657 26559 15691
rect 26559 15657 26568 15691
rect 26516 15648 26568 15657
rect 28816 15648 28868 15700
rect 29460 15648 29512 15700
rect 30196 15648 30248 15700
rect 39120 15648 39172 15700
rect 21364 15580 21416 15632
rect 24124 15512 24176 15564
rect 27344 15512 27396 15564
rect 27988 15512 28040 15564
rect 29644 15580 29696 15632
rect 29736 15555 29788 15564
rect 29736 15521 29745 15555
rect 29745 15521 29779 15555
rect 29779 15521 29788 15555
rect 29736 15512 29788 15521
rect 30564 15512 30616 15564
rect 33508 15512 33560 15564
rect 35808 15555 35860 15564
rect 35808 15521 35817 15555
rect 35817 15521 35851 15555
rect 35851 15521 35860 15555
rect 35808 15512 35860 15521
rect 37096 15512 37148 15564
rect 25320 15376 25372 15428
rect 25412 15376 25464 15428
rect 26884 15419 26936 15428
rect 26884 15385 26893 15419
rect 26893 15385 26927 15419
rect 26927 15385 26936 15419
rect 26884 15376 26936 15385
rect 27436 15376 27488 15428
rect 28264 15376 28316 15428
rect 28816 15376 28868 15428
rect 29184 15376 29236 15428
rect 22652 15308 22704 15360
rect 27344 15308 27396 15360
rect 32588 15487 32640 15496
rect 32588 15453 32597 15487
rect 32597 15453 32631 15487
rect 32631 15453 32640 15487
rect 32588 15444 32640 15453
rect 33416 15487 33468 15496
rect 33416 15453 33425 15487
rect 33425 15453 33459 15487
rect 33459 15453 33468 15487
rect 33416 15444 33468 15453
rect 46848 15444 46900 15496
rect 30472 15376 30524 15428
rect 32404 15351 32456 15360
rect 32404 15317 32413 15351
rect 32413 15317 32447 15351
rect 32447 15317 32456 15351
rect 32404 15308 32456 15317
rect 33600 15376 33652 15428
rect 36544 15376 36596 15428
rect 49148 15419 49200 15428
rect 49148 15385 49157 15419
rect 49157 15385 49191 15419
rect 49191 15385 49200 15419
rect 49148 15376 49200 15385
rect 34428 15308 34480 15360
rect 37740 15308 37792 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 20076 15104 20128 15156
rect 26148 15104 26200 15156
rect 29000 15104 29052 15156
rect 29460 15147 29512 15156
rect 29460 15113 29469 15147
rect 29469 15113 29503 15147
rect 29503 15113 29512 15147
rect 29460 15104 29512 15113
rect 29644 15104 29696 15156
rect 37648 15104 37700 15156
rect 24768 15036 24820 15088
rect 30104 15036 30156 15088
rect 31576 15079 31628 15088
rect 31576 15045 31585 15079
rect 31585 15045 31619 15079
rect 31619 15045 31628 15079
rect 31576 15036 31628 15045
rect 37556 15036 37608 15088
rect 17040 14968 17092 15020
rect 22468 15011 22520 15020
rect 22468 14977 22477 15011
rect 22477 14977 22511 15011
rect 22511 14977 22520 15011
rect 22468 14968 22520 14977
rect 27620 14968 27672 15020
rect 29092 14968 29144 15020
rect 32220 14968 32272 15020
rect 39764 14968 39816 15020
rect 46756 14968 46808 15020
rect 21180 14943 21232 14952
rect 21180 14909 21189 14943
rect 21189 14909 21223 14943
rect 21223 14909 21232 14943
rect 21180 14900 21232 14909
rect 26608 14900 26660 14952
rect 27712 14943 27764 14952
rect 27712 14909 27721 14943
rect 27721 14909 27755 14943
rect 27755 14909 27764 14943
rect 27712 14900 27764 14909
rect 27988 14943 28040 14952
rect 27988 14909 27997 14943
rect 27997 14909 28031 14943
rect 28031 14909 28040 14943
rect 27988 14900 28040 14909
rect 25872 14875 25924 14884
rect 25872 14841 25881 14875
rect 25881 14841 25915 14875
rect 25915 14841 25924 14875
rect 25872 14832 25924 14841
rect 31024 14900 31076 14952
rect 32864 14943 32916 14952
rect 32864 14909 32873 14943
rect 32873 14909 32907 14943
rect 32907 14909 32916 14943
rect 32864 14900 32916 14909
rect 36636 14900 36688 14952
rect 49148 14943 49200 14952
rect 49148 14909 49157 14943
rect 49157 14909 49191 14943
rect 49191 14909 49200 14943
rect 49148 14900 49200 14909
rect 30288 14832 30340 14884
rect 33784 14832 33836 14884
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 30196 14764 30248 14816
rect 37372 14764 37424 14816
rect 41328 14764 41380 14816
rect 44180 14764 44232 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 20536 14560 20588 14612
rect 30564 14560 30616 14612
rect 32220 14603 32272 14612
rect 32220 14569 32229 14603
rect 32229 14569 32263 14603
rect 32263 14569 32272 14603
rect 32220 14560 32272 14569
rect 27988 14492 28040 14544
rect 24860 14424 24912 14476
rect 27712 14424 27764 14476
rect 26148 14331 26200 14340
rect 26148 14297 26157 14331
rect 26157 14297 26191 14331
rect 26191 14297 26200 14331
rect 26148 14288 26200 14297
rect 24768 14220 24820 14272
rect 29092 14288 29144 14340
rect 30288 14492 30340 14544
rect 34428 14492 34480 14544
rect 39764 14492 39816 14544
rect 32496 14424 32548 14476
rect 33968 14424 34020 14476
rect 35440 14424 35492 14476
rect 37740 14467 37792 14476
rect 37740 14433 37749 14467
rect 37749 14433 37783 14467
rect 37783 14433 37792 14467
rect 37740 14424 37792 14433
rect 30196 14399 30248 14408
rect 30196 14365 30205 14399
rect 30205 14365 30239 14399
rect 30239 14365 30248 14399
rect 30196 14356 30248 14365
rect 30288 14356 30340 14408
rect 34612 14356 34664 14408
rect 39948 14356 40000 14408
rect 28816 14220 28868 14272
rect 35164 14331 35216 14340
rect 35164 14297 35173 14331
rect 35173 14297 35207 14331
rect 35207 14297 35216 14331
rect 35164 14288 35216 14297
rect 36912 14220 36964 14272
rect 44088 14220 44140 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 29276 13948 29328 14000
rect 34796 14016 34848 14068
rect 35808 14016 35860 14068
rect 38568 14016 38620 14068
rect 42708 14016 42760 14068
rect 5632 13880 5684 13932
rect 30564 13923 30616 13932
rect 30564 13889 30573 13923
rect 30573 13889 30607 13923
rect 30607 13889 30616 13923
rect 30564 13880 30616 13889
rect 36820 13948 36872 14000
rect 40040 13948 40092 14000
rect 35256 13880 35308 13932
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 29736 13812 29788 13864
rect 35532 13812 35584 13864
rect 36912 13923 36964 13932
rect 36912 13889 36921 13923
rect 36921 13889 36955 13923
rect 36955 13889 36964 13923
rect 36912 13880 36964 13889
rect 37832 13880 37884 13932
rect 39120 13923 39172 13932
rect 39120 13889 39129 13923
rect 39129 13889 39163 13923
rect 39163 13889 39172 13923
rect 39120 13880 39172 13889
rect 39488 13880 39540 13932
rect 46664 13880 46716 13932
rect 38384 13812 38436 13864
rect 40684 13812 40736 13864
rect 44364 13812 44416 13864
rect 49148 13855 49200 13864
rect 49148 13821 49157 13855
rect 49157 13821 49191 13855
rect 49191 13821 49200 13855
rect 49148 13812 49200 13821
rect 35440 13676 35492 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 27620 13472 27672 13524
rect 33968 13472 34020 13524
rect 28908 13404 28960 13456
rect 30564 13336 30616 13388
rect 34796 13336 34848 13388
rect 37740 13336 37792 13388
rect 25228 13268 25280 13320
rect 28908 13268 28960 13320
rect 33692 13268 33744 13320
rect 34152 13311 34204 13320
rect 34152 13277 34161 13311
rect 34161 13277 34195 13311
rect 34195 13277 34204 13311
rect 34152 13268 34204 13277
rect 37188 13311 37240 13320
rect 37188 13277 37197 13311
rect 37197 13277 37231 13311
rect 37231 13277 37240 13311
rect 37188 13268 37240 13277
rect 37372 13268 37424 13320
rect 40684 13311 40736 13320
rect 40684 13277 40693 13311
rect 40693 13277 40727 13311
rect 40727 13277 40736 13311
rect 40684 13268 40736 13277
rect 44548 13268 44600 13320
rect 36544 13200 36596 13252
rect 49148 13243 49200 13252
rect 49148 13209 49157 13243
rect 49157 13209 49191 13243
rect 49191 13209 49200 13243
rect 49148 13200 49200 13209
rect 24584 13132 24636 13184
rect 31760 13132 31812 13184
rect 32312 13132 32364 13184
rect 34244 13175 34296 13184
rect 34244 13141 34253 13175
rect 34253 13141 34287 13175
rect 34287 13141 34296 13175
rect 34244 13132 34296 13141
rect 37280 13175 37332 13184
rect 37280 13141 37289 13175
rect 37289 13141 37323 13175
rect 37323 13141 37332 13175
rect 37280 13132 37332 13141
rect 39856 13132 39908 13184
rect 46756 13132 46808 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 28724 12928 28776 12980
rect 29276 12971 29328 12980
rect 29276 12937 29285 12971
rect 29285 12937 29319 12971
rect 29319 12937 29328 12971
rect 29276 12928 29328 12937
rect 30288 12928 30340 12980
rect 30472 12971 30524 12980
rect 30472 12937 30481 12971
rect 30481 12937 30515 12971
rect 30515 12937 30524 12971
rect 30472 12928 30524 12937
rect 30656 12928 30708 12980
rect 31944 12928 31996 12980
rect 32312 12928 32364 12980
rect 26700 12860 26752 12912
rect 27804 12860 27856 12912
rect 32404 12860 32456 12912
rect 34888 12928 34940 12980
rect 35440 12971 35492 12980
rect 35440 12937 35449 12971
rect 35449 12937 35483 12971
rect 35483 12937 35492 12971
rect 35440 12928 35492 12937
rect 36176 12928 36228 12980
rect 36544 12928 36596 12980
rect 46020 12928 46072 12980
rect 33968 12903 34020 12912
rect 33968 12869 33977 12903
rect 33977 12869 34011 12903
rect 34011 12869 34020 12903
rect 33968 12860 34020 12869
rect 27804 12724 27856 12776
rect 28632 12724 28684 12776
rect 29552 12724 29604 12776
rect 30564 12767 30616 12776
rect 30564 12733 30573 12767
rect 30573 12733 30607 12767
rect 30607 12733 30616 12767
rect 30564 12724 30616 12733
rect 27160 12656 27212 12708
rect 29000 12656 29052 12708
rect 25228 12588 25280 12640
rect 35256 12792 35308 12844
rect 36176 12792 36228 12844
rect 36268 12835 36320 12844
rect 36268 12801 36277 12835
rect 36277 12801 36311 12835
rect 36311 12801 36320 12835
rect 36268 12792 36320 12801
rect 34428 12724 34480 12776
rect 38568 12860 38620 12912
rect 46756 12792 46808 12844
rect 49148 12767 49200 12776
rect 49148 12733 49157 12767
rect 49157 12733 49191 12767
rect 49191 12733 49200 12767
rect 49148 12724 49200 12733
rect 36544 12656 36596 12708
rect 44732 12656 44784 12708
rect 39948 12588 40000 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 36268 12384 36320 12436
rect 39856 12248 39908 12300
rect 3424 12180 3476 12232
rect 9404 12180 9456 12232
rect 28908 12180 28960 12232
rect 38292 12180 38344 12232
rect 41328 12180 41380 12232
rect 44732 12180 44784 12232
rect 29184 12112 29236 12164
rect 41880 12112 41932 12164
rect 49148 12155 49200 12164
rect 49148 12121 49157 12155
rect 49157 12121 49191 12155
rect 49191 12121 49200 12155
rect 49148 12112 49200 12121
rect 43352 12044 43404 12096
rect 44272 12087 44324 12096
rect 44272 12053 44281 12087
rect 44281 12053 44315 12087
rect 44315 12053 44324 12087
rect 44272 12044 44324 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 44180 11772 44232 11824
rect 39764 11704 39816 11756
rect 42708 11704 42760 11756
rect 44088 11636 44140 11688
rect 46756 11636 46808 11688
rect 46664 11568 46716 11620
rect 44180 11500 44232 11552
rect 46296 11543 46348 11552
rect 46296 11509 46305 11543
rect 46305 11509 46339 11543
rect 46339 11509 46348 11543
rect 46296 11500 46348 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 17040 11296 17092 11348
rect 19800 11160 19852 11212
rect 44272 11092 44324 11144
rect 49148 11135 49200 11144
rect 49148 11101 49157 11135
rect 49157 11101 49191 11135
rect 49191 11101 49200 11135
rect 49148 11092 49200 11101
rect 7564 11024 7616 11076
rect 44364 11024 44416 11076
rect 46480 11067 46532 11076
rect 46480 11033 46489 11067
rect 46489 11033 46523 11067
rect 46523 11033 46532 11067
rect 46480 11024 46532 11033
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 24308 10684 24360 10736
rect 39948 10616 40000 10668
rect 47768 10616 47820 10668
rect 49148 10591 49200 10600
rect 49148 10557 49157 10591
rect 49157 10557 49191 10591
rect 49191 10557 49200 10591
rect 49148 10548 49200 10557
rect 25136 10480 25188 10532
rect 42708 10412 42760 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 28448 10004 28500 10056
rect 31852 10047 31904 10056
rect 31852 10013 31861 10047
rect 31861 10013 31895 10047
rect 31895 10013 31904 10047
rect 31852 10004 31904 10013
rect 46756 10004 46808 10056
rect 30104 9936 30156 9988
rect 49148 9979 49200 9988
rect 49148 9945 49157 9979
rect 49157 9945 49191 9979
rect 49191 9945 49200 9979
rect 49148 9936 49200 9945
rect 29920 9868 29972 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 32036 9596 32088 9648
rect 34980 9596 35032 9648
rect 44180 9528 44232 9580
rect 46664 9528 46716 9580
rect 49148 9503 49200 9512
rect 49148 9469 49157 9503
rect 49157 9469 49191 9503
rect 49191 9469 49200 9503
rect 49148 9460 49200 9469
rect 33968 9392 34020 9444
rect 37372 9392 37424 9444
rect 47860 9324 47912 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 3332 9052 3384 9104
rect 9588 9052 9640 9104
rect 43352 8916 43404 8968
rect 46204 8891 46256 8900
rect 46204 8857 46213 8891
rect 46213 8857 46247 8891
rect 46247 8857 46256 8891
rect 46204 8848 46256 8857
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 5540 8508 5592 8560
rect 16488 8508 16540 8560
rect 19248 8508 19300 8560
rect 32312 8508 32364 8560
rect 38476 8508 38528 8560
rect 42708 8508 42760 8560
rect 18604 8440 18656 8492
rect 46480 8440 46532 8492
rect 21548 8372 21600 8424
rect 42616 8372 42668 8424
rect 49148 8415 49200 8424
rect 49148 8381 49157 8415
rect 49157 8381 49191 8415
rect 49191 8381 49200 8415
rect 49148 8372 49200 8381
rect 16488 8304 16540 8356
rect 37648 8304 37700 8356
rect 45928 8347 45980 8356
rect 45928 8313 45937 8347
rect 45937 8313 45971 8347
rect 45971 8313 45980 8347
rect 45928 8304 45980 8313
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 46296 7828 46348 7880
rect 49148 7803 49200 7812
rect 49148 7769 49157 7803
rect 49157 7769 49191 7803
rect 49191 7769 49200 7803
rect 49148 7760 49200 7769
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 31760 7420 31812 7472
rect 29368 7352 29420 7404
rect 47860 7352 47912 7404
rect 49148 7327 49200 7336
rect 49148 7293 49157 7327
rect 49157 7293 49191 7327
rect 49191 7293 49200 7327
rect 49148 7284 49200 7293
rect 45192 7216 45244 7268
rect 41420 7148 41472 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 3424 6808 3476 6860
rect 8944 6808 8996 6860
rect 45928 6808 45980 6860
rect 36544 6740 36596 6792
rect 32404 6672 32456 6724
rect 40132 6740 40184 6792
rect 47400 6783 47452 6792
rect 47400 6749 47409 6783
rect 47409 6749 47443 6783
rect 47443 6749 47452 6783
rect 47400 6740 47452 6749
rect 44456 6672 44508 6724
rect 49148 6715 49200 6724
rect 49148 6681 49157 6715
rect 49157 6681 49191 6715
rect 49191 6681 49200 6715
rect 49148 6672 49200 6681
rect 47492 6604 47544 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 48780 6264 48832 6316
rect 48320 6060 48372 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 46204 5652 46256 5704
rect 49148 5695 49200 5704
rect 49148 5661 49157 5695
rect 49157 5661 49191 5695
rect 49191 5661 49200 5695
rect 49148 5652 49200 5661
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 10048 5176 10100 5228
rect 3424 4972 3476 5024
rect 9036 4972 9088 5024
rect 47860 4972 47912 5024
rect 49332 5015 49384 5024
rect 49332 4981 49341 5015
rect 49341 4981 49375 5015
rect 49375 4981 49384 5015
rect 49332 4972 49384 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 24676 4564 24728 4616
rect 49148 4539 49200 4548
rect 49148 4505 49157 4539
rect 49157 4505 49191 4539
rect 49191 4505 49200 4539
rect 49148 4496 49200 4505
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 33968 4131 34020 4140
rect 33968 4097 33977 4131
rect 33977 4097 34011 4131
rect 34011 4097 34020 4131
rect 33968 4088 34020 4097
rect 38384 4088 38436 4140
rect 40132 4088 40184 4140
rect 46020 4131 46072 4140
rect 46020 4097 46029 4131
rect 46029 4097 46063 4131
rect 46063 4097 46072 4131
rect 46020 4088 46072 4097
rect 48780 4131 48832 4140
rect 48780 4097 48789 4131
rect 48789 4097 48823 4131
rect 48823 4097 48832 4131
rect 48780 4088 48832 4097
rect 33876 4020 33928 4072
rect 39028 4020 39080 4072
rect 43444 4020 43496 4072
rect 48596 4020 48648 4072
rect 47768 3884 47820 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 5540 3680 5592 3732
rect 24308 3544 24360 3596
rect 29460 3544 29512 3596
rect 30932 3544 30984 3596
rect 34612 3544 34664 3596
rect 36084 3544 36136 3596
rect 39764 3544 39816 3596
rect 41236 3544 41288 3596
rect 44180 3544 44232 3596
rect 2780 3476 2832 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 29736 3519 29788 3528
rect 29736 3485 29745 3519
rect 29745 3485 29779 3519
rect 29779 3485 29788 3519
rect 29736 3476 29788 3485
rect 30104 3476 30156 3528
rect 34244 3476 34296 3528
rect 36728 3519 36780 3528
rect 36728 3485 36737 3519
rect 36737 3485 36771 3519
rect 36771 3485 36780 3519
rect 36728 3476 36780 3485
rect 37372 3476 37424 3528
rect 41880 3519 41932 3528
rect 41880 3485 41889 3519
rect 41889 3485 41923 3519
rect 41923 3485 41932 3519
rect 41880 3476 41932 3485
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 48320 3476 48372 3528
rect 6920 3408 6972 3460
rect 21364 3408 21416 3460
rect 49332 3408 49384 3460
rect 12808 3340 12860 3392
rect 27252 3340 27304 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 12808 3179 12860 3188
rect 12808 3145 12817 3179
rect 12817 3145 12851 3179
rect 12851 3145 12860 3179
rect 12808 3136 12860 3145
rect 17224 3136 17276 3188
rect 17960 3179 18012 3188
rect 17960 3145 17969 3179
rect 17969 3145 18003 3179
rect 18003 3145 18012 3179
rect 17960 3136 18012 3145
rect 19984 3068 20036 3120
rect 1492 3000 1544 3052
rect 756 2932 808 2984
rect 3700 3000 3752 3052
rect 5172 3000 5224 3052
rect 6644 3000 6696 3052
rect 10324 3000 10376 3052
rect 12532 3000 12584 3052
rect 14004 3000 14056 3052
rect 17684 3000 17736 3052
rect 28356 3136 28408 3188
rect 17316 2932 17368 2984
rect 19156 2932 19208 2984
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 22100 2932 22152 2984
rect 5448 2907 5500 2916
rect 5448 2873 5457 2907
rect 5457 2873 5491 2907
rect 5491 2873 5500 2907
rect 5448 2864 5500 2873
rect 7564 2864 7616 2916
rect 14464 2864 14516 2916
rect 27436 3068 27488 3120
rect 37280 3068 37332 3120
rect 24124 3000 24176 3052
rect 25136 3043 25188 3052
rect 25136 3009 25145 3043
rect 25145 3009 25179 3043
rect 25179 3009 25188 3043
rect 25136 3000 25188 3009
rect 27344 3043 27396 3052
rect 27344 3009 27353 3043
rect 27353 3009 27387 3043
rect 27387 3009 27396 3043
rect 27344 3000 27396 3009
rect 29184 3043 29236 3052
rect 29184 3009 29193 3043
rect 29193 3009 29227 3043
rect 29227 3009 29236 3043
rect 29184 3000 29236 3009
rect 33324 3000 33376 3052
rect 34336 3043 34388 3052
rect 34336 3009 34345 3043
rect 34345 3009 34379 3043
rect 34379 3009 34388 3043
rect 34336 3000 34388 3009
rect 37648 3043 37700 3052
rect 37648 3009 37657 3043
rect 37657 3009 37691 3043
rect 37691 3009 37700 3043
rect 37648 3000 37700 3009
rect 42616 3043 42668 3052
rect 42616 3009 42625 3043
rect 42625 3009 42659 3043
rect 42659 3009 42668 3043
rect 42616 3000 42668 3009
rect 44456 3043 44508 3052
rect 44456 3009 44465 3043
rect 44465 3009 44499 3043
rect 44499 3009 44508 3043
rect 44456 3000 44508 3009
rect 47400 3000 47452 3052
rect 47492 3000 47544 3052
rect 23572 2932 23624 2984
rect 25044 2932 25096 2984
rect 27252 2932 27304 2984
rect 28724 2932 28776 2984
rect 31668 2932 31720 2984
rect 30472 2864 30524 2916
rect 32404 2864 32456 2916
rect 36820 2932 36872 2984
rect 37556 2864 37608 2916
rect 41972 2932 42024 2984
rect 42708 2864 42760 2916
rect 47124 2932 47176 2984
rect 47860 2932 47912 2984
rect 46388 2796 46440 2848
rect 48320 2796 48372 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 14464 2592 14516 2644
rect 18696 2592 18748 2644
rect 16396 2456 16448 2508
rect 2228 2388 2280 2440
rect 7380 2388 7432 2440
rect 2964 2320 3016 2372
rect 4436 2320 4488 2372
rect 5908 2320 5960 2372
rect 6000 2363 6052 2372
rect 6000 2329 6009 2363
rect 6009 2329 6043 2363
rect 6043 2329 6052 2363
rect 6000 2320 6052 2329
rect 7840 2320 7892 2372
rect 8852 2320 8904 2372
rect 9588 2388 9640 2440
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 14740 2388 14792 2440
rect 16580 2524 16632 2576
rect 20720 2592 20772 2644
rect 20812 2592 20864 2644
rect 22192 2592 22244 2644
rect 46020 2592 46072 2644
rect 27804 2524 27856 2576
rect 18420 2456 18472 2508
rect 21364 2456 21416 2508
rect 22836 2456 22888 2508
rect 25780 2499 25832 2508
rect 25780 2465 25789 2499
rect 25789 2465 25823 2499
rect 25823 2465 25832 2499
rect 25780 2456 25832 2465
rect 26516 2456 26568 2508
rect 28356 2456 28408 2508
rect 30288 2456 30340 2508
rect 35348 2456 35400 2508
rect 38292 2456 38344 2508
rect 40592 2456 40644 2508
rect 48320 2499 48372 2508
rect 48320 2465 48329 2499
rect 48329 2465 48363 2499
rect 48363 2465 48372 2499
rect 48320 2456 48372 2465
rect 2412 2295 2464 2304
rect 2412 2261 2421 2295
rect 2421 2261 2455 2295
rect 2455 2261 2464 2295
rect 2412 2252 2464 2261
rect 3332 2295 3384 2304
rect 3332 2261 3341 2295
rect 3341 2261 3375 2295
rect 3375 2261 3384 2295
rect 3332 2252 3384 2261
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 11060 2320 11112 2372
rect 11152 2363 11204 2372
rect 11152 2329 11161 2363
rect 11161 2329 11195 2363
rect 11195 2329 11204 2363
rect 11152 2320 11204 2329
rect 11796 2320 11848 2372
rect 13268 2320 13320 2372
rect 15476 2320 15528 2372
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 16212 2320 16264 2372
rect 16304 2363 16356 2372
rect 16304 2329 16313 2363
rect 16313 2329 16347 2363
rect 16347 2329 16356 2363
rect 16304 2320 16356 2329
rect 16948 2320 17000 2372
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 19892 2388 19944 2440
rect 20904 2431 20956 2440
rect 20904 2397 20913 2431
rect 20913 2397 20947 2431
rect 20947 2397 20956 2431
rect 20904 2388 20956 2397
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 29920 2431 29972 2440
rect 29920 2397 29929 2431
rect 29929 2397 29963 2431
rect 29963 2397 29972 2431
rect 29920 2388 29972 2397
rect 31024 2388 31076 2440
rect 33784 2388 33836 2440
rect 35256 2388 35308 2440
rect 40040 2431 40092 2440
rect 40040 2397 40049 2431
rect 40049 2397 40083 2431
rect 40083 2397 40092 2431
rect 40040 2388 40092 2397
rect 41420 2388 41472 2440
rect 47768 2431 47820 2440
rect 47768 2397 47777 2431
rect 47777 2397 47811 2431
rect 47811 2397 47820 2431
rect 47768 2388 47820 2397
rect 23664 2320 23716 2372
rect 20812 2252 20864 2304
rect 20996 2252 21048 2304
rect 23756 2252 23808 2304
rect 33140 2252 33192 2304
rect 45652 2320 45704 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
rect 13636 2048 13688 2100
rect 22560 2048 22612 2100
rect 14464 1980 14516 2032
rect 20996 1980 21048 2032
rect 16304 1912 16356 1964
rect 28540 1912 28592 1964
rect 18328 1844 18380 1896
rect 28816 1844 28868 1896
rect 2412 1776 2464 1828
rect 19524 1776 19576 1828
rect 20904 1776 20956 1828
rect 29276 1776 29328 1828
rect 3332 1708 3384 1760
rect 21088 1708 21140 1760
rect 17500 1640 17552 1692
rect 26056 1640 26108 1692
<< metal2 >>
rect 386 56200 442 57000
rect 1122 56200 1178 57000
rect 1858 56200 1914 57000
rect 2594 56200 2650 57000
rect 3330 56200 3386 57000
rect 4066 56200 4122 57000
rect 4802 56200 4858 57000
rect 5538 56200 5594 57000
rect 6274 56200 6330 57000
rect 7010 56200 7066 57000
rect 7746 56200 7802 57000
rect 8482 56200 8538 57000
rect 9218 56200 9274 57000
rect 9954 56200 10010 57000
rect 10690 56200 10746 57000
rect 11426 56200 11482 57000
rect 12162 56200 12218 57000
rect 12898 56200 12954 57000
rect 13634 56200 13690 57000
rect 14370 56200 14426 57000
rect 15106 56200 15162 57000
rect 15842 56200 15898 57000
rect 16578 56200 16634 57000
rect 17314 56200 17370 57000
rect 18050 56200 18106 57000
rect 18156 56222 18368 56250
rect 400 55758 428 56200
rect 388 55752 440 55758
rect 388 55694 440 55700
rect 940 53100 992 53106
rect 940 53042 992 53048
rect 952 52737 980 53042
rect 938 52728 994 52737
rect 938 52663 994 52672
rect 1136 52562 1164 56200
rect 1872 53650 1900 56200
rect 1860 53644 1912 53650
rect 1860 53586 1912 53592
rect 2608 53038 2636 56200
rect 2872 55752 2924 55758
rect 2872 55694 2924 55700
rect 2778 55040 2834 55049
rect 2778 54975 2834 54984
rect 2792 54194 2820 54975
rect 2780 54188 2832 54194
rect 2780 54130 2832 54136
rect 2596 53032 2648 53038
rect 2596 52974 2648 52980
rect 1952 52964 2004 52970
rect 1952 52906 2004 52912
rect 1124 52556 1176 52562
rect 1124 52498 1176 52504
rect 1584 52012 1636 52018
rect 1584 51954 1636 51960
rect 940 50924 992 50930
rect 940 50866 992 50872
rect 952 50425 980 50866
rect 938 50416 994 50425
rect 938 50351 994 50360
rect 938 48104 994 48113
rect 938 48039 940 48048
rect 992 48039 994 48048
rect 940 48010 992 48016
rect 940 45892 992 45898
rect 940 45834 992 45840
rect 952 45801 980 45834
rect 938 45792 994 45801
rect 938 45727 994 45736
rect 1596 41818 1624 51954
rect 1676 50720 1728 50726
rect 1676 50662 1728 50668
rect 1688 42242 1716 50662
rect 1860 48068 1912 48074
rect 1860 48010 1912 48016
rect 1768 45824 1820 45830
rect 1768 45766 1820 45772
rect 1780 45626 1808 45766
rect 1768 45620 1820 45626
rect 1768 45562 1820 45568
rect 1688 42214 1808 42242
rect 1584 41812 1636 41818
rect 1584 41754 1636 41760
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 1688 41177 1716 41482
rect 1674 41168 1730 41177
rect 1674 41103 1730 41112
rect 1780 39114 1808 42214
rect 1872 39302 1900 48010
rect 1964 41206 1992 52906
rect 2884 52086 2912 55694
rect 3344 54262 3372 56200
rect 3332 54256 3384 54262
rect 3332 54198 3384 54204
rect 3976 53984 4028 53990
rect 3976 53926 4028 53932
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 2872 52080 2924 52086
rect 2872 52022 2924 52028
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 3988 48074 4016 53926
rect 4080 52562 4108 56200
rect 4816 55214 4844 56200
rect 4816 55186 4936 55214
rect 4908 53038 4936 55186
rect 5552 53650 5580 56200
rect 6288 54262 6316 56200
rect 6276 54256 6328 54262
rect 6276 54198 6328 54204
rect 7024 53650 7052 56200
rect 5540 53644 5592 53650
rect 5540 53586 5592 53592
rect 7012 53644 7064 53650
rect 7012 53586 7064 53592
rect 6276 53508 6328 53514
rect 6276 53450 6328 53456
rect 4896 53032 4948 53038
rect 4896 52974 4948 52980
rect 5816 52624 5868 52630
rect 5816 52566 5868 52572
rect 4068 52556 4120 52562
rect 4068 52498 4120 52504
rect 3976 48068 4028 48074
rect 3976 48010 4028 48016
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 5828 41274 5856 52566
rect 6288 42362 6316 53450
rect 6368 53168 6420 53174
rect 6368 53110 6420 53116
rect 6276 42356 6328 42362
rect 6276 42298 6328 42304
rect 6380 42294 6408 53110
rect 7760 53038 7788 56200
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8496 54262 8524 56200
rect 8484 54256 8536 54262
rect 8484 54198 8536 54204
rect 8944 53576 8996 53582
rect 8944 53518 8996 53524
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7748 53032 7800 53038
rect 7748 52974 7800 52980
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8956 43246 8984 53518
rect 9036 53100 9088 53106
rect 9036 53042 9088 53048
rect 9048 43926 9076 53042
rect 9232 52562 9260 56200
rect 9864 53168 9916 53174
rect 9864 53110 9916 53116
rect 9772 53100 9824 53106
rect 9772 53042 9824 53048
rect 9220 52556 9272 52562
rect 9220 52498 9272 52504
rect 9128 52488 9180 52494
rect 9128 52430 9180 52436
rect 9036 43920 9088 43926
rect 9036 43862 9088 43868
rect 8944 43240 8996 43246
rect 8944 43182 8996 43188
rect 9140 42770 9168 52430
rect 9784 44538 9812 53042
rect 9772 44532 9824 44538
rect 9772 44474 9824 44480
rect 9128 42764 9180 42770
rect 9128 42706 9180 42712
rect 9220 42628 9272 42634
rect 9220 42570 9272 42576
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 6368 42288 6420 42294
rect 6368 42230 6420 42236
rect 7104 42220 7156 42226
rect 7104 42162 7156 42168
rect 7840 42220 7892 42226
rect 7840 42162 7892 42168
rect 5816 41268 5868 41274
rect 5816 41210 5868 41216
rect 1952 41200 2004 41206
rect 1952 41142 2004 41148
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 1860 39296 1912 39302
rect 1860 39238 1912 39244
rect 1780 39086 1900 39114
rect 1872 38962 1900 39086
rect 940 38956 992 38962
rect 940 38898 992 38904
rect 1860 38956 1912 38962
rect 1860 38898 1912 38904
rect 952 38865 980 38898
rect 938 38856 994 38865
rect 938 38791 994 38800
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 940 36780 992 36786
rect 940 36722 992 36728
rect 952 36553 980 36722
rect 938 36544 994 36553
rect 938 36479 994 36488
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1780 34241 1808 34546
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 1766 34232 1822 34241
rect 2950 34235 3258 34244
rect 1766 34167 1822 34176
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 940 32428 992 32434
rect 940 32370 992 32376
rect 952 31929 980 32370
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 938 31920 994 31929
rect 938 31855 994 31864
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 1308 29708 1360 29714
rect 1308 29650 1360 29656
rect 1320 29617 1348 29650
rect 4804 29640 4856 29646
rect 1306 29608 1362 29617
rect 4804 29582 4856 29588
rect 1306 29543 1362 29552
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 4816 28218 4844 29582
rect 7116 28422 7144 42162
rect 7380 38752 7432 38758
rect 7380 38694 7432 38700
rect 7392 30258 7420 38694
rect 7564 36576 7616 36582
rect 7564 36518 7616 36524
rect 7472 32224 7524 32230
rect 7472 32166 7524 32172
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 4804 28212 4856 28218
rect 4804 28154 4856 28160
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 1308 27532 1360 27538
rect 1308 27474 1360 27480
rect 1320 27305 1348 27474
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 4896 27396 4948 27402
rect 4896 27338 4948 27344
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 1308 25356 1360 25362
rect 1308 25298 1360 25304
rect 1320 24993 1348 25298
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 1306 24984 1362 24993
rect 1306 24919 1362 24928
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 4172 23322 4200 25230
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 1308 23180 1360 23186
rect 1308 23122 1360 23128
rect 1320 22681 1348 23122
rect 4908 23118 4936 27338
rect 5000 25498 5028 27406
rect 7484 25906 7512 32166
rect 7576 28082 7604 36518
rect 7852 35894 7880 42162
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 7760 35866 7880 35894
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 7656 30184 7708 30190
rect 7656 30126 7708 30132
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7668 27606 7696 30126
rect 7760 29034 7788 35866
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 7840 34740 7892 34746
rect 7840 34682 7892 34688
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7748 28008 7800 28014
rect 7748 27950 7800 27956
rect 7656 27600 7708 27606
rect 7656 27542 7708 27548
rect 7760 26586 7788 27950
rect 7852 26994 7880 34682
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 9232 30598 9260 42570
rect 9876 41274 9904 53110
rect 9968 53038 9996 56200
rect 10048 54324 10100 54330
rect 10048 54266 10100 54272
rect 9956 53032 10008 53038
rect 9956 52974 10008 52980
rect 10060 51610 10088 54266
rect 10704 53650 10732 56200
rect 11440 54262 11468 56200
rect 11428 54256 11480 54262
rect 11428 54198 11480 54204
rect 11704 54188 11756 54194
rect 11704 54130 11756 54136
rect 10692 53644 10744 53650
rect 10692 53586 10744 53592
rect 10416 53576 10468 53582
rect 10416 53518 10468 53524
rect 10048 51604 10100 51610
rect 10048 51546 10100 51552
rect 10428 45558 10456 53518
rect 10784 53508 10836 53514
rect 10784 53450 10836 53456
rect 10416 45552 10468 45558
rect 10416 45494 10468 45500
rect 10600 41472 10652 41478
rect 10600 41414 10652 41420
rect 9864 41268 9916 41274
rect 9864 41210 9916 41216
rect 9772 41132 9824 41138
rect 9772 41074 9824 41080
rect 9784 31385 9812 41074
rect 9770 31376 9826 31385
rect 9770 31311 9826 31320
rect 9220 30592 9272 30598
rect 9220 30534 9272 30540
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 9128 30184 9180 30190
rect 9128 30126 9180 30132
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7748 26376 7800 26382
rect 7748 26318 7800 26324
rect 7760 26234 7788 26318
rect 7760 26206 7880 26234
rect 7472 25900 7524 25906
rect 7472 25842 7524 25848
rect 4988 25492 5040 25498
rect 4988 25434 5040 25440
rect 6000 25288 6052 25294
rect 6000 25230 6052 25236
rect 6012 23866 6040 25230
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 7852 23662 7880 26206
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 8312 24750 8340 26862
rect 9036 25832 9088 25838
rect 9036 25774 9088 25780
rect 8942 24984 8998 24993
rect 8942 24919 8998 24928
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 1306 22672 1362 22681
rect 1306 22607 1362 22616
rect 2792 20466 2820 22918
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 5552 22166 5580 23122
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 7852 20942 7880 23598
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 1308 20392 1360 20398
rect 1306 20360 1308 20369
rect 1360 20360 1362 20369
rect 1306 20295 1362 20304
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 1308 18216 1360 18222
rect 1308 18158 1360 18164
rect 1320 18057 1348 18158
rect 1306 18048 1362 18057
rect 1306 17983 1362 17992
rect 2792 16114 2820 18566
rect 2884 18290 2912 20742
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15745 1348 15982
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 1306 15736 1362 15745
rect 2950 15739 3258 15748
rect 1306 15671 1362 15680
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 5644 13938 5672 16390
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13433 2820 13806
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2778 13424 2834 13433
rect 2778 13359 2834 13368
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3436 11121 3464 12174
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 3422 11112 3478 11121
rect 3422 11047 3478 11056
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3344 8809 3372 9046
rect 3330 8800 3386 8809
rect 3330 8735 3386 8744
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3436 4185 3464 4966
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 5552 3738 5580 8502
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 756 2984 808 2990
rect 756 2926 808 2932
rect 768 800 796 2926
rect 1504 800 1532 2994
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2240 800 2268 2382
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2424 1834 2452 2246
rect 2792 1873 2820 3470
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6932 3194 6960 3402
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2778 1864 2834 1873
rect 2412 1828 2464 1834
rect 2778 1799 2834 1808
rect 2412 1770 2464 1776
rect 2976 800 3004 2314
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 1766 3372 2246
rect 3332 1760 3384 1766
rect 3332 1702 3384 1708
rect 3712 800 3740 2994
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4448 800 4476 2314
rect 5184 800 5212 2994
rect 5446 2952 5502 2961
rect 5446 2887 5448 2896
rect 5500 2887 5502 2896
rect 5448 2858 5500 2864
rect 5998 2408 6054 2417
rect 5908 2372 5960 2378
rect 5998 2343 6000 2352
rect 5908 2314 5960 2320
rect 6052 2343 6054 2352
rect 6000 2314 6052 2320
rect 5920 800 5948 2314
rect 6656 800 6684 2994
rect 7576 2922 7604 11018
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8956 6866 8984 24919
rect 9048 23186 9076 25774
rect 9036 23180 9088 23186
rect 9036 23122 9088 23128
rect 9140 22030 9168 30126
rect 9496 28008 9548 28014
rect 9496 27950 9548 27956
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9416 24954 9444 25774
rect 9508 25265 9536 27950
rect 9680 27940 9732 27946
rect 9680 27882 9732 27888
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9494 25256 9550 25265
rect 9494 25191 9550 25200
rect 9508 24993 9536 25191
rect 9494 24984 9550 24993
rect 9404 24948 9456 24954
rect 9494 24919 9550 24928
rect 9404 24890 9456 24896
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9140 6914 9168 21966
rect 9324 21894 9352 24754
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9324 20942 9352 21830
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9324 18766 9352 20878
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9416 12238 9444 24890
rect 9600 22681 9628 26862
rect 9692 26586 9720 27882
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9784 26382 9812 27406
rect 9772 26376 9824 26382
rect 9772 26318 9824 26324
rect 10612 25294 10640 41414
rect 10796 41274 10824 53450
rect 11716 43994 11744 54130
rect 12176 53650 12204 56200
rect 12912 55214 12940 56200
rect 12820 55186 12940 55214
rect 12348 53984 12400 53990
rect 12348 53926 12400 53932
rect 12164 53644 12216 53650
rect 12164 53586 12216 53592
rect 12360 49978 12388 53926
rect 12820 53038 12848 55186
rect 13648 54262 13676 56200
rect 13636 54256 13688 54262
rect 13636 54198 13688 54204
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12808 53032 12860 53038
rect 12808 52974 12860 52980
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 14384 52562 14412 56200
rect 14556 54188 14608 54194
rect 14556 54130 14608 54136
rect 14372 52556 14424 52562
rect 14372 52498 14424 52504
rect 14464 52488 14516 52494
rect 14464 52430 14516 52436
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 14476 51610 14504 52430
rect 14464 51604 14516 51610
rect 14464 51546 14516 51552
rect 14280 51332 14332 51338
rect 14280 51274 14332 51280
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12348 49972 12400 49978
rect 12348 49914 12400 49920
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 14292 45898 14320 51274
rect 14280 45892 14332 45898
rect 14280 45834 14332 45840
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 14464 44396 14516 44402
rect 14464 44338 14516 44344
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 11704 43988 11756 43994
rect 11704 43930 11756 43936
rect 12164 43716 12216 43722
rect 12164 43658 12216 43664
rect 13452 43716 13504 43722
rect 13452 43658 13504 43664
rect 12176 43382 12204 43658
rect 12164 43376 12216 43382
rect 12164 43318 12216 43324
rect 12072 43308 12124 43314
rect 12072 43250 12124 43256
rect 10784 41268 10836 41274
rect 10784 41210 10836 41216
rect 10692 41132 10744 41138
rect 10692 41074 10744 41080
rect 10704 29850 10732 41074
rect 12084 32774 12112 43250
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12072 32768 12124 32774
rect 12072 32710 12124 32716
rect 13464 32502 13492 43658
rect 14476 37194 14504 44338
rect 14568 42770 14596 54130
rect 14648 54052 14700 54058
rect 14648 53994 14700 54000
rect 14660 43994 14688 53994
rect 14740 53576 14792 53582
rect 14740 53518 14792 53524
rect 14752 49978 14780 53518
rect 15120 53038 15148 56200
rect 15856 53718 15884 56200
rect 16592 54262 16620 56200
rect 16580 54256 16632 54262
rect 16580 54198 16632 54204
rect 15844 53712 15896 53718
rect 15844 53654 15896 53660
rect 16948 53168 17000 53174
rect 16948 53110 17000 53116
rect 15200 53100 15252 53106
rect 15200 53042 15252 53048
rect 15108 53032 15160 53038
rect 15108 52974 15160 52980
rect 14740 49972 14792 49978
rect 14740 49914 14792 49920
rect 15212 49434 15240 53042
rect 15936 51332 15988 51338
rect 15936 51274 15988 51280
rect 15200 49428 15252 49434
rect 15200 49370 15252 49376
rect 15948 46170 15976 51274
rect 16856 49836 16908 49842
rect 16856 49778 16908 49784
rect 15936 46164 15988 46170
rect 15936 46106 15988 46112
rect 14648 43988 14700 43994
rect 14648 43930 14700 43936
rect 16120 43716 16172 43722
rect 16120 43658 16172 43664
rect 14556 42764 14608 42770
rect 14556 42706 14608 42712
rect 14464 37188 14516 37194
rect 14464 37130 14516 37136
rect 13452 32496 13504 32502
rect 13452 32438 13504 32444
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 10692 29844 10744 29850
rect 10692 29786 10744 29792
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 10876 26444 10928 26450
rect 10876 26386 10928 26392
rect 10888 25430 10916 26386
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10980 25498 11008 26318
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 10876 25424 10928 25430
rect 10876 25366 10928 25372
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10612 24206 10640 25230
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 11072 23866 11100 25298
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11164 23662 11192 24006
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9586 22672 9642 22681
rect 9586 22607 9642 22616
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9600 9110 9628 22607
rect 9692 21146 9720 22986
rect 9784 21486 9812 23054
rect 10232 21956 10284 21962
rect 10232 21898 10284 21904
rect 10244 21690 10272 21898
rect 12176 21690 12204 23666
rect 12636 22030 12664 24142
rect 14108 23594 14136 24346
rect 14096 23588 14148 23594
rect 14096 23530 14148 23536
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13372 22234 13400 22374
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 14108 22166 14136 23530
rect 14096 22160 14148 22166
rect 14096 22102 14148 22108
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9784 18902 9812 21422
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10980 20058 11008 20946
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9784 16522 9812 18838
rect 12636 18766 12664 21966
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13556 21554 13584 21830
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 9048 6886 9168 6914
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 9048 5030 9076 6886
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 7392 800 7420 2382
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 754 0 810 800
rect 1490 0 1546 800
rect 2226 0 2282 800
rect 2962 0 3018 800
rect 3698 0 3754 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7378 0 7434 800
rect 7852 762 7880 2314
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8864 800 8892 2314
rect 9600 800 9628 2382
rect 10060 2310 10088 5170
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 3194 12848 3334
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10336 800 10364 2994
rect 12346 2544 12402 2553
rect 12346 2479 12402 2488
rect 12360 2446 12388 2479
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 11072 800 11100 2314
rect 11164 1873 11192 2314
rect 11150 1864 11206 1873
rect 11150 1799 11206 1808
rect 11808 800 11836 2314
rect 12544 800 12572 2994
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 13280 800 13308 2314
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13648 2106 13676 2246
rect 13636 2100 13688 2106
rect 13636 2042 13688 2048
rect 14016 800 14044 2994
rect 14476 2922 14504 37130
rect 16132 35834 16160 43658
rect 16868 43450 16896 49778
rect 16960 43994 16988 53110
rect 17328 53038 17356 56200
rect 18064 56114 18092 56200
rect 18156 56114 18184 56222
rect 18064 56086 18184 56114
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 17684 54188 17736 54194
rect 17684 54130 17736 54136
rect 17316 53032 17368 53038
rect 17316 52974 17368 52980
rect 17696 50522 17724 54130
rect 18340 53650 18368 56222
rect 18786 56200 18842 57000
rect 19522 56200 19578 57000
rect 20258 56200 20314 57000
rect 20994 56200 21050 57000
rect 21730 56200 21786 57000
rect 22466 56200 22522 57000
rect 23202 56200 23258 57000
rect 23938 56200 23994 57000
rect 24674 56200 24730 57000
rect 25410 56200 25466 57000
rect 26146 56200 26202 57000
rect 26882 56200 26938 57000
rect 27618 56200 27674 57000
rect 28354 56200 28410 57000
rect 29090 56200 29146 57000
rect 29826 56200 29882 57000
rect 30562 56200 30618 57000
rect 31298 56200 31354 57000
rect 32034 56200 32090 57000
rect 32770 56200 32826 57000
rect 33506 56200 33562 57000
rect 34242 56200 34298 57000
rect 34978 56200 35034 57000
rect 35714 56200 35770 57000
rect 36450 56200 36506 57000
rect 37186 56200 37242 57000
rect 37922 56200 37978 57000
rect 38658 56200 38714 57000
rect 39394 56200 39450 57000
rect 40130 56200 40186 57000
rect 40866 56200 40922 57000
rect 41602 56200 41658 57000
rect 42338 56200 42394 57000
rect 43074 56200 43130 57000
rect 43810 56200 43866 57000
rect 43916 56222 44128 56250
rect 18800 54262 18828 56200
rect 18788 54256 18840 54262
rect 18788 54198 18840 54204
rect 18328 53644 18380 53650
rect 18328 53586 18380 53592
rect 18420 53576 18472 53582
rect 18420 53518 18472 53524
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17684 50516 17736 50522
rect 17684 50458 17736 50464
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 18432 49434 18460 53518
rect 19536 53038 19564 56200
rect 20168 54120 20220 54126
rect 20168 54062 20220 54068
rect 19616 53100 19668 53106
rect 19616 53042 19668 53048
rect 19524 53032 19576 53038
rect 19524 52974 19576 52980
rect 19156 52488 19208 52494
rect 19156 52430 19208 52436
rect 18420 49428 18472 49434
rect 18420 49370 18472 49376
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 16948 43988 17000 43994
rect 16948 43930 17000 43936
rect 17040 43716 17092 43722
rect 17040 43658 17092 43664
rect 16856 43444 16908 43450
rect 16856 43386 16908 43392
rect 16120 35828 16172 35834
rect 16120 35770 16172 35776
rect 17052 35193 17080 43658
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 19168 43450 19196 52430
rect 19628 43926 19656 53042
rect 20180 45554 20208 54062
rect 20272 53650 20300 56200
rect 21008 54262 21036 56200
rect 20996 54256 21048 54262
rect 20996 54198 21048 54204
rect 20352 54188 20404 54194
rect 20352 54130 20404 54136
rect 20260 53644 20312 53650
rect 20260 53586 20312 53592
rect 20364 50998 20392 54130
rect 21744 53650 21772 56200
rect 22480 54126 22508 56200
rect 23216 55214 23244 56200
rect 23216 55186 23336 55214
rect 22744 54188 22796 54194
rect 22744 54130 22796 54136
rect 22468 54120 22520 54126
rect 22468 54062 22520 54068
rect 21732 53644 21784 53650
rect 21732 53586 21784 53592
rect 22192 53508 22244 53514
rect 22192 53450 22244 53456
rect 20444 53440 20496 53446
rect 20444 53382 20496 53388
rect 20352 50992 20404 50998
rect 20352 50934 20404 50940
rect 20180 45526 20392 45554
rect 19616 43920 19668 43926
rect 19616 43862 19668 43868
rect 20364 43450 20392 45526
rect 20456 43994 20484 53382
rect 21272 53168 21324 53174
rect 21272 53110 21324 53116
rect 20904 49904 20956 49910
rect 20904 49846 20956 49852
rect 20720 49224 20772 49230
rect 20720 49166 20772 49172
rect 20536 48000 20588 48006
rect 20536 47942 20588 47948
rect 20444 43988 20496 43994
rect 20444 43930 20496 43936
rect 19156 43444 19208 43450
rect 19156 43386 19208 43392
rect 20352 43444 20404 43450
rect 20352 43386 20404 43392
rect 19064 43308 19116 43314
rect 19064 43250 19116 43256
rect 20260 43308 20312 43314
rect 20260 43250 20312 43256
rect 17408 42628 17460 42634
rect 17408 42570 17460 42576
rect 17224 36780 17276 36786
rect 17224 36722 17276 36728
rect 17038 35184 17094 35193
rect 17038 35119 17094 35128
rect 17236 32570 17264 36722
rect 17224 32564 17276 32570
rect 17224 32506 17276 32512
rect 17420 31754 17448 42570
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17684 41064 17736 41070
rect 17684 41006 17736 41012
rect 17696 32570 17724 41006
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 17684 32564 17736 32570
rect 17684 32506 17736 32512
rect 17236 31726 17448 31754
rect 17236 29238 17264 31726
rect 17224 29232 17276 29238
rect 17224 29174 17276 29180
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16500 23866 16528 25230
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 15292 23792 15344 23798
rect 15292 23734 15344 23740
rect 15304 23050 15332 23734
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16224 23186 16252 23462
rect 16212 23180 16264 23186
rect 16212 23122 16264 23128
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 16212 23044 16264 23050
rect 16212 22986 16264 22992
rect 16224 22030 16252 22986
rect 16500 22642 16528 23598
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 14844 21554 14872 21966
rect 16500 21962 16528 22102
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16592 21894 16620 22374
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15672 18086 15700 19790
rect 16040 19514 16068 21422
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 16592 16182 16620 21830
rect 16580 16176 16632 16182
rect 16580 16118 16632 16124
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17052 11354 17080 14962
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16500 8362 16528 8502
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 17236 3194 17264 29174
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17420 22710 17448 22986
rect 17408 22704 17460 22710
rect 17408 22646 17460 22652
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17420 21962 17448 22374
rect 17408 21956 17460 21962
rect 17408 21898 17460 21904
rect 17696 19854 17724 32506
rect 19076 31754 19104 43250
rect 19432 43240 19484 43246
rect 19432 43182 19484 43188
rect 19444 36922 19472 43182
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 20272 32230 20300 43250
rect 20548 42022 20576 47942
rect 20628 45892 20680 45898
rect 20628 45834 20680 45840
rect 20536 42016 20588 42022
rect 20536 41958 20588 41964
rect 20640 40662 20668 45834
rect 20732 42362 20760 49166
rect 20916 43450 20944 49846
rect 21088 48204 21140 48210
rect 21088 48146 21140 48152
rect 20904 43444 20956 43450
rect 20904 43386 20956 43392
rect 20720 42356 20772 42362
rect 20720 42298 20772 42304
rect 20996 42220 21048 42226
rect 20996 42162 21048 42168
rect 20628 40656 20680 40662
rect 20628 40598 20680 40604
rect 20720 38412 20772 38418
rect 20720 38354 20772 38360
rect 20732 37210 20760 38354
rect 20548 37182 20760 37210
rect 20548 36242 20576 37182
rect 20536 36236 20588 36242
rect 20536 36178 20588 36184
rect 20548 35494 20576 36178
rect 20536 35488 20588 35494
rect 20536 35430 20588 35436
rect 20548 35086 20576 35430
rect 20536 35080 20588 35086
rect 20536 35022 20588 35028
rect 21008 34202 21036 42162
rect 21100 38418 21128 48146
rect 21284 43994 21312 53110
rect 22204 51066 22232 53450
rect 22756 52154 22784 54130
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23308 53582 23336 55186
rect 23952 53582 23980 56200
rect 24688 54262 24716 56200
rect 24676 54256 24728 54262
rect 24676 54198 24728 54204
rect 25424 54194 25452 56200
rect 26160 54210 26188 56200
rect 26160 54194 26280 54210
rect 26896 54194 26924 56200
rect 27632 54194 27660 56200
rect 27950 54428 28258 54437
rect 27950 54426 27956 54428
rect 28012 54426 28036 54428
rect 28092 54426 28116 54428
rect 28172 54426 28196 54428
rect 28252 54426 28258 54428
rect 28012 54374 28014 54426
rect 28194 54374 28196 54426
rect 27950 54372 27956 54374
rect 28012 54372 28036 54374
rect 28092 54372 28116 54374
rect 28172 54372 28196 54374
rect 28252 54372 28258 54374
rect 27950 54363 28258 54372
rect 28368 54262 28396 56200
rect 28908 54324 28960 54330
rect 28908 54266 28960 54272
rect 28356 54256 28408 54262
rect 28356 54198 28408 54204
rect 25412 54188 25464 54194
rect 26160 54188 26292 54194
rect 26160 54182 26240 54188
rect 25412 54130 25464 54136
rect 26240 54130 26292 54136
rect 26884 54188 26936 54194
rect 26884 54130 26936 54136
rect 27620 54188 27672 54194
rect 27620 54130 27672 54136
rect 25228 54052 25280 54058
rect 25228 53994 25280 54000
rect 22836 53576 22888 53582
rect 22836 53518 22888 53524
rect 23296 53576 23348 53582
rect 23296 53518 23348 53524
rect 23940 53576 23992 53582
rect 23940 53518 23992 53524
rect 22744 52148 22796 52154
rect 22744 52090 22796 52096
rect 22848 51610 22876 53518
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 23756 52012 23808 52018
rect 23756 51954 23808 51960
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22836 51604 22888 51610
rect 22836 51546 22888 51552
rect 22192 51060 22244 51066
rect 22192 51002 22244 51008
rect 22744 50924 22796 50930
rect 22744 50866 22796 50872
rect 21824 50244 21876 50250
rect 21824 50186 21876 50192
rect 21548 45484 21600 45490
rect 21548 45426 21600 45432
rect 21272 43988 21324 43994
rect 21272 43930 21324 43936
rect 21180 43716 21232 43722
rect 21180 43658 21232 43664
rect 21088 38412 21140 38418
rect 21088 38354 21140 38360
rect 21192 35894 21220 43658
rect 21364 38276 21416 38282
rect 21364 38218 21416 38224
rect 21376 36718 21404 38218
rect 21560 37466 21588 45426
rect 21836 43994 21864 50186
rect 22100 49156 22152 49162
rect 22100 49098 22152 49104
rect 21916 48068 21968 48074
rect 21916 48010 21968 48016
rect 21824 43988 21876 43994
rect 21824 43930 21876 43936
rect 21928 43466 21956 48010
rect 22008 45960 22060 45966
rect 22008 45902 22060 45908
rect 21836 43438 21956 43466
rect 21836 41070 21864 43438
rect 21916 43376 21968 43382
rect 21916 43318 21968 43324
rect 21824 41064 21876 41070
rect 21824 41006 21876 41012
rect 21548 37460 21600 37466
rect 21548 37402 21600 37408
rect 21824 36848 21876 36854
rect 21824 36790 21876 36796
rect 21364 36712 21416 36718
rect 21364 36654 21416 36660
rect 21192 35866 21312 35894
rect 21180 35828 21232 35834
rect 21180 35770 21232 35776
rect 21192 35494 21220 35770
rect 21180 35488 21232 35494
rect 21180 35430 21232 35436
rect 20996 34196 21048 34202
rect 20996 34138 21048 34144
rect 21088 33448 21140 33454
rect 21284 33425 21312 35866
rect 21376 35834 21404 36654
rect 21836 36106 21864 36790
rect 21928 36310 21956 43318
rect 22020 40730 22048 45902
rect 22112 42362 22140 49098
rect 22468 45620 22520 45626
rect 22468 45562 22520 45568
rect 22284 43784 22336 43790
rect 22284 43726 22336 43732
rect 22100 42356 22152 42362
rect 22100 42298 22152 42304
rect 22296 41414 22324 43726
rect 22376 42016 22428 42022
rect 22376 41958 22428 41964
rect 22388 41546 22416 41958
rect 22376 41540 22428 41546
rect 22376 41482 22428 41488
rect 22480 41414 22508 45562
rect 22756 45082 22784 50866
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 23768 47802 23796 51954
rect 24124 50924 24176 50930
rect 24124 50866 24176 50872
rect 23756 47796 23808 47802
rect 23756 47738 23808 47744
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 24136 45082 24164 50866
rect 22744 45076 22796 45082
rect 22744 45018 22796 45024
rect 24124 45076 24176 45082
rect 24124 45018 24176 45024
rect 24492 44872 24544 44878
rect 24492 44814 24544 44820
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22744 43716 22796 43722
rect 22744 43658 22796 43664
rect 22560 42220 22612 42226
rect 22560 42162 22612 42168
rect 22112 41386 22324 41414
rect 22388 41386 22508 41414
rect 22008 40724 22060 40730
rect 22008 40666 22060 40672
rect 22112 38554 22140 41386
rect 22388 41070 22416 41386
rect 22468 41200 22520 41206
rect 22468 41142 22520 41148
rect 22376 41064 22428 41070
rect 22376 41006 22428 41012
rect 22192 40384 22244 40390
rect 22192 40326 22244 40332
rect 22100 38548 22152 38554
rect 22100 38490 22152 38496
rect 22100 38276 22152 38282
rect 22100 38218 22152 38224
rect 22112 37942 22140 38218
rect 22100 37936 22152 37942
rect 22100 37878 22152 37884
rect 22112 36854 22140 37878
rect 22204 37126 22232 40326
rect 22284 39500 22336 39506
rect 22284 39442 22336 39448
rect 22192 37120 22244 37126
rect 22192 37062 22244 37068
rect 22100 36848 22152 36854
rect 22100 36790 22152 36796
rect 22008 36780 22060 36786
rect 22008 36722 22060 36728
rect 21916 36304 21968 36310
rect 21916 36246 21968 36252
rect 21824 36100 21876 36106
rect 21824 36042 21876 36048
rect 21836 35894 21864 36042
rect 21836 35866 21956 35894
rect 21364 35828 21416 35834
rect 21364 35770 21416 35776
rect 21928 35766 21956 35866
rect 21916 35760 21968 35766
rect 21916 35702 21968 35708
rect 21732 35080 21784 35086
rect 21732 35022 21784 35028
rect 21744 33454 21772 35022
rect 21928 34950 21956 35702
rect 22020 35290 22048 36722
rect 22008 35284 22060 35290
rect 22008 35226 22060 35232
rect 22100 35148 22152 35154
rect 22296 35136 22324 39442
rect 22480 39438 22508 41142
rect 22468 39432 22520 39438
rect 22468 39374 22520 39380
rect 22376 38412 22428 38418
rect 22376 38354 22428 38360
rect 22388 36378 22416 38354
rect 22468 37664 22520 37670
rect 22468 37606 22520 37612
rect 22480 37262 22508 37606
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22376 36372 22428 36378
rect 22376 36314 22428 36320
rect 22152 35108 22324 35136
rect 22100 35090 22152 35096
rect 21916 34944 21968 34950
rect 21916 34886 21968 34892
rect 22388 34406 22416 36314
rect 22466 35048 22522 35057
rect 22466 34983 22522 34992
rect 22376 34400 22428 34406
rect 22376 34342 22428 34348
rect 21732 33448 21784 33454
rect 21088 33390 21140 33396
rect 21270 33416 21326 33425
rect 21100 32910 21128 33390
rect 21732 33390 21784 33396
rect 21270 33351 21326 33360
rect 22376 33312 22428 33318
rect 22376 33254 22428 33260
rect 22388 32978 22416 33254
rect 22376 32972 22428 32978
rect 22376 32914 22428 32920
rect 21088 32904 21140 32910
rect 21088 32846 21140 32852
rect 20260 32224 20312 32230
rect 20260 32166 20312 32172
rect 18708 31726 19104 31754
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18708 30122 18736 31726
rect 18696 30116 18748 30122
rect 18696 30058 18748 30064
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18604 20324 18656 20330
rect 18604 20266 18656 20272
rect 18616 19922 18644 20266
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17328 2990 17356 19790
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18616 8498 18644 16594
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17972 3097 18000 3130
rect 17958 3088 18014 3097
rect 17684 3052 17736 3058
rect 17958 3023 18014 3032
rect 17684 2994 17736 3000
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14476 2038 14504 2586
rect 16580 2576 16632 2582
rect 16408 2524 16580 2530
rect 16408 2518 16632 2524
rect 16408 2514 16620 2518
rect 16396 2508 16620 2514
rect 16448 2502 16620 2508
rect 16396 2450 16448 2456
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 14752 800 14780 2382
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 16212 2372 16264 2378
rect 16212 2314 16264 2320
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 2009 15332 2246
rect 15290 2000 15346 2009
rect 15290 1935 15346 1944
rect 15488 800 15516 2314
rect 16224 800 16252 2314
rect 16316 1970 16344 2314
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16960 800 16988 2314
rect 17512 1698 17540 2382
rect 17500 1692 17552 1698
rect 17500 1634 17552 1640
rect 17696 800 17724 2994
rect 18708 2650 18736 30058
rect 21100 29714 21128 32846
rect 22480 31754 22508 34983
rect 22572 34134 22600 42162
rect 22652 41676 22704 41682
rect 22652 41618 22704 41624
rect 22664 40050 22692 41618
rect 22652 40044 22704 40050
rect 22652 39986 22704 39992
rect 22664 36786 22692 39986
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 22664 34610 22692 36722
rect 22756 35193 22784 43658
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 24400 42152 24452 42158
rect 24400 42094 24452 42100
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 23664 41812 23716 41818
rect 23664 41754 23716 41760
rect 22928 41744 22980 41750
rect 22928 41686 22980 41692
rect 22940 41274 22968 41686
rect 23676 41682 23704 41754
rect 23664 41676 23716 41682
rect 23664 41618 23716 41624
rect 24412 41414 24440 42094
rect 24320 41386 24440 41414
rect 22928 41268 22980 41274
rect 22928 41210 22980 41216
rect 24320 41070 24348 41386
rect 24308 41064 24360 41070
rect 24308 41006 24360 41012
rect 23388 40928 23440 40934
rect 23388 40870 23440 40876
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 23400 39030 23428 40870
rect 23480 40452 23532 40458
rect 23480 40394 23532 40400
rect 23388 39024 23440 39030
rect 23388 38966 23440 38972
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23296 37256 23348 37262
rect 23294 37224 23296 37233
rect 23348 37224 23350 37233
rect 23294 37159 23350 37168
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 23400 36242 23428 38966
rect 23492 37126 23520 40394
rect 23572 39976 23624 39982
rect 23572 39918 23624 39924
rect 23584 39302 23612 39918
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 23572 39296 23624 39302
rect 23572 39238 23624 39244
rect 23584 37330 23612 39238
rect 23676 39098 23704 39782
rect 23664 39092 23716 39098
rect 23664 39034 23716 39040
rect 24124 38004 24176 38010
rect 24124 37946 24176 37952
rect 23572 37324 23624 37330
rect 23572 37266 23624 37272
rect 23480 37120 23532 37126
rect 23480 37062 23532 37068
rect 24136 36854 24164 37946
rect 24124 36848 24176 36854
rect 24124 36790 24176 36796
rect 23664 36576 23716 36582
rect 23664 36518 23716 36524
rect 23572 36304 23624 36310
rect 23572 36246 23624 36252
rect 23388 36236 23440 36242
rect 23388 36178 23440 36184
rect 23584 36038 23612 36246
rect 23676 36174 23704 36518
rect 24320 36242 24348 41006
rect 24400 39568 24452 39574
rect 24400 39510 24452 39516
rect 24412 37194 24440 39510
rect 24504 39098 24532 44814
rect 24676 42696 24728 42702
rect 24676 42638 24728 42644
rect 24688 42294 24716 42638
rect 24860 42560 24912 42566
rect 24860 42502 24912 42508
rect 24872 42294 24900 42502
rect 24676 42288 24728 42294
rect 24676 42230 24728 42236
rect 24860 42288 24912 42294
rect 24860 42230 24912 42236
rect 24688 41478 24716 42230
rect 24872 42022 24900 42230
rect 24860 42016 24912 42022
rect 24860 41958 24912 41964
rect 24676 41472 24728 41478
rect 24676 41414 24728 41420
rect 24596 41386 24716 41414
rect 24596 41070 24624 41386
rect 24872 41274 24900 41958
rect 24860 41268 24912 41274
rect 24860 41210 24912 41216
rect 24584 41064 24636 41070
rect 24584 41006 24636 41012
rect 25044 41064 25096 41070
rect 25044 41006 25096 41012
rect 24596 39506 24624 41006
rect 25056 40594 25084 41006
rect 25044 40588 25096 40594
rect 25044 40530 25096 40536
rect 25056 40186 25084 40530
rect 25044 40180 25096 40186
rect 25044 40122 25096 40128
rect 24584 39500 24636 39506
rect 24584 39442 24636 39448
rect 24952 39500 25004 39506
rect 24952 39442 25004 39448
rect 24492 39092 24544 39098
rect 24492 39034 24544 39040
rect 24964 38978 24992 39442
rect 25136 39364 25188 39370
rect 25136 39306 25188 39312
rect 24860 38956 24912 38962
rect 24964 38950 25084 38978
rect 25148 38962 25176 39306
rect 24860 38898 24912 38904
rect 24768 38888 24820 38894
rect 24768 38830 24820 38836
rect 24780 38350 24808 38830
rect 24768 38344 24820 38350
rect 24768 38286 24820 38292
rect 24676 37664 24728 37670
rect 24676 37606 24728 37612
rect 24688 37398 24716 37606
rect 24676 37392 24728 37398
rect 24676 37334 24728 37340
rect 24584 37324 24636 37330
rect 24584 37266 24636 37272
rect 24400 37188 24452 37194
rect 24400 37130 24452 37136
rect 24308 36236 24360 36242
rect 24308 36178 24360 36184
rect 23664 36168 23716 36174
rect 23664 36110 23716 36116
rect 23572 36032 23624 36038
rect 23572 35974 23624 35980
rect 23296 35624 23348 35630
rect 23296 35566 23348 35572
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 22742 35184 22798 35193
rect 23308 35154 23336 35566
rect 22742 35119 22798 35128
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 22652 34604 22704 34610
rect 22652 34546 22704 34552
rect 22560 34128 22612 34134
rect 22560 34070 22612 34076
rect 22664 32434 22692 34546
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22652 32428 22704 32434
rect 22652 32370 22704 32376
rect 22664 32026 22692 32370
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 22480 31726 22600 31754
rect 22468 31272 22520 31278
rect 22466 31240 22468 31249
rect 22520 31240 22522 31249
rect 22466 31175 22522 31184
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 21836 30734 21864 31078
rect 22098 30832 22154 30841
rect 22098 30767 22100 30776
rect 22152 30767 22154 30776
rect 22100 30738 22152 30744
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 22192 30660 22244 30666
rect 22192 30602 22244 30608
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 21180 30252 21232 30258
rect 21180 30194 21232 30200
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 21192 29578 21220 30194
rect 21180 29572 21232 29578
rect 21180 29514 21232 29520
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22642 18920 22918
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 19352 20942 19380 28358
rect 21192 28150 21220 29514
rect 21180 28144 21232 28150
rect 21180 28086 21232 28092
rect 21456 28008 21508 28014
rect 21456 27950 21508 27956
rect 21364 24880 21416 24886
rect 21364 24822 21416 24828
rect 19708 24744 19760 24750
rect 19708 24686 19760 24692
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 19720 24274 19748 24686
rect 21088 24676 21140 24682
rect 21088 24618 21140 24624
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19720 23186 19748 24210
rect 21100 24138 21128 24618
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19616 21616 19668 21622
rect 19616 21558 19668 21564
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 21026 19564 21286
rect 19444 20998 19564 21026
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19444 19922 19472 20998
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19260 17134 19288 17614
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19260 16658 19288 17070
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19260 8566 19288 16390
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18340 1902 18368 2382
rect 18328 1896 18380 1902
rect 18328 1838 18380 1844
rect 18432 800 18460 2450
rect 19168 800 19196 2926
rect 19536 1834 19564 20878
rect 19628 19922 19656 21558
rect 19720 21010 19748 22986
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19904 21146 19932 22510
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 19892 21140 19944 21146
rect 19892 21082 19944 21088
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19892 20800 19944 20806
rect 19892 20742 19944 20748
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19812 16522 19840 19722
rect 19904 18970 19932 20742
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19996 17762 20024 19994
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20088 17882 20116 19382
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19996 17734 20116 17762
rect 20548 17746 20576 19994
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 19812 11218 19840 16458
rect 19996 16250 20024 17478
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19996 3126 20024 16186
rect 20088 15162 20116 17734
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 14618 20576 14758
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 19524 1828 19576 1834
rect 19524 1770 19576 1776
rect 19904 800 19932 2382
rect 20640 800 20668 2926
rect 20732 2650 20760 21898
rect 20824 21622 20852 23054
rect 20916 21894 20944 23598
rect 21008 21962 21036 23734
rect 21100 22166 21128 24074
rect 21284 24070 21312 24686
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21284 23662 21312 24006
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 21376 23186 21404 24822
rect 21468 24274 21496 27950
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21468 23730 21496 24210
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21560 23594 21588 24550
rect 21836 24410 21864 30534
rect 22204 28762 22232 30602
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 22388 29034 22416 29106
rect 22376 29028 22428 29034
rect 22376 28970 22428 28976
rect 22192 28756 22244 28762
rect 22192 28698 22244 28704
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22112 26450 22140 28018
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 22388 25838 22416 28970
rect 22572 28626 22600 31726
rect 22756 30938 22784 33798
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23308 33114 23336 35090
rect 22836 33108 22888 33114
rect 22836 33050 22888 33056
rect 23296 33108 23348 33114
rect 23296 33050 23348 33056
rect 22848 32366 22876 33050
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 22836 32360 22888 32366
rect 22836 32302 22888 32308
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23204 31680 23256 31686
rect 23204 31622 23256 31628
rect 22836 31340 22888 31346
rect 22836 31282 22888 31288
rect 22744 30932 22796 30938
rect 22744 30874 22796 30880
rect 22848 30870 22876 31282
rect 23216 31142 23244 31622
rect 23492 31414 23520 32370
rect 23480 31408 23532 31414
rect 23480 31350 23532 31356
rect 23584 31362 23612 35974
rect 24320 34474 24348 36178
rect 24596 36106 24624 37266
rect 24584 36100 24636 36106
rect 24584 36042 24636 36048
rect 24596 34950 24624 36042
rect 24688 35698 24716 37334
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 24676 35692 24728 35698
rect 24676 35634 24728 35640
rect 24780 35018 24808 35770
rect 24768 35012 24820 35018
rect 24768 34954 24820 34960
rect 24584 34944 24636 34950
rect 24584 34886 24636 34892
rect 24308 34468 24360 34474
rect 24308 34410 24360 34416
rect 24032 34060 24084 34066
rect 24032 34002 24084 34008
rect 24044 33658 24072 34002
rect 24032 33652 24084 33658
rect 24032 33594 24084 33600
rect 23664 32972 23716 32978
rect 23664 32914 23716 32920
rect 23676 32774 23704 32914
rect 23664 32768 23716 32774
rect 23664 32710 23716 32716
rect 23676 31822 23704 32710
rect 23756 32496 23808 32502
rect 23756 32438 23808 32444
rect 23768 31958 23796 32438
rect 24044 32026 24072 33594
rect 24596 33454 24624 34886
rect 24780 34678 24808 34954
rect 24872 34746 24900 38898
rect 24952 38888 25004 38894
rect 24952 38830 25004 38836
rect 24964 37670 24992 38830
rect 25056 38486 25084 38950
rect 25136 38956 25188 38962
rect 25136 38898 25188 38904
rect 25044 38480 25096 38486
rect 25044 38422 25096 38428
rect 25044 38344 25096 38350
rect 25044 38286 25096 38292
rect 25056 38010 25084 38286
rect 25136 38276 25188 38282
rect 25136 38218 25188 38224
rect 25044 38004 25096 38010
rect 25044 37946 25096 37952
rect 24952 37664 25004 37670
rect 24952 37606 25004 37612
rect 24964 36718 24992 37606
rect 24952 36712 25004 36718
rect 24952 36654 25004 36660
rect 25056 35630 25084 37946
rect 25044 35624 25096 35630
rect 25044 35566 25096 35572
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 24768 34672 24820 34678
rect 24768 34614 24820 34620
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 24584 33448 24636 33454
rect 24584 33390 24636 33396
rect 24124 32360 24176 32366
rect 24124 32302 24176 32308
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 23756 31952 23808 31958
rect 23756 31894 23808 31900
rect 23940 31884 23992 31890
rect 23940 31826 23992 31832
rect 24032 31884 24084 31890
rect 24032 31826 24084 31832
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 23848 31816 23900 31822
rect 23848 31758 23900 31764
rect 23860 31482 23888 31758
rect 23952 31482 23980 31826
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23940 31476 23992 31482
rect 23940 31418 23992 31424
rect 23296 31340 23348 31346
rect 23584 31334 23704 31362
rect 23296 31282 23348 31288
rect 23204 31136 23256 31142
rect 23204 31078 23256 31084
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22836 30864 22888 30870
rect 22836 30806 22888 30812
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22560 28620 22612 28626
rect 22560 28562 22612 28568
rect 22572 28506 22600 28562
rect 22480 28478 22600 28506
rect 22376 25832 22428 25838
rect 22376 25774 22428 25780
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21836 23798 21864 24346
rect 21824 23792 21876 23798
rect 21824 23734 21876 23740
rect 21548 23588 21600 23594
rect 21548 23530 21600 23536
rect 22100 23520 22152 23526
rect 22100 23462 22152 23468
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21192 22574 21220 22918
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20812 21616 20864 21622
rect 20864 21576 20944 21604
rect 20812 21558 20864 21564
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20824 2774 20852 20402
rect 20916 19786 20944 21576
rect 21192 20602 21220 22374
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21008 18970 21036 19314
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21192 18426 21220 20198
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 19310 21312 19654
rect 21376 19514 21404 22442
rect 22112 21894 22140 23462
rect 22192 23044 22244 23050
rect 22192 22986 22244 22992
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21468 19378 21496 19654
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20916 17338 20944 18090
rect 21008 17746 21036 18158
rect 20996 17740 21048 17746
rect 20996 17682 21048 17688
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21100 16454 21128 17138
rect 21284 17066 21312 18294
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 14958 21220 16390
rect 21376 15638 21404 18566
rect 21468 18358 21496 19314
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21468 17338 21496 17682
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21364 15632 21416 15638
rect 21364 15574 21416 15580
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21376 3466 21404 15574
rect 21560 8430 21588 19246
rect 21744 18766 21772 19382
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21928 17134 21956 20334
rect 21916 17128 21968 17134
rect 21916 17070 21968 17076
rect 21928 16658 21956 17070
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 20824 2746 21128 2774
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20824 2310 20852 2586
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20916 1834 20944 2382
rect 20996 2304 21048 2310
rect 20996 2246 21048 2252
rect 21008 2038 21036 2246
rect 20996 2032 21048 2038
rect 20996 1974 21048 1980
rect 20904 1828 20956 1834
rect 20904 1770 20956 1776
rect 21100 1766 21128 2746
rect 21364 2508 21416 2514
rect 21364 2450 21416 2456
rect 21088 1760 21140 1766
rect 21088 1702 21140 1708
rect 21376 800 21404 2450
rect 22112 800 22140 2926
rect 22204 2650 22232 22986
rect 22296 22778 22324 25094
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22296 19378 22324 21898
rect 22388 20466 22416 25774
rect 22480 23526 22508 28478
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 22572 27062 22600 28358
rect 22560 27056 22612 27062
rect 22560 26998 22612 27004
rect 22652 25152 22704 25158
rect 22652 25094 22704 25100
rect 22664 24818 22692 25094
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22480 21570 22508 23462
rect 22572 22166 22600 24006
rect 22756 23050 22784 29446
rect 23308 29306 23336 31282
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 23296 29300 23348 29306
rect 23296 29242 23348 29248
rect 23294 29200 23350 29209
rect 23294 29135 23296 29144
rect 23348 29135 23350 29144
rect 23296 29106 23348 29112
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 23400 28626 23428 30670
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23584 30190 23612 30534
rect 23572 30184 23624 30190
rect 23572 30126 23624 30132
rect 23676 29510 23704 31334
rect 23952 30802 23980 31418
rect 23940 30796 23992 30802
rect 23940 30738 23992 30744
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23388 28620 23440 28626
rect 23388 28562 23440 28568
rect 23846 28112 23902 28121
rect 23846 28047 23848 28056
rect 23900 28047 23902 28056
rect 23848 28018 23900 28024
rect 23388 28008 23440 28014
rect 23388 27950 23440 27956
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 23124 27130 23152 27406
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 23400 26926 23428 27950
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 23768 26382 23796 26454
rect 23756 26376 23808 26382
rect 23756 26318 23808 26324
rect 23664 26308 23716 26314
rect 23664 26250 23716 26256
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22560 22160 22612 22166
rect 22560 22102 22612 22108
rect 22664 21672 22692 22918
rect 22664 21644 22784 21672
rect 22480 21542 22692 21570
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22480 20466 22508 21422
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22480 19922 22508 20402
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22480 19446 22508 19858
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22388 17746 22416 18770
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22480 18086 22508 18634
rect 22572 18222 22600 18634
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22572 17490 22600 18158
rect 22480 17462 22600 17490
rect 22480 16794 22508 17462
rect 22664 17354 22692 21542
rect 22756 17542 22784 21644
rect 22848 21486 22876 24142
rect 23308 23866 23336 25094
rect 23676 24886 23704 26250
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23676 24138 23704 24822
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23676 23798 23704 24074
rect 23664 23792 23716 23798
rect 23492 23752 23664 23780
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22234 23336 22578
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 22848 18834 22876 21422
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23308 19446 23336 20470
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 23308 19310 23336 19382
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23400 18970 23428 22646
rect 23492 21622 23520 23752
rect 23664 23734 23716 23740
rect 23664 23588 23716 23594
rect 23664 23530 23716 23536
rect 23676 23186 23704 23530
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23584 21690 23612 21898
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23676 21570 23704 22714
rect 23768 21672 23796 26318
rect 23860 26314 23888 28018
rect 24044 26874 24072 31826
rect 24136 31278 24164 32302
rect 24124 31272 24176 31278
rect 24124 31214 24176 31220
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24136 30870 24164 31214
rect 24124 30864 24176 30870
rect 24124 30806 24176 30812
rect 24596 30734 24624 31214
rect 24688 31210 24716 33798
rect 24780 33590 24808 34614
rect 24860 34536 24912 34542
rect 24860 34478 24912 34484
rect 24768 33584 24820 33590
rect 24768 33526 24820 33532
rect 24780 32774 24808 33526
rect 24768 32768 24820 32774
rect 24768 32710 24820 32716
rect 24780 32502 24808 32710
rect 24768 32496 24820 32502
rect 24768 32438 24820 32444
rect 24780 32366 24808 32438
rect 24768 32360 24820 32366
rect 24768 32302 24820 32308
rect 24872 31754 24900 34478
rect 24860 31748 24912 31754
rect 24860 31690 24912 31696
rect 24768 31408 24820 31414
rect 24768 31350 24820 31356
rect 24676 31204 24728 31210
rect 24676 31146 24728 31152
rect 24780 30802 24808 31350
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24780 30326 24808 30738
rect 24872 30666 24900 31690
rect 24952 31136 25004 31142
rect 25056 31124 25084 35566
rect 25148 33658 25176 38218
rect 25136 33652 25188 33658
rect 25136 33594 25188 33600
rect 25136 33516 25188 33522
rect 25136 33458 25188 33464
rect 25004 31096 25084 31124
rect 24952 31078 25004 31084
rect 25148 30938 25176 33458
rect 25240 32586 25268 53994
rect 26056 53984 26108 53990
rect 26056 53926 26108 53932
rect 26240 53984 26292 53990
rect 26240 53926 26292 53932
rect 27436 53984 27488 53990
rect 27436 53926 27488 53932
rect 28540 53984 28592 53990
rect 28540 53926 28592 53932
rect 25780 53508 25832 53514
rect 25780 53450 25832 53456
rect 25320 41200 25372 41206
rect 25320 41142 25372 41148
rect 25332 40118 25360 41142
rect 25320 40112 25372 40118
rect 25320 40054 25372 40060
rect 25332 39370 25360 40054
rect 25320 39364 25372 39370
rect 25320 39306 25372 39312
rect 25504 38208 25556 38214
rect 25504 38150 25556 38156
rect 25516 37126 25544 38150
rect 25412 37120 25464 37126
rect 25412 37062 25464 37068
rect 25504 37120 25556 37126
rect 25504 37062 25556 37068
rect 25424 36768 25452 37062
rect 25504 36780 25556 36786
rect 25424 36740 25504 36768
rect 25504 36722 25556 36728
rect 25596 36712 25648 36718
rect 25596 36654 25648 36660
rect 25608 35018 25636 36654
rect 25596 35012 25648 35018
rect 25596 34954 25648 34960
rect 25608 34746 25636 34954
rect 25596 34740 25648 34746
rect 25596 34682 25648 34688
rect 25688 34604 25740 34610
rect 25688 34546 25740 34552
rect 25596 34060 25648 34066
rect 25596 34002 25648 34008
rect 25240 32558 25360 32586
rect 25608 32570 25636 34002
rect 25332 31754 25360 32558
rect 25596 32564 25648 32570
rect 25596 32506 25648 32512
rect 25332 31726 25452 31754
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 25136 30660 25188 30666
rect 25136 30602 25188 30608
rect 24768 30320 24820 30326
rect 24768 30262 24820 30268
rect 25148 29102 25176 30602
rect 25424 30598 25452 31726
rect 25700 31686 25728 34546
rect 25688 31680 25740 31686
rect 25688 31622 25740 31628
rect 25792 31142 25820 53450
rect 25872 47660 25924 47666
rect 25872 47602 25924 47608
rect 25884 43450 25912 47602
rect 25872 43444 25924 43450
rect 25872 43386 25924 43392
rect 25964 43308 26016 43314
rect 25964 43250 26016 43256
rect 25872 42628 25924 42634
rect 25872 42570 25924 42576
rect 25884 42022 25912 42570
rect 25872 42016 25924 42022
rect 25872 41958 25924 41964
rect 25884 41750 25912 41958
rect 25872 41744 25924 41750
rect 25872 41686 25924 41692
rect 25884 38894 25912 41686
rect 25976 39098 26004 43250
rect 25964 39092 26016 39098
rect 25964 39034 26016 39040
rect 25872 38888 25924 38894
rect 25872 38830 25924 38836
rect 25964 38820 26016 38826
rect 25964 38762 26016 38768
rect 25872 36576 25924 36582
rect 25872 36518 25924 36524
rect 25780 31136 25832 31142
rect 25780 31078 25832 31084
rect 25412 30592 25464 30598
rect 25412 30534 25464 30540
rect 25136 29096 25188 29102
rect 25136 29038 25188 29044
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 24964 28150 24992 28494
rect 24952 28144 25004 28150
rect 24952 28086 25004 28092
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 24044 26846 24164 26874
rect 24032 26784 24084 26790
rect 24032 26726 24084 26732
rect 23848 26308 23900 26314
rect 23848 26250 23900 26256
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23860 21962 23888 24006
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23768 21644 23980 21672
rect 23492 20534 23520 21558
rect 23676 21542 23796 21570
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23492 19786 23520 20470
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23584 19174 23612 19654
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23584 18834 23612 19110
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22572 17326 22692 17354
rect 22848 17338 22876 18226
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23216 17338 23244 17614
rect 23584 17610 23612 18294
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 22836 17332 22888 17338
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22480 16046 22508 16730
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 22480 15026 22508 15982
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22572 2106 22600 17326
rect 22836 17274 22888 17280
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23308 17218 23336 17546
rect 23216 17202 23336 17218
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23204 17196 23336 17202
rect 23256 17190 23336 17196
rect 23204 17138 23256 17144
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 16522 23336 17190
rect 23400 16794 23428 17206
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22664 2446 22692 15302
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22560 2100 22612 2106
rect 22560 2042 22612 2048
rect 22848 800 22876 2450
rect 23584 800 23612 2926
rect 23676 2378 23704 19382
rect 23664 2372 23716 2378
rect 23664 2314 23716 2320
rect 23768 2310 23796 21542
rect 23952 21350 23980 21644
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 23952 19378 23980 19790
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 24044 17202 24072 26726
rect 24136 19446 24164 26846
rect 24228 26518 24256 27814
rect 24964 27538 24992 28086
rect 24952 27532 25004 27538
rect 24952 27474 25004 27480
rect 25228 27396 25280 27402
rect 25228 27338 25280 27344
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 24216 26512 24268 26518
rect 24216 26454 24268 26460
rect 25056 26450 25084 26522
rect 25044 26444 25096 26450
rect 25044 26386 25096 26392
rect 24584 26240 24636 26246
rect 24584 26182 24636 26188
rect 24216 25356 24268 25362
rect 24216 25298 24268 25304
rect 24228 22098 24256 25298
rect 24216 22092 24268 22098
rect 24216 22034 24268 22040
rect 24228 21350 24256 22034
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24228 21010 24256 21286
rect 24216 21004 24268 21010
rect 24216 20946 24268 20952
rect 24596 20262 24624 26182
rect 25240 25838 25268 27338
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 25228 25832 25280 25838
rect 25228 25774 25280 25780
rect 25240 25498 25268 25774
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25136 25356 25188 25362
rect 25136 25298 25188 25304
rect 25148 24682 25176 25298
rect 25136 24676 25188 24682
rect 25136 24618 25188 24624
rect 24676 23588 24728 23594
rect 24676 23530 24728 23536
rect 24584 20256 24636 20262
rect 24584 20198 24636 20204
rect 24688 20074 24716 23530
rect 24952 23520 25004 23526
rect 24858 23488 24914 23497
rect 24952 23462 25004 23468
rect 24858 23423 24914 23432
rect 24872 23118 24900 23423
rect 24964 23118 24992 23462
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24780 22642 24808 22986
rect 24952 22976 25004 22982
rect 25044 22976 25096 22982
rect 24952 22918 25004 22924
rect 25042 22944 25044 22953
rect 25096 22944 25098 22953
rect 24964 22778 24992 22918
rect 25042 22879 25098 22888
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 25044 22432 25096 22438
rect 25044 22374 25096 22380
rect 25056 22234 25084 22374
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 24952 21888 25004 21894
rect 24952 21830 25004 21836
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24596 20046 24716 20074
rect 24216 19780 24268 19786
rect 24216 19722 24268 19728
rect 24228 19446 24256 19722
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24228 19334 24256 19382
rect 24400 19372 24452 19378
rect 24228 19306 24348 19334
rect 24400 19314 24452 19320
rect 24320 18426 24348 19306
rect 24308 18420 24360 18426
rect 24308 18362 24360 18368
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 24308 17196 24360 17202
rect 24308 17138 24360 17144
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24136 3058 24164 15506
rect 24320 10742 24348 17138
rect 24412 16658 24440 19314
rect 24596 19242 24624 20046
rect 24584 19236 24636 19242
rect 24584 19178 24636 19184
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24688 16182 24716 18838
rect 24780 18834 24808 21286
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 24872 18766 24900 20198
rect 24964 20058 24992 21830
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24964 18426 24992 18566
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 25056 18358 25084 22170
rect 25148 21554 25176 24618
rect 25228 23180 25280 23186
rect 25228 23122 25280 23128
rect 25240 22438 25268 23122
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 25228 22160 25280 22166
rect 25228 22102 25280 22108
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25148 20602 25176 21490
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25148 19922 25176 20538
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 25056 17270 25084 18294
rect 25044 17264 25096 17270
rect 25044 17206 25096 17212
rect 25056 16658 25084 17206
rect 24768 16652 24820 16658
rect 25044 16652 25096 16658
rect 24820 16612 24900 16640
rect 24768 16594 24820 16600
rect 24768 16516 24820 16522
rect 24768 16458 24820 16464
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24584 13184 24636 13190
rect 24584 13126 24636 13132
rect 24308 10736 24360 10742
rect 24308 10678 24360 10684
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 24320 800 24348 3538
rect 24596 3534 24624 13126
rect 24688 4622 24716 16118
rect 24780 16046 24808 16458
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24780 15094 24808 15982
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24780 14278 24808 15030
rect 24872 14482 24900 16612
rect 25044 16594 25096 16600
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 25240 13326 25268 22102
rect 25332 15434 25360 26522
rect 25424 15434 25452 30534
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25516 28490 25544 30194
rect 25608 29850 25636 30194
rect 25596 29844 25648 29850
rect 25596 29786 25648 29792
rect 25504 28484 25556 28490
rect 25504 28426 25556 28432
rect 25504 25220 25556 25226
rect 25504 25162 25556 25168
rect 25516 24562 25544 25162
rect 25608 24750 25636 29786
rect 25688 29028 25740 29034
rect 25688 28970 25740 28976
rect 25700 25226 25728 28970
rect 25792 26586 25820 31078
rect 25884 27062 25912 36518
rect 25976 35290 26004 38762
rect 26068 35850 26096 53926
rect 26252 43790 26280 53926
rect 27068 53712 27120 53718
rect 27068 53654 27120 53660
rect 26700 51400 26752 51406
rect 26700 51342 26752 51348
rect 26712 46170 26740 51342
rect 26700 46164 26752 46170
rect 26700 46106 26752 46112
rect 26240 43784 26292 43790
rect 26240 43726 26292 43732
rect 26332 43240 26384 43246
rect 26332 43182 26384 43188
rect 26344 41818 26372 43182
rect 26332 41812 26384 41818
rect 26332 41754 26384 41760
rect 26424 41608 26476 41614
rect 26424 41550 26476 41556
rect 26148 39364 26200 39370
rect 26148 39306 26200 39312
rect 26160 38962 26188 39306
rect 26240 39092 26292 39098
rect 26292 39052 26372 39080
rect 26240 39034 26292 39040
rect 26148 38956 26200 38962
rect 26148 38898 26200 38904
rect 26240 38956 26292 38962
rect 26240 38898 26292 38904
rect 26252 36378 26280 38898
rect 26344 38554 26372 39052
rect 26332 38548 26384 38554
rect 26332 38490 26384 38496
rect 26436 36718 26464 41550
rect 26608 40928 26660 40934
rect 26608 40870 26660 40876
rect 26620 40594 26648 40870
rect 26608 40588 26660 40594
rect 26608 40530 26660 40536
rect 27080 40526 27108 53654
rect 27160 44872 27212 44878
rect 27160 44814 27212 44820
rect 26976 40520 27028 40526
rect 26976 40462 27028 40468
rect 27068 40520 27120 40526
rect 27068 40462 27120 40468
rect 26884 40384 26936 40390
rect 26884 40326 26936 40332
rect 26700 38344 26752 38350
rect 26700 38286 26752 38292
rect 26712 37806 26740 38286
rect 26700 37800 26752 37806
rect 26700 37742 26752 37748
rect 26792 37800 26844 37806
rect 26792 37742 26844 37748
rect 26424 36712 26476 36718
rect 26424 36654 26476 36660
rect 26240 36372 26292 36378
rect 26240 36314 26292 36320
rect 26608 36168 26660 36174
rect 26608 36110 26660 36116
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 26068 35822 26188 35850
rect 25964 35284 26016 35290
rect 25964 35226 26016 35232
rect 26056 33924 26108 33930
rect 26056 33866 26108 33872
rect 26068 33046 26096 33866
rect 26056 33040 26108 33046
rect 26056 32982 26108 32988
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 25964 32224 26016 32230
rect 25964 32166 26016 32172
rect 25976 31754 26004 32166
rect 26068 31890 26096 32506
rect 26056 31884 26108 31890
rect 26056 31826 26108 31832
rect 25976 31726 26096 31754
rect 26068 30326 26096 31726
rect 26056 30320 26108 30326
rect 26056 30262 26108 30268
rect 26068 28200 26096 30262
rect 26160 29034 26188 35822
rect 26252 35086 26280 35974
rect 26424 35828 26476 35834
rect 26424 35770 26476 35776
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 26332 35012 26384 35018
rect 26332 34954 26384 34960
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 26252 30734 26280 31282
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26148 29028 26200 29034
rect 26148 28970 26200 28976
rect 26068 28172 26188 28200
rect 25872 27056 25924 27062
rect 25872 26998 25924 27004
rect 25780 26580 25832 26586
rect 25780 26522 25832 26528
rect 25780 25696 25832 25702
rect 25780 25638 25832 25644
rect 25872 25696 25924 25702
rect 25872 25638 25924 25644
rect 25792 25362 25820 25638
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25688 25220 25740 25226
rect 25688 25162 25740 25168
rect 25884 24886 25912 25638
rect 25964 25288 26016 25294
rect 26160 25276 26188 28172
rect 26252 28150 26280 30670
rect 26344 30122 26372 34954
rect 26436 34542 26464 35770
rect 26620 35018 26648 36110
rect 26712 35834 26740 37742
rect 26804 37262 26832 37742
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26700 35828 26752 35834
rect 26700 35770 26752 35776
rect 26804 35698 26832 37198
rect 26792 35692 26844 35698
rect 26792 35634 26844 35640
rect 26804 35154 26832 35634
rect 26896 35578 26924 40326
rect 26988 38486 27016 40462
rect 27172 39098 27200 44814
rect 27344 43240 27396 43246
rect 27344 43182 27396 43188
rect 27356 42906 27384 43182
rect 27344 42900 27396 42906
rect 27344 42842 27396 42848
rect 27356 42294 27384 42842
rect 27344 42288 27396 42294
rect 27344 42230 27396 42236
rect 27252 42152 27304 42158
rect 27252 42094 27304 42100
rect 27264 41478 27292 42094
rect 27252 41472 27304 41478
rect 27252 41414 27304 41420
rect 27448 41414 27476 53926
rect 27950 53340 28258 53349
rect 27950 53338 27956 53340
rect 28012 53338 28036 53340
rect 28092 53338 28116 53340
rect 28172 53338 28196 53340
rect 28252 53338 28258 53340
rect 28012 53286 28014 53338
rect 28194 53286 28196 53338
rect 27950 53284 27956 53286
rect 28012 53284 28036 53286
rect 28092 53284 28116 53286
rect 28172 53284 28196 53286
rect 28252 53284 28258 53286
rect 27950 53275 28258 53284
rect 27950 52252 28258 52261
rect 27950 52250 27956 52252
rect 28012 52250 28036 52252
rect 28092 52250 28116 52252
rect 28172 52250 28196 52252
rect 28252 52250 28258 52252
rect 28012 52198 28014 52250
rect 28194 52198 28196 52250
rect 27950 52196 27956 52198
rect 28012 52196 28036 52198
rect 28092 52196 28116 52198
rect 28172 52196 28196 52198
rect 28252 52196 28258 52198
rect 27950 52187 28258 52196
rect 27950 51164 28258 51173
rect 27950 51162 27956 51164
rect 28012 51162 28036 51164
rect 28092 51162 28116 51164
rect 28172 51162 28196 51164
rect 28252 51162 28258 51164
rect 28012 51110 28014 51162
rect 28194 51110 28196 51162
rect 27950 51108 27956 51110
rect 28012 51108 28036 51110
rect 28092 51108 28116 51110
rect 28172 51108 28196 51110
rect 28252 51108 28258 51110
rect 27950 51099 28258 51108
rect 27950 50076 28258 50085
rect 27950 50074 27956 50076
rect 28012 50074 28036 50076
rect 28092 50074 28116 50076
rect 28172 50074 28196 50076
rect 28252 50074 28258 50076
rect 28012 50022 28014 50074
rect 28194 50022 28196 50074
rect 27950 50020 27956 50022
rect 28012 50020 28036 50022
rect 28092 50020 28116 50022
rect 28172 50020 28196 50022
rect 28252 50020 28258 50022
rect 27950 50011 28258 50020
rect 27950 48988 28258 48997
rect 27950 48986 27956 48988
rect 28012 48986 28036 48988
rect 28092 48986 28116 48988
rect 28172 48986 28196 48988
rect 28252 48986 28258 48988
rect 28012 48934 28014 48986
rect 28194 48934 28196 48986
rect 27950 48932 27956 48934
rect 28012 48932 28036 48934
rect 28092 48932 28116 48934
rect 28172 48932 28196 48934
rect 28252 48932 28258 48934
rect 27950 48923 28258 48932
rect 27950 47900 28258 47909
rect 27950 47898 27956 47900
rect 28012 47898 28036 47900
rect 28092 47898 28116 47900
rect 28172 47898 28196 47900
rect 28252 47898 28258 47900
rect 28012 47846 28014 47898
rect 28194 47846 28196 47898
rect 27950 47844 27956 47846
rect 28012 47844 28036 47846
rect 28092 47844 28116 47846
rect 28172 47844 28196 47846
rect 28252 47844 28258 47846
rect 27950 47835 28258 47844
rect 27950 46812 28258 46821
rect 27950 46810 27956 46812
rect 28012 46810 28036 46812
rect 28092 46810 28116 46812
rect 28172 46810 28196 46812
rect 28252 46810 28258 46812
rect 28012 46758 28014 46810
rect 28194 46758 28196 46810
rect 27950 46756 27956 46758
rect 28012 46756 28036 46758
rect 28092 46756 28116 46758
rect 28172 46756 28196 46758
rect 28252 46756 28258 46758
rect 27950 46747 28258 46756
rect 27804 45960 27856 45966
rect 27804 45902 27856 45908
rect 27620 43648 27672 43654
rect 27620 43590 27672 43596
rect 27264 41138 27292 41414
rect 27356 41386 27476 41414
rect 27252 41132 27304 41138
rect 27252 41074 27304 41080
rect 27252 40996 27304 41002
rect 27252 40938 27304 40944
rect 27160 39092 27212 39098
rect 27160 39034 27212 39040
rect 27264 38554 27292 40938
rect 27252 38548 27304 38554
rect 27252 38490 27304 38496
rect 26976 38480 27028 38486
rect 26976 38422 27028 38428
rect 27264 37466 27292 38490
rect 27252 37460 27304 37466
rect 27252 37402 27304 37408
rect 27068 37324 27120 37330
rect 27068 37266 27120 37272
rect 26976 37188 27028 37194
rect 26976 37130 27028 37136
rect 26988 36106 27016 37130
rect 26976 36100 27028 36106
rect 26976 36042 27028 36048
rect 26896 35550 27016 35578
rect 27080 35562 27108 37266
rect 26884 35488 26936 35494
rect 26884 35430 26936 35436
rect 26896 35290 26924 35430
rect 26884 35284 26936 35290
rect 26884 35226 26936 35232
rect 26792 35148 26844 35154
rect 26792 35090 26844 35096
rect 26608 35012 26660 35018
rect 26608 34954 26660 34960
rect 26804 34610 26832 35090
rect 26792 34604 26844 34610
rect 26792 34546 26844 34552
rect 26424 34536 26476 34542
rect 26424 34478 26476 34484
rect 26804 33930 26832 34546
rect 26988 34082 27016 35550
rect 27068 35556 27120 35562
rect 27068 35498 27120 35504
rect 27080 35222 27108 35498
rect 27356 35476 27384 41386
rect 27436 40588 27488 40594
rect 27436 40530 27488 40536
rect 27264 35448 27384 35476
rect 27068 35216 27120 35222
rect 27068 35158 27120 35164
rect 26988 34054 27108 34082
rect 26792 33924 26844 33930
rect 26792 33866 26844 33872
rect 27080 33454 27108 34054
rect 27068 33448 27120 33454
rect 26790 33416 26846 33425
rect 27068 33390 27120 33396
rect 26790 33351 26846 33360
rect 26804 32978 26832 33351
rect 26792 32972 26844 32978
rect 26792 32914 26844 32920
rect 26804 32881 26832 32914
rect 26884 32904 26936 32910
rect 26790 32872 26846 32881
rect 26884 32846 26936 32852
rect 26790 32807 26846 32816
rect 26608 32768 26660 32774
rect 26608 32710 26660 32716
rect 26620 32502 26648 32710
rect 26608 32496 26660 32502
rect 26608 32438 26660 32444
rect 26424 32292 26476 32298
rect 26424 32234 26476 32240
rect 26436 31754 26464 32234
rect 26436 31748 26568 31754
rect 26436 31726 26516 31748
rect 26516 31690 26568 31696
rect 26528 31346 26556 31690
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26332 30116 26384 30122
rect 26332 30058 26384 30064
rect 26240 28144 26292 28150
rect 26238 28112 26240 28121
rect 26292 28112 26294 28121
rect 26238 28047 26294 28056
rect 26252 27402 26280 28047
rect 26700 28008 26752 28014
rect 26700 27950 26752 27956
rect 26240 27396 26292 27402
rect 26292 27356 26372 27384
rect 26240 27338 26292 27344
rect 26240 25764 26292 25770
rect 26240 25706 26292 25712
rect 25964 25230 26016 25236
rect 26068 25248 26188 25276
rect 25976 24886 26004 25230
rect 25872 24880 25924 24886
rect 25872 24822 25924 24828
rect 25964 24880 26016 24886
rect 25964 24822 26016 24828
rect 25596 24744 25648 24750
rect 25964 24744 26016 24750
rect 25596 24686 25648 24692
rect 25962 24712 25964 24721
rect 26016 24712 26018 24721
rect 25962 24647 26018 24656
rect 25516 24534 25636 24562
rect 25502 24304 25558 24313
rect 25502 24239 25504 24248
rect 25556 24239 25558 24248
rect 25504 24210 25556 24216
rect 25504 22568 25556 22574
rect 25504 22510 25556 22516
rect 25516 20398 25544 22510
rect 25608 22166 25636 24534
rect 26068 23610 26096 25248
rect 26148 25152 26200 25158
rect 26148 25094 26200 25100
rect 26160 24886 26188 25094
rect 26148 24880 26200 24886
rect 26148 24822 26200 24828
rect 26252 24750 26280 25706
rect 26344 25226 26372 27356
rect 26712 27334 26740 27950
rect 26700 27328 26752 27334
rect 26700 27270 26752 27276
rect 26700 27124 26752 27130
rect 26700 27066 26752 27072
rect 26332 25220 26384 25226
rect 26332 25162 26384 25168
rect 26344 24857 26372 25162
rect 26330 24848 26386 24857
rect 26330 24783 26386 24792
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 26608 24064 26660 24070
rect 26608 24006 26660 24012
rect 26160 23730 26188 24006
rect 26620 23798 26648 24006
rect 26608 23792 26660 23798
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 26344 23718 26556 23746
rect 26608 23734 26660 23740
rect 26344 23610 26372 23718
rect 26528 23662 26556 23718
rect 26068 23582 26372 23610
rect 26424 23656 26476 23662
rect 26424 23598 26476 23604
rect 26516 23656 26568 23662
rect 26516 23598 26568 23604
rect 25872 23520 25924 23526
rect 25872 23462 25924 23468
rect 25596 22160 25648 22166
rect 25596 22102 25648 22108
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25608 21622 25636 21830
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25792 21486 25820 22034
rect 25884 21690 25912 23462
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 25780 21480 25832 21486
rect 25780 21422 25832 21428
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 25516 19990 25544 20334
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 25608 18834 25636 21422
rect 25596 18828 25648 18834
rect 25596 18770 25648 18776
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25976 17338 26004 18566
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25412 15428 25464 15434
rect 25412 15370 25464 15376
rect 25884 14890 25912 17138
rect 25872 14884 25924 14890
rect 25872 14826 25924 14832
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25228 12640 25280 12646
rect 25228 12582 25280 12588
rect 25136 10532 25188 10538
rect 25136 10474 25188 10480
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 25148 3058 25176 10474
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 25056 800 25084 2926
rect 25240 2446 25268 12582
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25792 800 25820 2450
rect 26068 1698 26096 23582
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 26160 20602 26188 23462
rect 26436 22094 26464 23598
rect 26712 23508 26740 27066
rect 26896 26246 26924 32846
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 27068 32020 27120 32026
rect 27068 31962 27120 31968
rect 27080 30802 27108 31962
rect 27172 31958 27200 32166
rect 27160 31952 27212 31958
rect 27160 31894 27212 31900
rect 27264 31754 27292 35448
rect 27448 35272 27476 40530
rect 27528 40520 27580 40526
rect 27526 40488 27528 40497
rect 27580 40488 27582 40497
rect 27526 40423 27582 40432
rect 27528 38752 27580 38758
rect 27528 38694 27580 38700
rect 27540 38418 27568 38694
rect 27528 38412 27580 38418
rect 27528 38354 27580 38360
rect 27632 37330 27660 43590
rect 27816 41274 27844 45902
rect 27950 45724 28258 45733
rect 27950 45722 27956 45724
rect 28012 45722 28036 45724
rect 28092 45722 28116 45724
rect 28172 45722 28196 45724
rect 28252 45722 28258 45724
rect 28012 45670 28014 45722
rect 28194 45670 28196 45722
rect 27950 45668 27956 45670
rect 28012 45668 28036 45670
rect 28092 45668 28116 45670
rect 28172 45668 28196 45670
rect 28252 45668 28258 45670
rect 27950 45659 28258 45668
rect 27950 44636 28258 44645
rect 27950 44634 27956 44636
rect 28012 44634 28036 44636
rect 28092 44634 28116 44636
rect 28172 44634 28196 44636
rect 28252 44634 28258 44636
rect 28012 44582 28014 44634
rect 28194 44582 28196 44634
rect 27950 44580 27956 44582
rect 28012 44580 28036 44582
rect 28092 44580 28116 44582
rect 28172 44580 28196 44582
rect 28252 44580 28258 44582
rect 27950 44571 28258 44580
rect 28448 43852 28500 43858
rect 28448 43794 28500 43800
rect 27950 43548 28258 43557
rect 27950 43546 27956 43548
rect 28012 43546 28036 43548
rect 28092 43546 28116 43548
rect 28172 43546 28196 43548
rect 28252 43546 28258 43548
rect 28012 43494 28014 43546
rect 28194 43494 28196 43546
rect 27950 43492 27956 43494
rect 28012 43492 28036 43494
rect 28092 43492 28116 43494
rect 28172 43492 28196 43494
rect 28252 43492 28258 43494
rect 27950 43483 28258 43492
rect 28460 43110 28488 43794
rect 28448 43104 28500 43110
rect 28448 43046 28500 43052
rect 27950 42460 28258 42469
rect 27950 42458 27956 42460
rect 28012 42458 28036 42460
rect 28092 42458 28116 42460
rect 28172 42458 28196 42460
rect 28252 42458 28258 42460
rect 28012 42406 28014 42458
rect 28194 42406 28196 42458
rect 27950 42404 27956 42406
rect 28012 42404 28036 42406
rect 28092 42404 28116 42406
rect 28172 42404 28196 42406
rect 28252 42404 28258 42406
rect 27950 42395 28258 42404
rect 27950 41372 28258 41381
rect 27950 41370 27956 41372
rect 28012 41370 28036 41372
rect 28092 41370 28116 41372
rect 28172 41370 28196 41372
rect 28252 41370 28258 41372
rect 28012 41318 28014 41370
rect 28194 41318 28196 41370
rect 27950 41316 27956 41318
rect 28012 41316 28036 41318
rect 28092 41316 28116 41318
rect 28172 41316 28196 41318
rect 28252 41316 28258 41318
rect 27950 41307 28258 41316
rect 27804 41268 27856 41274
rect 27804 41210 27856 41216
rect 27712 40588 27764 40594
rect 27712 40530 27764 40536
rect 27724 38350 27752 40530
rect 27950 40284 28258 40293
rect 27950 40282 27956 40284
rect 28012 40282 28036 40284
rect 28092 40282 28116 40284
rect 28172 40282 28196 40284
rect 28252 40282 28258 40284
rect 28012 40230 28014 40282
rect 28194 40230 28196 40282
rect 27950 40228 27956 40230
rect 28012 40228 28036 40230
rect 28092 40228 28116 40230
rect 28172 40228 28196 40230
rect 28252 40228 28258 40230
rect 27950 40219 28258 40228
rect 28460 39982 28488 43046
rect 28448 39976 28500 39982
rect 28448 39918 28500 39924
rect 27804 39840 27856 39846
rect 27804 39782 27856 39788
rect 27816 38978 27844 39782
rect 28356 39500 28408 39506
rect 28356 39442 28408 39448
rect 27950 39196 28258 39205
rect 27950 39194 27956 39196
rect 28012 39194 28036 39196
rect 28092 39194 28116 39196
rect 28172 39194 28196 39196
rect 28252 39194 28258 39196
rect 28012 39142 28014 39194
rect 28194 39142 28196 39194
rect 27950 39140 27956 39142
rect 28012 39140 28036 39142
rect 28092 39140 28116 39142
rect 28172 39140 28196 39142
rect 28252 39140 28258 39142
rect 27950 39131 28258 39140
rect 27816 38950 28028 38978
rect 28368 38962 28396 39442
rect 28448 39432 28500 39438
rect 28448 39374 28500 39380
rect 28460 39030 28488 39374
rect 28448 39024 28500 39030
rect 28448 38966 28500 38972
rect 27896 38888 27948 38894
rect 27896 38830 27948 38836
rect 27712 38344 27764 38350
rect 27712 38286 27764 38292
rect 27620 37324 27672 37330
rect 27620 37266 27672 37272
rect 27724 37210 27752 38286
rect 27908 38196 27936 38830
rect 28000 38808 28028 38950
rect 28356 38956 28408 38962
rect 28356 38898 28408 38904
rect 28552 38842 28580 53926
rect 28724 43784 28776 43790
rect 28724 43726 28776 43732
rect 28736 43246 28764 43726
rect 28920 43654 28948 54266
rect 29104 53582 29132 56200
rect 29840 54194 29868 56200
rect 30576 54194 30604 56200
rect 31312 54194 31340 56200
rect 29828 54188 29880 54194
rect 29828 54130 29880 54136
rect 30564 54188 30616 54194
rect 30564 54130 30616 54136
rect 31300 54188 31352 54194
rect 31300 54130 31352 54136
rect 29644 54052 29696 54058
rect 29644 53994 29696 54000
rect 29092 53576 29144 53582
rect 29092 53518 29144 53524
rect 28908 43648 28960 43654
rect 28908 43590 28960 43596
rect 28724 43240 28776 43246
rect 28724 43182 28776 43188
rect 28736 42158 28764 43182
rect 28724 42152 28776 42158
rect 28724 42094 28776 42100
rect 28920 40594 28948 43590
rect 29184 43376 29236 43382
rect 29184 43318 29236 43324
rect 28908 40588 28960 40594
rect 28908 40530 28960 40536
rect 28908 40452 28960 40458
rect 28908 40394 28960 40400
rect 28724 39636 28776 39642
rect 28724 39578 28776 39584
rect 28632 39296 28684 39302
rect 28632 39238 28684 39244
rect 28080 38820 28132 38826
rect 28000 38780 28080 38808
rect 28080 38762 28132 38768
rect 28356 38820 28408 38826
rect 28356 38762 28408 38768
rect 28460 38814 28580 38842
rect 27816 38168 27936 38196
rect 27816 37806 27844 38168
rect 27950 38108 28258 38117
rect 27950 38106 27956 38108
rect 28012 38106 28036 38108
rect 28092 38106 28116 38108
rect 28172 38106 28196 38108
rect 28252 38106 28258 38108
rect 28012 38054 28014 38106
rect 28194 38054 28196 38106
rect 27950 38052 27956 38054
rect 28012 38052 28036 38054
rect 28092 38052 28116 38054
rect 28172 38052 28196 38054
rect 28252 38052 28258 38054
rect 27950 38043 28258 38052
rect 28172 37936 28224 37942
rect 28172 37878 28224 37884
rect 27804 37800 27856 37806
rect 27804 37742 27856 37748
rect 27816 37466 27844 37742
rect 27804 37460 27856 37466
rect 27804 37402 27856 37408
rect 28184 37262 28212 37878
rect 27632 37182 27752 37210
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 27528 36780 27580 36786
rect 27528 36722 27580 36728
rect 27540 36378 27568 36722
rect 27528 36372 27580 36378
rect 27528 36314 27580 36320
rect 27528 35284 27580 35290
rect 27448 35244 27528 35272
rect 27528 35226 27580 35232
rect 27540 34202 27568 35226
rect 27528 34196 27580 34202
rect 27528 34138 27580 34144
rect 27528 34060 27580 34066
rect 27528 34002 27580 34008
rect 27540 33946 27568 34002
rect 27172 31726 27292 31754
rect 27356 33918 27568 33946
rect 27172 31346 27200 31726
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27068 30796 27120 30802
rect 27068 30738 27120 30744
rect 27080 29646 27108 30738
rect 27068 29640 27120 29646
rect 27068 29582 27120 29588
rect 27080 29170 27108 29582
rect 27068 29164 27120 29170
rect 27068 29106 27120 29112
rect 27068 28484 27120 28490
rect 27068 28426 27120 28432
rect 26976 26784 27028 26790
rect 26976 26726 27028 26732
rect 26988 26382 27016 26726
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 26884 26240 26936 26246
rect 26884 26182 26936 26188
rect 26792 24404 26844 24410
rect 26792 24346 26844 24352
rect 26804 23866 26832 24346
rect 26792 23860 26844 23866
rect 26792 23802 26844 23808
rect 26528 23480 26740 23508
rect 26528 22506 26556 23480
rect 26896 22710 26924 26182
rect 26976 26036 27028 26042
rect 26976 25978 27028 25984
rect 26988 24886 27016 25978
rect 26976 24880 27028 24886
rect 26976 24822 27028 24828
rect 26988 23322 27016 24822
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 26884 22704 26936 22710
rect 26884 22646 26936 22652
rect 26516 22500 26568 22506
rect 26516 22442 26568 22448
rect 26344 22066 26464 22094
rect 26528 22094 26556 22442
rect 26608 22228 26660 22234
rect 26804 22222 26924 22250
rect 26804 22216 26832 22222
rect 26660 22188 26832 22216
rect 26608 22170 26660 22176
rect 26896 22166 26924 22222
rect 26884 22160 26936 22166
rect 26884 22102 26936 22108
rect 26528 22066 26740 22094
rect 26148 20596 26200 20602
rect 26148 20538 26200 20544
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 26160 18970 26188 20402
rect 26344 19174 26372 22066
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26148 18964 26200 18970
rect 26148 18906 26200 18912
rect 26436 18834 26464 21830
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26252 16640 26280 18702
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26344 17338 26372 18566
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 26252 16612 26372 16640
rect 26344 16454 26372 16612
rect 26332 16448 26384 16454
rect 26332 16390 26384 16396
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26160 15162 26188 15982
rect 26528 15706 26556 19654
rect 26620 19378 26648 20334
rect 26608 19372 26660 19378
rect 26608 19314 26660 19320
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26620 17066 26648 18770
rect 26608 17060 26660 17066
rect 26608 17002 26660 17008
rect 26620 16794 26648 17002
rect 26608 16788 26660 16794
rect 26608 16730 26660 16736
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26148 15156 26200 15162
rect 26148 15098 26200 15104
rect 26160 14346 26188 15098
rect 26620 14958 26648 16730
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 26712 12918 26740 22066
rect 26792 21956 26844 21962
rect 26792 21898 26844 21904
rect 26804 20058 26832 21898
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 27080 19990 27108 28426
rect 27172 27130 27200 31282
rect 27356 30666 27384 33918
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27436 33516 27488 33522
rect 27436 33458 27488 33464
rect 27344 30660 27396 30666
rect 27344 30602 27396 30608
rect 27356 29714 27384 30602
rect 27448 30122 27476 33458
rect 27540 33114 27568 33798
rect 27528 33108 27580 33114
rect 27528 33050 27580 33056
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27540 31822 27568 31962
rect 27528 31816 27580 31822
rect 27528 31758 27580 31764
rect 27540 31278 27568 31758
rect 27528 31272 27580 31278
rect 27528 31214 27580 31220
rect 27528 30184 27580 30190
rect 27528 30126 27580 30132
rect 27436 30116 27488 30122
rect 27436 30058 27488 30064
rect 27540 29714 27568 30126
rect 27344 29708 27396 29714
rect 27344 29650 27396 29656
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27632 28694 27660 37182
rect 27950 37020 28258 37029
rect 27950 37018 27956 37020
rect 28012 37018 28036 37020
rect 28092 37018 28116 37020
rect 28172 37018 28196 37020
rect 28252 37018 28258 37020
rect 28012 36966 28014 37018
rect 28194 36966 28196 37018
rect 27950 36964 27956 36966
rect 28012 36964 28036 36966
rect 28092 36964 28116 36966
rect 28172 36964 28196 36966
rect 28252 36964 28258 36966
rect 27950 36955 28258 36964
rect 28368 36904 28396 38762
rect 28276 36876 28396 36904
rect 28276 36174 28304 36876
rect 28356 36236 28408 36242
rect 28356 36178 28408 36184
rect 28264 36168 28316 36174
rect 28264 36110 28316 36116
rect 27950 35932 28258 35941
rect 27950 35930 27956 35932
rect 28012 35930 28036 35932
rect 28092 35930 28116 35932
rect 28172 35930 28196 35932
rect 28252 35930 28258 35932
rect 28012 35878 28014 35930
rect 28194 35878 28196 35930
rect 27950 35876 27956 35878
rect 28012 35876 28036 35878
rect 28092 35876 28116 35878
rect 28172 35876 28196 35878
rect 28252 35876 28258 35878
rect 27950 35867 28258 35876
rect 27710 35728 27766 35737
rect 27710 35663 27766 35672
rect 27724 35630 27752 35663
rect 27712 35624 27764 35630
rect 27712 35566 27764 35572
rect 27804 34944 27856 34950
rect 27804 34886 27856 34892
rect 27712 34400 27764 34406
rect 27712 34342 27764 34348
rect 27724 31906 27752 34342
rect 27816 32026 27844 34886
rect 27950 34844 28258 34853
rect 27950 34842 27956 34844
rect 28012 34842 28036 34844
rect 28092 34842 28116 34844
rect 28172 34842 28196 34844
rect 28252 34842 28258 34844
rect 28012 34790 28014 34842
rect 28194 34790 28196 34842
rect 27950 34788 27956 34790
rect 28012 34788 28036 34790
rect 28092 34788 28116 34790
rect 28172 34788 28196 34790
rect 28252 34788 28258 34790
rect 27950 34779 28258 34788
rect 28264 34740 28316 34746
rect 28264 34682 28316 34688
rect 28276 34649 28304 34682
rect 28262 34640 28318 34649
rect 28262 34575 28318 34584
rect 27950 33756 28258 33765
rect 27950 33754 27956 33756
rect 28012 33754 28036 33756
rect 28092 33754 28116 33756
rect 28172 33754 28196 33756
rect 28252 33754 28258 33756
rect 28012 33702 28014 33754
rect 28194 33702 28196 33754
rect 27950 33700 27956 33702
rect 28012 33700 28036 33702
rect 28092 33700 28116 33702
rect 28172 33700 28196 33702
rect 28252 33700 28258 33702
rect 27950 33691 28258 33700
rect 28368 33318 28396 36178
rect 28356 33312 28408 33318
rect 28356 33254 28408 33260
rect 28368 32978 28396 33254
rect 28356 32972 28408 32978
rect 28356 32914 28408 32920
rect 27950 32668 28258 32677
rect 27950 32666 27956 32668
rect 28012 32666 28036 32668
rect 28092 32666 28116 32668
rect 28172 32666 28196 32668
rect 28252 32666 28258 32668
rect 28012 32614 28014 32666
rect 28194 32614 28196 32666
rect 27950 32612 27956 32614
rect 28012 32612 28036 32614
rect 28092 32612 28116 32614
rect 28172 32612 28196 32614
rect 28252 32612 28258 32614
rect 27950 32603 28258 32612
rect 28460 32552 28488 38814
rect 28540 38752 28592 38758
rect 28540 38694 28592 38700
rect 28552 38418 28580 38694
rect 28644 38486 28672 39238
rect 28736 38894 28764 39578
rect 28816 39432 28868 39438
rect 28816 39374 28868 39380
rect 28724 38888 28776 38894
rect 28724 38830 28776 38836
rect 28632 38480 28684 38486
rect 28632 38422 28684 38428
rect 28540 38412 28592 38418
rect 28540 38354 28592 38360
rect 28540 38276 28592 38282
rect 28540 38218 28592 38224
rect 28552 37738 28580 38218
rect 28540 37732 28592 37738
rect 28540 37674 28592 37680
rect 28540 37324 28592 37330
rect 28540 37266 28592 37272
rect 28276 32524 28488 32552
rect 28276 32366 28304 32524
rect 27896 32360 27948 32366
rect 27896 32302 27948 32308
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 27804 32020 27856 32026
rect 27804 31962 27856 31968
rect 27908 31906 27936 32302
rect 28356 32292 28408 32298
rect 28356 32234 28408 32240
rect 27724 31878 27936 31906
rect 27712 31680 27764 31686
rect 27712 31622 27764 31628
rect 27620 28688 27672 28694
rect 27620 28630 27672 28636
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27632 28014 27660 28494
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27620 27396 27672 27402
rect 27620 27338 27672 27344
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 27160 27124 27212 27130
rect 27160 27066 27212 27072
rect 27160 26580 27212 26586
rect 27160 26522 27212 26528
rect 27172 26450 27200 26522
rect 27160 26444 27212 26450
rect 27160 26386 27212 26392
rect 27264 25430 27292 27270
rect 27436 25696 27488 25702
rect 27436 25638 27488 25644
rect 27252 25424 27304 25430
rect 27252 25366 27304 25372
rect 27448 24954 27476 25638
rect 27632 25242 27660 27338
rect 27540 25214 27660 25242
rect 27436 24948 27488 24954
rect 27436 24890 27488 24896
rect 27448 24342 27476 24890
rect 27540 24614 27568 25214
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 27632 24614 27660 25094
rect 27528 24608 27580 24614
rect 27528 24550 27580 24556
rect 27620 24608 27672 24614
rect 27620 24550 27672 24556
rect 27436 24336 27488 24342
rect 27436 24278 27488 24284
rect 27540 24274 27568 24550
rect 27528 24268 27580 24274
rect 27528 24210 27580 24216
rect 27540 23610 27568 24210
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27632 23798 27660 24006
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 27540 23582 27660 23610
rect 27632 23322 27660 23582
rect 27528 23316 27580 23322
rect 27528 23258 27580 23264
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 27540 23202 27568 23258
rect 27160 23180 27212 23186
rect 27540 23174 27660 23202
rect 27160 23122 27212 23128
rect 27172 22642 27200 23122
rect 27528 23044 27580 23050
rect 27528 22986 27580 22992
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27540 22574 27568 22986
rect 27528 22568 27580 22574
rect 27528 22510 27580 22516
rect 27160 20324 27212 20330
rect 27160 20266 27212 20272
rect 27068 19984 27120 19990
rect 27068 19926 27120 19932
rect 27172 19854 27200 20266
rect 27528 19916 27580 19922
rect 27528 19858 27580 19864
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27344 19780 27396 19786
rect 27344 19722 27396 19728
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26804 16658 26832 19314
rect 27264 19281 27292 19654
rect 27250 19272 27306 19281
rect 27250 19207 27306 19216
rect 27160 18692 27212 18698
rect 27160 18634 27212 18640
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 27172 16250 27200 18634
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 27264 18358 27292 18566
rect 27252 18352 27304 18358
rect 27252 18294 27304 18300
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 26884 16176 26936 16182
rect 26884 16118 26936 16124
rect 26896 15434 26924 16118
rect 26884 15428 26936 15434
rect 26884 15370 26936 15376
rect 26700 12912 26752 12918
rect 26700 12854 26752 12860
rect 27160 12708 27212 12714
rect 27160 12650 27212 12656
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26056 1692 26108 1698
rect 26056 1634 26108 1640
rect 26528 800 26556 2450
rect 27172 2446 27200 12650
rect 27264 3398 27292 18294
rect 27356 17882 27384 19722
rect 27436 19168 27488 19174
rect 27436 19110 27488 19116
rect 27344 17876 27396 17882
rect 27344 17818 27396 17824
rect 27448 17814 27476 19110
rect 27540 18222 27568 19858
rect 27632 18578 27660 23174
rect 27724 18737 27752 31622
rect 27950 31580 28258 31589
rect 27950 31578 27956 31580
rect 28012 31578 28036 31580
rect 28092 31578 28116 31580
rect 28172 31578 28196 31580
rect 28252 31578 28258 31580
rect 28012 31526 28014 31578
rect 28194 31526 28196 31578
rect 27950 31524 27956 31526
rect 28012 31524 28036 31526
rect 28092 31524 28116 31526
rect 28172 31524 28196 31526
rect 28252 31524 28258 31526
rect 27950 31515 28258 31524
rect 28368 30938 28396 32234
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 27950 30492 28258 30501
rect 27950 30490 27956 30492
rect 28012 30490 28036 30492
rect 28092 30490 28116 30492
rect 28172 30490 28196 30492
rect 28252 30490 28258 30492
rect 28012 30438 28014 30490
rect 28194 30438 28196 30490
rect 27950 30436 27956 30438
rect 28012 30436 28036 30438
rect 28092 30436 28116 30438
rect 28172 30436 28196 30438
rect 28252 30436 28258 30438
rect 27950 30427 28258 30436
rect 27950 29404 28258 29413
rect 27950 29402 27956 29404
rect 28012 29402 28036 29404
rect 28092 29402 28116 29404
rect 28172 29402 28196 29404
rect 28252 29402 28258 29404
rect 28012 29350 28014 29402
rect 28194 29350 28196 29402
rect 27950 29348 27956 29350
rect 28012 29348 28036 29350
rect 28092 29348 28116 29350
rect 28172 29348 28196 29350
rect 28252 29348 28258 29350
rect 27950 29339 28258 29348
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 27950 28316 28258 28325
rect 27950 28314 27956 28316
rect 28012 28314 28036 28316
rect 28092 28314 28116 28316
rect 28172 28314 28196 28316
rect 28252 28314 28258 28316
rect 28012 28262 28014 28314
rect 28194 28262 28196 28314
rect 27950 28260 27956 28262
rect 28012 28260 28036 28262
rect 28092 28260 28116 28262
rect 28172 28260 28196 28262
rect 28252 28260 28258 28262
rect 27950 28251 28258 28260
rect 27804 28144 27856 28150
rect 27804 28086 27856 28092
rect 27816 26586 27844 28086
rect 28368 27674 28396 28358
rect 28460 27962 28488 32302
rect 28552 29578 28580 37266
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 28644 35766 28672 37198
rect 28724 36780 28776 36786
rect 28724 36722 28776 36728
rect 28632 35760 28684 35766
rect 28632 35702 28684 35708
rect 28644 35086 28672 35702
rect 28632 35080 28684 35086
rect 28632 35022 28684 35028
rect 28632 34672 28684 34678
rect 28632 34614 28684 34620
rect 28644 30054 28672 34614
rect 28736 33658 28764 36722
rect 28828 36242 28856 39374
rect 28920 37806 28948 40394
rect 29000 39364 29052 39370
rect 29000 39306 29052 39312
rect 28908 37800 28960 37806
rect 28908 37742 28960 37748
rect 28816 36236 28868 36242
rect 28816 36178 28868 36184
rect 28908 35216 28960 35222
rect 28908 35158 28960 35164
rect 28816 35080 28868 35086
rect 28816 35022 28868 35028
rect 28828 33930 28856 35022
rect 28816 33924 28868 33930
rect 28816 33866 28868 33872
rect 28724 33652 28776 33658
rect 28724 33594 28776 33600
rect 28920 33114 28948 35158
rect 28908 33108 28960 33114
rect 28908 33050 28960 33056
rect 28724 32972 28776 32978
rect 28724 32914 28776 32920
rect 28736 31906 28764 32914
rect 29012 32774 29040 39306
rect 29092 38276 29144 38282
rect 29092 38218 29144 38224
rect 29104 34202 29132 38218
rect 29196 36650 29224 43318
rect 29368 42288 29420 42294
rect 29368 42230 29420 42236
rect 29276 37392 29328 37398
rect 29276 37334 29328 37340
rect 29184 36644 29236 36650
rect 29184 36586 29236 36592
rect 29184 35284 29236 35290
rect 29184 35226 29236 35232
rect 29196 34746 29224 35226
rect 29184 34740 29236 34746
rect 29184 34682 29236 34688
rect 29288 34406 29316 37334
rect 29380 36718 29408 42230
rect 29460 42016 29512 42022
rect 29460 41958 29512 41964
rect 29472 39370 29500 41958
rect 29460 39364 29512 39370
rect 29460 39306 29512 39312
rect 29368 36712 29420 36718
rect 29368 36654 29420 36660
rect 29460 36576 29512 36582
rect 29460 36518 29512 36524
rect 29472 36378 29500 36518
rect 29460 36372 29512 36378
rect 29460 36314 29512 36320
rect 29368 35624 29420 35630
rect 29368 35566 29420 35572
rect 29276 34400 29328 34406
rect 29276 34342 29328 34348
rect 29092 34196 29144 34202
rect 29092 34138 29144 34144
rect 29092 33992 29144 33998
rect 29092 33934 29144 33940
rect 29104 33658 29132 33934
rect 29092 33652 29144 33658
rect 29092 33594 29144 33600
rect 29184 33448 29236 33454
rect 29184 33390 29236 33396
rect 29000 32768 29052 32774
rect 29000 32710 29052 32716
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 28736 31890 29040 31906
rect 28736 31884 29052 31890
rect 28736 31878 29000 31884
rect 29000 31826 29052 31832
rect 29104 31770 29132 32370
rect 29196 32298 29224 33390
rect 29276 32972 29328 32978
rect 29276 32914 29328 32920
rect 29288 32366 29316 32914
rect 29276 32360 29328 32366
rect 29276 32302 29328 32308
rect 29184 32292 29236 32298
rect 29184 32234 29236 32240
rect 28920 31742 29132 31770
rect 28724 31680 28776 31686
rect 28722 31648 28724 31657
rect 28776 31648 28778 31657
rect 28722 31583 28778 31592
rect 28722 31512 28778 31521
rect 28920 31482 28948 31742
rect 28722 31447 28778 31456
rect 28908 31476 28960 31482
rect 28736 30841 28764 31447
rect 28908 31418 28960 31424
rect 28722 30832 28778 30841
rect 28722 30767 28778 30776
rect 28736 30258 28764 30767
rect 28816 30592 28868 30598
rect 28816 30534 28868 30540
rect 28908 30592 28960 30598
rect 28908 30534 28960 30540
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28632 30048 28684 30054
rect 28632 29990 28684 29996
rect 28828 29850 28856 30534
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 28540 29572 28592 29578
rect 28540 29514 28592 29520
rect 28724 29572 28776 29578
rect 28724 29514 28776 29520
rect 28540 28960 28592 28966
rect 28540 28902 28592 28908
rect 28552 28150 28580 28902
rect 28540 28144 28592 28150
rect 28540 28086 28592 28092
rect 28460 27934 28580 27962
rect 28448 27872 28500 27878
rect 28448 27814 28500 27820
rect 28356 27668 28408 27674
rect 28356 27610 28408 27616
rect 27950 27228 28258 27237
rect 27950 27226 27956 27228
rect 28012 27226 28036 27228
rect 28092 27226 28116 27228
rect 28172 27226 28196 27228
rect 28252 27226 28258 27228
rect 28012 27174 28014 27226
rect 28194 27174 28196 27226
rect 27950 27172 27956 27174
rect 28012 27172 28036 27174
rect 28092 27172 28116 27174
rect 28172 27172 28196 27174
rect 28252 27172 28258 27174
rect 27950 27163 28258 27172
rect 28172 26852 28224 26858
rect 28172 26794 28224 26800
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 28184 26382 28212 26794
rect 28172 26376 28224 26382
rect 28172 26318 28224 26324
rect 27804 26240 27856 26246
rect 27804 26182 27856 26188
rect 27816 22098 27844 26182
rect 27950 26140 28258 26149
rect 27950 26138 27956 26140
rect 28012 26138 28036 26140
rect 28092 26138 28116 26140
rect 28172 26138 28196 26140
rect 28252 26138 28258 26140
rect 28012 26086 28014 26138
rect 28194 26086 28196 26138
rect 27950 26084 27956 26086
rect 28012 26084 28036 26086
rect 28092 26084 28116 26086
rect 28172 26084 28196 26086
rect 28252 26084 28258 26086
rect 27950 26075 28258 26084
rect 27950 25052 28258 25061
rect 27950 25050 27956 25052
rect 28012 25050 28036 25052
rect 28092 25050 28116 25052
rect 28172 25050 28196 25052
rect 28252 25050 28258 25052
rect 28012 24998 28014 25050
rect 28194 24998 28196 25050
rect 27950 24996 27956 24998
rect 28012 24996 28036 24998
rect 28092 24996 28116 24998
rect 28172 24996 28196 24998
rect 28252 24996 28258 24998
rect 27950 24987 28258 24996
rect 27896 24880 27948 24886
rect 27894 24848 27896 24857
rect 27948 24848 27950 24857
rect 27894 24783 27950 24792
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 28092 24070 28120 24210
rect 28080 24064 28132 24070
rect 28080 24006 28132 24012
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27804 22092 27856 22098
rect 27804 22034 27856 22040
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27816 19854 27844 21286
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 27710 18728 27766 18737
rect 27816 18714 27844 19790
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 28368 19446 28396 27610
rect 28460 26926 28488 27814
rect 28552 27577 28580 27934
rect 28632 27872 28684 27878
rect 28632 27814 28684 27820
rect 28538 27568 28594 27577
rect 28538 27503 28594 27512
rect 28540 27328 28592 27334
rect 28540 27270 28592 27276
rect 28448 26920 28500 26926
rect 28448 26862 28500 26868
rect 28460 25838 28488 26862
rect 28448 25832 28500 25838
rect 28448 25774 28500 25780
rect 28460 24954 28488 25774
rect 28552 25702 28580 27270
rect 28540 25696 28592 25702
rect 28540 25638 28592 25644
rect 28448 24948 28500 24954
rect 28448 24890 28500 24896
rect 28538 24848 28594 24857
rect 28538 24783 28594 24792
rect 28448 24064 28500 24070
rect 28448 24006 28500 24012
rect 28460 22030 28488 24006
rect 28552 23118 28580 24783
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28552 22642 28580 23054
rect 28540 22636 28592 22642
rect 28540 22578 28592 22584
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 28644 21554 28672 27814
rect 28736 21894 28764 29514
rect 28828 29306 28856 29786
rect 28816 29300 28868 29306
rect 28816 29242 28868 29248
rect 28816 28688 28868 28694
rect 28816 28630 28868 28636
rect 28828 23497 28856 28630
rect 28920 26382 28948 30534
rect 29380 29714 29408 35566
rect 29656 35442 29684 53994
rect 30104 53984 30156 53990
rect 30104 53926 30156 53932
rect 30472 53984 30524 53990
rect 30472 53926 30524 53932
rect 29736 53440 29788 53446
rect 29736 53382 29788 53388
rect 29748 45490 29776 53382
rect 29736 45484 29788 45490
rect 29736 45426 29788 45432
rect 29736 42084 29788 42090
rect 29736 42026 29788 42032
rect 29748 41614 29776 42026
rect 29736 41608 29788 41614
rect 29736 41550 29788 41556
rect 29748 40526 29776 41550
rect 30116 41414 30144 53926
rect 30380 43376 30432 43382
rect 30380 43318 30432 43324
rect 30196 42356 30248 42362
rect 30392 42344 30420 43318
rect 30248 42316 30420 42344
rect 30196 42298 30248 42304
rect 30484 41414 30512 53926
rect 32048 53582 32076 56200
rect 32784 54262 32812 56200
rect 33520 54262 33548 56200
rect 32772 54256 32824 54262
rect 32772 54198 32824 54204
rect 33508 54256 33560 54262
rect 33508 54198 33560 54204
rect 34256 54194 34284 56200
rect 34244 54188 34296 54194
rect 34244 54130 34296 54136
rect 33416 54052 33468 54058
rect 33416 53994 33468 54000
rect 33968 54052 34020 54058
rect 33968 53994 34020 54000
rect 32950 53884 33258 53893
rect 32950 53882 32956 53884
rect 33012 53882 33036 53884
rect 33092 53882 33116 53884
rect 33172 53882 33196 53884
rect 33252 53882 33258 53884
rect 33012 53830 33014 53882
rect 33194 53830 33196 53882
rect 32950 53828 32956 53830
rect 33012 53828 33036 53830
rect 33092 53828 33116 53830
rect 33172 53828 33196 53830
rect 33252 53828 33258 53830
rect 32950 53819 33258 53828
rect 32036 53576 32088 53582
rect 32036 53518 32088 53524
rect 32128 53440 32180 53446
rect 32128 53382 32180 53388
rect 32140 45558 32168 53382
rect 32950 52796 33258 52805
rect 32950 52794 32956 52796
rect 33012 52794 33036 52796
rect 33092 52794 33116 52796
rect 33172 52794 33196 52796
rect 33252 52794 33258 52796
rect 33012 52742 33014 52794
rect 33194 52742 33196 52794
rect 32950 52740 32956 52742
rect 33012 52740 33036 52742
rect 33092 52740 33116 52742
rect 33172 52740 33196 52742
rect 33252 52740 33258 52742
rect 32950 52731 33258 52740
rect 32950 51708 33258 51717
rect 32950 51706 32956 51708
rect 33012 51706 33036 51708
rect 33092 51706 33116 51708
rect 33172 51706 33196 51708
rect 33252 51706 33258 51708
rect 33012 51654 33014 51706
rect 33194 51654 33196 51706
rect 32950 51652 32956 51654
rect 33012 51652 33036 51654
rect 33092 51652 33116 51654
rect 33172 51652 33196 51654
rect 33252 51652 33258 51654
rect 32950 51643 33258 51652
rect 32950 50620 33258 50629
rect 32950 50618 32956 50620
rect 33012 50618 33036 50620
rect 33092 50618 33116 50620
rect 33172 50618 33196 50620
rect 33252 50618 33258 50620
rect 33012 50566 33014 50618
rect 33194 50566 33196 50618
rect 32950 50564 32956 50566
rect 33012 50564 33036 50566
rect 33092 50564 33116 50566
rect 33172 50564 33196 50566
rect 33252 50564 33258 50566
rect 32950 50555 33258 50564
rect 32950 49532 33258 49541
rect 32950 49530 32956 49532
rect 33012 49530 33036 49532
rect 33092 49530 33116 49532
rect 33172 49530 33196 49532
rect 33252 49530 33258 49532
rect 33012 49478 33014 49530
rect 33194 49478 33196 49530
rect 32950 49476 32956 49478
rect 33012 49476 33036 49478
rect 33092 49476 33116 49478
rect 33172 49476 33196 49478
rect 33252 49476 33258 49478
rect 32950 49467 33258 49476
rect 32950 48444 33258 48453
rect 32950 48442 32956 48444
rect 33012 48442 33036 48444
rect 33092 48442 33116 48444
rect 33172 48442 33196 48444
rect 33252 48442 33258 48444
rect 33012 48390 33014 48442
rect 33194 48390 33196 48442
rect 32950 48388 32956 48390
rect 33012 48388 33036 48390
rect 33092 48388 33116 48390
rect 33172 48388 33196 48390
rect 33252 48388 33258 48390
rect 32950 48379 33258 48388
rect 32950 47356 33258 47365
rect 32950 47354 32956 47356
rect 33012 47354 33036 47356
rect 33092 47354 33116 47356
rect 33172 47354 33196 47356
rect 33252 47354 33258 47356
rect 33012 47302 33014 47354
rect 33194 47302 33196 47354
rect 32950 47300 32956 47302
rect 33012 47300 33036 47302
rect 33092 47300 33116 47302
rect 33172 47300 33196 47302
rect 33252 47300 33258 47302
rect 32950 47291 33258 47300
rect 32950 46268 33258 46277
rect 32950 46266 32956 46268
rect 33012 46266 33036 46268
rect 33092 46266 33116 46268
rect 33172 46266 33196 46268
rect 33252 46266 33258 46268
rect 33012 46214 33014 46266
rect 33194 46214 33196 46266
rect 32950 46212 32956 46214
rect 33012 46212 33036 46214
rect 33092 46212 33116 46214
rect 33172 46212 33196 46214
rect 33252 46212 33258 46214
rect 32950 46203 33258 46212
rect 32128 45552 32180 45558
rect 32128 45494 32180 45500
rect 33428 45490 33456 53994
rect 33416 45484 33468 45490
rect 33416 45426 33468 45432
rect 32864 45416 32916 45422
rect 32864 45358 32916 45364
rect 32680 45280 32732 45286
rect 32680 45222 32732 45228
rect 32588 43988 32640 43994
rect 32588 43930 32640 43936
rect 32220 43784 32272 43790
rect 32220 43726 32272 43732
rect 31300 43716 31352 43722
rect 31300 43658 31352 43664
rect 31312 43382 31340 43658
rect 31760 43648 31812 43654
rect 31760 43590 31812 43596
rect 31300 43376 31352 43382
rect 31300 43318 31352 43324
rect 31312 42294 31340 43318
rect 31772 42362 31800 43590
rect 32232 43314 32260 43726
rect 32220 43308 32272 43314
rect 32220 43250 32272 43256
rect 31944 43240 31996 43246
rect 31944 43182 31996 43188
rect 31760 42356 31812 42362
rect 31760 42298 31812 42304
rect 31300 42288 31352 42294
rect 31300 42230 31352 42236
rect 31208 41540 31260 41546
rect 31208 41482 31260 41488
rect 30116 41386 30236 41414
rect 30484 41386 30696 41414
rect 30012 41064 30064 41070
rect 30012 41006 30064 41012
rect 30024 40594 30052 41006
rect 30012 40588 30064 40594
rect 30012 40530 30064 40536
rect 29736 40520 29788 40526
rect 29736 40462 29788 40468
rect 29748 39846 29776 40462
rect 29736 39840 29788 39846
rect 29736 39782 29788 39788
rect 29828 39840 29880 39846
rect 29828 39782 29880 39788
rect 29748 38350 29776 39782
rect 29736 38344 29788 38350
rect 29736 38286 29788 38292
rect 29748 38010 29776 38286
rect 29736 38004 29788 38010
rect 29736 37946 29788 37952
rect 29840 37398 29868 39782
rect 29920 39024 29972 39030
rect 29920 38966 29972 38972
rect 29828 37392 29880 37398
rect 29828 37334 29880 37340
rect 29826 37224 29882 37233
rect 29826 37159 29882 37168
rect 29840 37126 29868 37159
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 29564 35414 29684 35442
rect 29460 30184 29512 30190
rect 29460 30126 29512 30132
rect 29368 29708 29420 29714
rect 29368 29650 29420 29656
rect 29472 29578 29500 30126
rect 29460 29572 29512 29578
rect 29460 29514 29512 29520
rect 29564 29170 29592 35414
rect 29932 34610 29960 38966
rect 30024 38282 30052 40530
rect 30104 39840 30156 39846
rect 30104 39782 30156 39788
rect 30116 39098 30144 39782
rect 30104 39092 30156 39098
rect 30104 39034 30156 39040
rect 30012 38276 30064 38282
rect 30012 38218 30064 38224
rect 30102 35592 30158 35601
rect 30102 35527 30158 35536
rect 30012 35148 30064 35154
rect 30012 35090 30064 35096
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 30024 34406 30052 35090
rect 30116 35086 30144 35527
rect 30104 35080 30156 35086
rect 30104 35022 30156 35028
rect 30012 34400 30064 34406
rect 30012 34342 30064 34348
rect 29644 33516 29696 33522
rect 29644 33458 29696 33464
rect 29276 29164 29328 29170
rect 29276 29106 29328 29112
rect 29552 29164 29604 29170
rect 29552 29106 29604 29112
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 28908 26376 28960 26382
rect 28908 26318 28960 26324
rect 29012 25294 29040 28970
rect 29092 26376 29144 26382
rect 29092 26318 29144 26324
rect 29104 26042 29132 26318
rect 29092 26036 29144 26042
rect 29092 25978 29144 25984
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 29092 25288 29144 25294
rect 29092 25230 29144 25236
rect 29104 24138 29132 25230
rect 29184 25220 29236 25226
rect 29184 25162 29236 25168
rect 29196 24750 29224 25162
rect 29184 24744 29236 24750
rect 29184 24686 29236 24692
rect 29288 24562 29316 29106
rect 29460 28960 29512 28966
rect 29460 28902 29512 28908
rect 29472 28626 29500 28902
rect 29460 28620 29512 28626
rect 29460 28562 29512 28568
rect 29552 28076 29604 28082
rect 29552 28018 29604 28024
rect 29564 27606 29592 28018
rect 29552 27600 29604 27606
rect 29552 27542 29604 27548
rect 29368 26444 29420 26450
rect 29368 26386 29420 26392
rect 29196 24534 29316 24562
rect 29092 24132 29144 24138
rect 29092 24074 29144 24080
rect 28814 23488 28870 23497
rect 28814 23423 28870 23432
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 28828 22710 28856 23054
rect 28816 22704 28868 22710
rect 28816 22646 28868 22652
rect 29196 22094 29224 24534
rect 29276 22976 29328 22982
rect 29380 22964 29408 26386
rect 29328 22936 29408 22964
rect 29276 22918 29328 22924
rect 29012 22066 29224 22094
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28356 19440 28408 19446
rect 28356 19382 28408 19388
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27908 18834 27936 19246
rect 27896 18828 27948 18834
rect 27896 18770 27948 18776
rect 27816 18686 28396 18714
rect 27710 18663 27766 18672
rect 27632 18550 27844 18578
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27528 18216 27580 18222
rect 27528 18158 27580 18164
rect 27436 17808 27488 17814
rect 27356 17756 27436 17762
rect 27356 17750 27488 17756
rect 27356 17734 27476 17750
rect 27540 17746 27568 18158
rect 27528 17740 27580 17746
rect 27356 15570 27384 17734
rect 27528 17682 27580 17688
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27448 16250 27476 16730
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27344 15564 27396 15570
rect 27344 15506 27396 15512
rect 27448 15434 27476 16186
rect 27540 16046 27568 17682
rect 27632 17678 27660 18226
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27712 17128 27764 17134
rect 27710 17096 27712 17105
rect 27764 17096 27766 17105
rect 27710 17031 27766 17040
rect 27816 16130 27844 18550
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27896 18080 27948 18086
rect 27894 18048 27896 18057
rect 27948 18048 27950 18057
rect 27894 17983 27950 17992
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 28368 17218 28396 18686
rect 28460 18426 28488 19314
rect 28736 18986 28764 21830
rect 28816 19304 28868 19310
rect 28816 19246 28868 19252
rect 28552 18958 28764 18986
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 28460 17678 28488 18362
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28276 17190 28396 17218
rect 28172 17128 28224 17134
rect 28172 17070 28224 17076
rect 28184 16658 28212 17070
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28276 16454 28304 17190
rect 28356 17128 28408 17134
rect 28356 17070 28408 17076
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28368 16250 28396 17070
rect 28448 16992 28500 16998
rect 28448 16934 28500 16940
rect 28460 16590 28488 16934
rect 28448 16584 28500 16590
rect 28448 16526 28500 16532
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 28356 16244 28408 16250
rect 28356 16186 28408 16192
rect 27816 16102 27936 16130
rect 27528 16040 27580 16046
rect 27804 16040 27856 16046
rect 27528 15982 27580 15988
rect 27724 15988 27804 15994
rect 27724 15982 27856 15988
rect 27724 15966 27844 15982
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27252 3392 27304 3398
rect 27252 3334 27304 3340
rect 27356 3058 27384 15302
rect 27448 3126 27476 15370
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27632 13530 27660 14962
rect 27724 14958 27752 15966
rect 27908 15858 27936 16102
rect 27816 15830 27936 15858
rect 28264 15904 28316 15910
rect 28264 15846 28316 15852
rect 27712 14952 27764 14958
rect 27712 14894 27764 14900
rect 27724 14482 27752 14894
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27816 12918 27844 15830
rect 27986 15600 28042 15609
rect 27986 15535 27988 15544
rect 28040 15535 28042 15544
rect 27988 15506 28040 15512
rect 28276 15434 28304 15846
rect 28264 15428 28316 15434
rect 28264 15370 28316 15376
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27988 14952 28040 14958
rect 27988 14894 28040 14900
rect 28000 14550 28028 14894
rect 27988 14544 28040 14550
rect 27988 14486 28040 14492
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27804 12912 27856 12918
rect 27804 12854 27856 12860
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27436 3120 27488 3126
rect 27436 3062 27488 3068
rect 27344 3052 27396 3058
rect 27344 2994 27396 3000
rect 27252 2984 27304 2990
rect 27252 2926 27304 2932
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 27264 800 27292 2926
rect 27816 2582 27844 12718
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28368 3194 28396 16186
rect 28460 10062 28488 16390
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28356 3188 28408 3194
rect 28356 3130 28408 3136
rect 27804 2576 27856 2582
rect 27804 2518 27856 2524
rect 28356 2508 28408 2514
rect 28356 2450 28408 2456
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28000 870 28120 898
rect 28000 800 28028 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8850 0 8906 800
rect 9586 0 9642 800
rect 10322 0 10378 800
rect 11058 0 11114 800
rect 11794 0 11850 800
rect 12530 0 12586 800
rect 13266 0 13322 800
rect 14002 0 14058 800
rect 14738 0 14794 800
rect 15474 0 15530 800
rect 16210 0 16266 800
rect 16946 0 17002 800
rect 17682 0 17738 800
rect 18418 0 18474 800
rect 19154 0 19210 800
rect 19890 0 19946 800
rect 20626 0 20682 800
rect 21362 0 21418 800
rect 22098 0 22154 800
rect 22834 0 22890 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25042 0 25098 800
rect 25778 0 25834 800
rect 26514 0 26570 800
rect 27250 0 27306 800
rect 27986 0 28042 800
rect 28092 762 28120 870
rect 28368 762 28396 2450
rect 28552 1970 28580 18958
rect 28722 18864 28778 18873
rect 28632 18828 28684 18834
rect 28722 18799 28724 18808
rect 28632 18770 28684 18776
rect 28776 18799 28778 18808
rect 28724 18770 28776 18776
rect 28644 18714 28672 18770
rect 28644 18686 28764 18714
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28644 12782 28672 17614
rect 28736 17202 28764 18686
rect 28724 17196 28776 17202
rect 28724 17138 28776 17144
rect 28724 16516 28776 16522
rect 28724 16458 28776 16464
rect 28736 12986 28764 16458
rect 28828 16454 28856 19246
rect 28908 18828 28960 18834
rect 28908 18770 28960 18776
rect 28920 17814 28948 18770
rect 29012 18748 29040 22066
rect 29012 18720 29224 18748
rect 28908 17808 28960 17814
rect 28908 17750 28960 17756
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 28816 16448 28868 16454
rect 28816 16390 28868 16396
rect 28828 16046 28856 16390
rect 28816 16040 28868 16046
rect 28816 15982 28868 15988
rect 28816 15700 28868 15706
rect 28816 15642 28868 15648
rect 28828 15609 28856 15642
rect 28814 15600 28870 15609
rect 28814 15535 28870 15544
rect 28816 15428 28868 15434
rect 28816 15370 28868 15376
rect 28828 14278 28856 15370
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28920 13462 28948 16594
rect 29196 15434 29224 18720
rect 29184 15428 29236 15434
rect 29184 15370 29236 15376
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 28908 13456 28960 13462
rect 28908 13398 28960 13404
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28724 12980 28776 12986
rect 28920 12968 28948 13262
rect 28724 12922 28776 12928
rect 28828 12940 28948 12968
rect 28632 12776 28684 12782
rect 28632 12718 28684 12724
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 28540 1964 28592 1970
rect 28540 1906 28592 1912
rect 28736 800 28764 2926
rect 28828 1902 28856 12940
rect 28906 12880 28962 12889
rect 28906 12815 28962 12824
rect 28920 12238 28948 12815
rect 29012 12714 29040 15098
rect 29092 15020 29144 15026
rect 29092 14962 29144 14968
rect 29104 14346 29132 14962
rect 29092 14340 29144 14346
rect 29092 14282 29144 14288
rect 29288 14006 29316 22918
rect 29368 17536 29420 17542
rect 29368 17478 29420 17484
rect 29380 16182 29408 17478
rect 29552 17196 29604 17202
rect 29552 17138 29604 17144
rect 29368 16176 29420 16182
rect 29368 16118 29420 16124
rect 29276 14000 29328 14006
rect 29276 13942 29328 13948
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 29000 12708 29052 12714
rect 29000 12650 29052 12656
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 29184 12164 29236 12170
rect 29184 12106 29236 12112
rect 29196 3058 29224 12106
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 28816 1896 28868 1902
rect 28816 1838 28868 1844
rect 29288 1834 29316 12922
rect 29380 7410 29408 16118
rect 29460 16040 29512 16046
rect 29460 15982 29512 15988
rect 29472 15706 29500 15982
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29472 15162 29500 15642
rect 29460 15156 29512 15162
rect 29460 15098 29512 15104
rect 29564 12782 29592 17138
rect 29656 15910 29684 33458
rect 29920 33312 29972 33318
rect 29920 33254 29972 33260
rect 29932 29510 29960 33254
rect 30012 30320 30064 30326
rect 30012 30262 30064 30268
rect 30024 29646 30052 30262
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 29920 29504 29972 29510
rect 29920 29446 29972 29452
rect 30104 29300 30156 29306
rect 30104 29242 30156 29248
rect 29736 29232 29788 29238
rect 29736 29174 29788 29180
rect 29748 28150 29776 29174
rect 30010 29064 30066 29073
rect 30010 28999 30066 29008
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 29736 28144 29788 28150
rect 29736 28086 29788 28092
rect 29736 28008 29788 28014
rect 29736 27950 29788 27956
rect 29748 19378 29776 27950
rect 29828 27872 29880 27878
rect 29828 27814 29880 27820
rect 29840 26926 29868 27814
rect 29932 27470 29960 28494
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 29828 26920 29880 26926
rect 29828 26862 29880 26868
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 29932 25344 29960 25638
rect 30024 25498 30052 28999
rect 30116 26790 30144 29242
rect 30208 28490 30236 41386
rect 30380 40928 30432 40934
rect 30380 40870 30432 40876
rect 30392 39914 30420 40870
rect 30668 40497 30696 41386
rect 30748 41200 30800 41206
rect 30748 41142 30800 41148
rect 30654 40488 30710 40497
rect 30472 40452 30524 40458
rect 30654 40423 30710 40432
rect 30472 40394 30524 40400
rect 30484 40186 30512 40394
rect 30472 40180 30524 40186
rect 30472 40122 30524 40128
rect 30380 39908 30432 39914
rect 30380 39850 30432 39856
rect 30484 39522 30512 40122
rect 30484 39494 30604 39522
rect 30576 39370 30604 39494
rect 30472 39364 30524 39370
rect 30472 39306 30524 39312
rect 30564 39364 30616 39370
rect 30564 39306 30616 39312
rect 30484 39098 30512 39306
rect 30668 39250 30696 40423
rect 30576 39222 30696 39250
rect 30472 39092 30524 39098
rect 30472 39034 30524 39040
rect 30472 38276 30524 38282
rect 30392 38236 30472 38264
rect 30392 35766 30420 38236
rect 30472 38218 30524 38224
rect 30472 36848 30524 36854
rect 30472 36790 30524 36796
rect 30484 36242 30512 36790
rect 30472 36236 30524 36242
rect 30472 36178 30524 36184
rect 30576 36122 30604 39222
rect 30656 37936 30708 37942
rect 30656 37878 30708 37884
rect 30668 37466 30696 37878
rect 30656 37460 30708 37466
rect 30656 37402 30708 37408
rect 30484 36094 30604 36122
rect 30380 35760 30432 35766
rect 30380 35702 30432 35708
rect 30288 35148 30340 35154
rect 30288 35090 30340 35096
rect 30300 31754 30328 35090
rect 30392 34921 30420 35702
rect 30378 34912 30434 34921
rect 30378 34847 30434 34856
rect 30392 34678 30420 34847
rect 30380 34672 30432 34678
rect 30380 34614 30432 34620
rect 30380 34060 30432 34066
rect 30380 34002 30432 34008
rect 30392 33590 30420 34002
rect 30380 33584 30432 33590
rect 30380 33526 30432 33532
rect 30380 32972 30432 32978
rect 30380 32914 30432 32920
rect 30392 32434 30420 32914
rect 30380 32428 30432 32434
rect 30380 32370 30432 32376
rect 30484 31754 30512 36094
rect 30564 35012 30616 35018
rect 30564 34954 30616 34960
rect 30576 33386 30604 34954
rect 30564 33380 30616 33386
rect 30564 33322 30616 33328
rect 30288 31748 30340 31754
rect 30288 31690 30340 31696
rect 30380 31748 30432 31754
rect 30484 31726 30604 31754
rect 30380 31690 30432 31696
rect 30300 30954 30328 31690
rect 30392 31142 30420 31690
rect 30380 31136 30432 31142
rect 30380 31078 30432 31084
rect 30300 30926 30512 30954
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30196 28484 30248 28490
rect 30196 28426 30248 28432
rect 30300 28218 30328 30738
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30288 28212 30340 28218
rect 30288 28154 30340 28160
rect 30196 28144 30248 28150
rect 30196 28086 30248 28092
rect 30208 27418 30236 28086
rect 30288 27532 30340 27538
rect 30392 27520 30420 30670
rect 30484 30394 30512 30926
rect 30472 30388 30524 30394
rect 30472 30330 30524 30336
rect 30472 30252 30524 30258
rect 30472 30194 30524 30200
rect 30484 29850 30512 30194
rect 30472 29844 30524 29850
rect 30472 29786 30524 29792
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30484 29306 30512 29650
rect 30472 29300 30524 29306
rect 30472 29242 30524 29248
rect 30472 29096 30524 29102
rect 30470 29064 30472 29073
rect 30524 29064 30526 29073
rect 30470 28999 30526 29008
rect 30340 27492 30420 27520
rect 30288 27474 30340 27480
rect 30208 27390 30328 27418
rect 30196 27328 30248 27334
rect 30196 27270 30248 27276
rect 30104 26784 30156 26790
rect 30104 26726 30156 26732
rect 30116 25838 30144 26726
rect 30104 25832 30156 25838
rect 30104 25774 30156 25780
rect 30012 25492 30064 25498
rect 30012 25434 30064 25440
rect 30012 25356 30064 25362
rect 29932 25316 30012 25344
rect 29932 24886 29960 25316
rect 30012 25298 30064 25304
rect 29920 24880 29972 24886
rect 29920 24822 29972 24828
rect 30208 24274 30236 27270
rect 30300 26994 30328 27390
rect 30288 26988 30340 26994
rect 30288 26930 30340 26936
rect 30300 25974 30328 26930
rect 30576 26874 30604 31726
rect 30668 27674 30696 37402
rect 30760 37126 30788 41142
rect 30840 41132 30892 41138
rect 30840 41074 30892 41080
rect 30852 39642 30880 41074
rect 31024 40724 31076 40730
rect 30944 40684 31024 40712
rect 30840 39636 30892 39642
rect 30840 39578 30892 39584
rect 30838 37904 30894 37913
rect 30838 37839 30894 37848
rect 30852 37806 30880 37839
rect 30840 37800 30892 37806
rect 30840 37742 30892 37748
rect 30748 37120 30800 37126
rect 30748 37062 30800 37068
rect 30748 35760 30800 35766
rect 30748 35702 30800 35708
rect 30760 35290 30788 35702
rect 30748 35284 30800 35290
rect 30748 35226 30800 35232
rect 30746 35184 30802 35193
rect 30746 35119 30802 35128
rect 30760 28014 30788 35119
rect 30944 34474 30972 40684
rect 31024 40666 31076 40672
rect 31116 39296 31168 39302
rect 31116 39238 31168 39244
rect 31024 38480 31076 38486
rect 31024 38422 31076 38428
rect 31036 37874 31064 38422
rect 31024 37868 31076 37874
rect 31024 37810 31076 37816
rect 31128 37210 31156 39238
rect 31220 37330 31248 41482
rect 31312 41002 31340 42230
rect 31956 42022 31984 43182
rect 31944 42016 31996 42022
rect 31944 41958 31996 41964
rect 31668 41676 31720 41682
rect 31668 41618 31720 41624
rect 31680 41546 31708 41618
rect 31668 41540 31720 41546
rect 31668 41482 31720 41488
rect 31956 41414 31984 41958
rect 32600 41414 32628 43930
rect 31956 41386 32076 41414
rect 31300 40996 31352 41002
rect 31300 40938 31352 40944
rect 31312 40186 31340 40938
rect 31484 40384 31536 40390
rect 31484 40326 31536 40332
rect 31300 40180 31352 40186
rect 31300 40122 31352 40128
rect 31496 39574 31524 40326
rect 31484 39568 31536 39574
rect 31484 39510 31536 39516
rect 31300 37664 31352 37670
rect 31300 37606 31352 37612
rect 31208 37324 31260 37330
rect 31208 37266 31260 37272
rect 31312 37262 31340 37606
rect 31496 37330 31524 39510
rect 31944 38820 31996 38826
rect 31944 38762 31996 38768
rect 31576 38548 31628 38554
rect 31628 38508 31800 38536
rect 31576 38490 31628 38496
rect 31668 38344 31720 38350
rect 31668 38286 31720 38292
rect 31576 38276 31628 38282
rect 31576 38218 31628 38224
rect 31484 37324 31536 37330
rect 31484 37266 31536 37272
rect 31300 37256 31352 37262
rect 31128 37182 31248 37210
rect 31300 37198 31352 37204
rect 31116 37120 31168 37126
rect 31116 37062 31168 37068
rect 31024 34944 31076 34950
rect 31024 34886 31076 34892
rect 30932 34468 30984 34474
rect 30932 34410 30984 34416
rect 31036 32994 31064 34886
rect 30944 32966 31064 32994
rect 30944 32774 30972 32966
rect 31024 32904 31076 32910
rect 31024 32846 31076 32852
rect 30932 32768 30984 32774
rect 30932 32710 30984 32716
rect 31036 31249 31064 32846
rect 31128 32502 31156 37062
rect 31220 35154 31248 37182
rect 31588 35698 31616 38218
rect 31680 37942 31708 38286
rect 31668 37936 31720 37942
rect 31668 37878 31720 37884
rect 31680 37466 31708 37878
rect 31772 37738 31800 38508
rect 31956 38282 31984 38762
rect 32048 38282 32076 41386
rect 32508 41386 32628 41414
rect 32312 41064 32364 41070
rect 32312 41006 32364 41012
rect 32324 39982 32352 41006
rect 32312 39976 32364 39982
rect 32312 39918 32364 39924
rect 31944 38276 31996 38282
rect 31944 38218 31996 38224
rect 32036 38276 32088 38282
rect 32036 38218 32088 38224
rect 32220 38208 32272 38214
rect 32220 38150 32272 38156
rect 31760 37732 31812 37738
rect 31760 37674 31812 37680
rect 31668 37460 31720 37466
rect 31668 37402 31720 37408
rect 32128 37120 32180 37126
rect 32128 37062 32180 37068
rect 32036 36916 32088 36922
rect 32036 36858 32088 36864
rect 31668 36712 31720 36718
rect 31668 36654 31720 36660
rect 31680 36224 31708 36654
rect 32048 36378 32076 36858
rect 32036 36372 32088 36378
rect 32036 36314 32088 36320
rect 31852 36304 31904 36310
rect 31850 36272 31852 36281
rect 31904 36272 31906 36281
rect 31760 36236 31812 36242
rect 31680 36196 31760 36224
rect 31850 36207 31906 36216
rect 31760 36178 31812 36184
rect 31576 35692 31628 35698
rect 31576 35634 31628 35640
rect 31298 35184 31354 35193
rect 31208 35148 31260 35154
rect 31298 35119 31354 35128
rect 31208 35090 31260 35096
rect 31206 35048 31262 35057
rect 31206 34983 31262 34992
rect 31220 34950 31248 34983
rect 31208 34944 31260 34950
rect 31208 34886 31260 34892
rect 31312 34746 31340 35119
rect 31392 35080 31444 35086
rect 31390 35048 31392 35057
rect 31444 35048 31446 35057
rect 31390 34983 31446 34992
rect 31300 34740 31352 34746
rect 31300 34682 31352 34688
rect 31484 34400 31536 34406
rect 31484 34342 31536 34348
rect 31208 33856 31260 33862
rect 31208 33798 31260 33804
rect 31116 32496 31168 32502
rect 31116 32438 31168 32444
rect 31022 31240 31078 31249
rect 31022 31175 31078 31184
rect 31220 29209 31248 33798
rect 31496 32978 31524 34342
rect 31588 33318 31616 35634
rect 31760 35488 31812 35494
rect 31760 35430 31812 35436
rect 31668 35148 31720 35154
rect 31668 35090 31720 35096
rect 31576 33312 31628 33318
rect 31576 33254 31628 33260
rect 31484 32972 31536 32978
rect 31484 32914 31536 32920
rect 31300 32768 31352 32774
rect 31300 32710 31352 32716
rect 31312 32570 31340 32710
rect 31300 32564 31352 32570
rect 31300 32506 31352 32512
rect 31576 32564 31628 32570
rect 31576 32506 31628 32512
rect 31300 30728 31352 30734
rect 31300 30670 31352 30676
rect 31312 30326 31340 30670
rect 31588 30666 31616 32506
rect 31680 31822 31708 35090
rect 31772 34746 31800 35430
rect 31760 34740 31812 34746
rect 31760 34682 31812 34688
rect 31852 33108 31904 33114
rect 31852 33050 31904 33056
rect 31668 31816 31720 31822
rect 31668 31758 31720 31764
rect 31680 31278 31708 31758
rect 31668 31272 31720 31278
rect 31668 31214 31720 31220
rect 31576 30660 31628 30666
rect 31576 30602 31628 30608
rect 31300 30320 31352 30326
rect 31300 30262 31352 30268
rect 31206 29200 31262 29209
rect 31206 29135 31262 29144
rect 31116 28416 31168 28422
rect 31116 28358 31168 28364
rect 31300 28416 31352 28422
rect 31300 28358 31352 28364
rect 30748 28008 30800 28014
rect 30748 27950 30800 27956
rect 30760 27674 30788 27950
rect 30656 27668 30708 27674
rect 30656 27610 30708 27616
rect 30748 27668 30800 27674
rect 30748 27610 30800 27616
rect 31022 27568 31078 27577
rect 31022 27503 31078 27512
rect 30656 27328 30708 27334
rect 30656 27270 30708 27276
rect 30748 27328 30800 27334
rect 30748 27270 30800 27276
rect 30668 27130 30696 27270
rect 30656 27124 30708 27130
rect 30656 27066 30708 27072
rect 30760 26874 30788 27270
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30576 26846 30788 26874
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30288 25968 30340 25974
rect 30288 25910 30340 25916
rect 30300 24954 30328 25910
rect 30288 24948 30340 24954
rect 30288 24890 30340 24896
rect 30288 24608 30340 24614
rect 30288 24550 30340 24556
rect 30300 24274 30328 24550
rect 30196 24268 30248 24274
rect 30196 24210 30248 24216
rect 30288 24268 30340 24274
rect 30288 24210 30340 24216
rect 30196 24064 30248 24070
rect 30196 24006 30248 24012
rect 30102 23488 30158 23497
rect 30102 23423 30158 23432
rect 29828 23180 29880 23186
rect 29828 23122 29880 23128
rect 29840 21486 29868 23122
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 29932 21690 29960 21966
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 29828 21480 29880 21486
rect 29828 21422 29880 21428
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 29840 19310 29868 21422
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29736 17740 29788 17746
rect 29736 17682 29788 17688
rect 29748 17134 29776 17682
rect 29736 17128 29788 17134
rect 29736 17070 29788 17076
rect 29748 16454 29776 17070
rect 29736 16448 29788 16454
rect 29736 16390 29788 16396
rect 29644 15904 29696 15910
rect 29644 15846 29696 15852
rect 29644 15632 29696 15638
rect 29644 15574 29696 15580
rect 29656 15162 29684 15574
rect 29748 15570 29776 16390
rect 29736 15564 29788 15570
rect 29736 15506 29788 15512
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 30116 15094 30144 23423
rect 30208 21622 30236 24006
rect 30392 22778 30420 26726
rect 30760 26450 30788 26846
rect 30748 26444 30800 26450
rect 30748 26386 30800 26392
rect 30564 25900 30616 25906
rect 30564 25842 30616 25848
rect 30472 24200 30524 24206
rect 30472 24142 30524 24148
rect 30484 23866 30512 24142
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 30576 23798 30604 25842
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 30380 22772 30432 22778
rect 30380 22714 30432 22720
rect 30472 22704 30524 22710
rect 30470 22672 30472 22681
rect 30524 22672 30526 22681
rect 30380 22636 30432 22642
rect 30470 22607 30526 22616
rect 30380 22578 30432 22584
rect 30392 22166 30420 22578
rect 30380 22160 30432 22166
rect 30380 22102 30432 22108
rect 30668 22094 30696 25094
rect 30484 22066 30696 22094
rect 30484 21690 30512 22066
rect 30472 21684 30524 21690
rect 30472 21626 30524 21632
rect 30196 21616 30248 21622
rect 30196 21558 30248 21564
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30668 20942 30696 21286
rect 30656 20936 30708 20942
rect 30656 20878 30708 20884
rect 30748 20936 30800 20942
rect 30748 20878 30800 20884
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 30196 18148 30248 18154
rect 30196 18090 30248 18096
rect 30208 17746 30236 18090
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 30300 17610 30328 20742
rect 30470 20632 30526 20641
rect 30470 20567 30472 20576
rect 30524 20567 30526 20576
rect 30472 20538 30524 20544
rect 30760 20534 30788 20878
rect 30748 20528 30800 20534
rect 30748 20470 30800 20476
rect 30852 18358 30880 27066
rect 31036 26926 31064 27503
rect 31024 26920 31076 26926
rect 31024 26862 31076 26868
rect 31036 26382 31064 26862
rect 31128 26432 31156 28358
rect 31206 27160 31262 27169
rect 31206 27095 31208 27104
rect 31260 27095 31262 27104
rect 31208 27066 31260 27072
rect 31312 26994 31340 28358
rect 31484 27396 31536 27402
rect 31484 27338 31536 27344
rect 31300 26988 31352 26994
rect 31300 26930 31352 26936
rect 31312 26897 31340 26930
rect 31392 26920 31444 26926
rect 31298 26888 31354 26897
rect 31392 26862 31444 26868
rect 31298 26823 31354 26832
rect 31300 26784 31352 26790
rect 31300 26726 31352 26732
rect 31312 26450 31340 26726
rect 31208 26444 31260 26450
rect 31128 26404 31208 26432
rect 31208 26386 31260 26392
rect 31300 26444 31352 26450
rect 31300 26386 31352 26392
rect 31024 26376 31076 26382
rect 31024 26318 31076 26324
rect 31024 25696 31076 25702
rect 31024 25638 31076 25644
rect 31036 24954 31064 25638
rect 31404 25242 31432 26862
rect 31496 26858 31524 27338
rect 31760 27328 31812 27334
rect 31760 27270 31812 27276
rect 31484 26852 31536 26858
rect 31484 26794 31536 26800
rect 31312 25214 31432 25242
rect 31116 25152 31168 25158
rect 31116 25094 31168 25100
rect 31024 24948 31076 24954
rect 31024 24890 31076 24896
rect 31128 22098 31156 25094
rect 31312 24750 31340 25214
rect 31392 25152 31444 25158
rect 31392 25094 31444 25100
rect 31300 24744 31352 24750
rect 31300 24686 31352 24692
rect 31208 24608 31260 24614
rect 31208 24550 31260 24556
rect 31220 24342 31248 24550
rect 31208 24336 31260 24342
rect 31208 24278 31260 24284
rect 31312 22438 31340 24686
rect 31300 22432 31352 22438
rect 31300 22374 31352 22380
rect 31116 22092 31168 22098
rect 31116 22034 31168 22040
rect 31404 20806 31432 25094
rect 31392 20800 31444 20806
rect 31392 20742 31444 20748
rect 31298 19272 31354 19281
rect 31298 19207 31354 19216
rect 31312 18766 31340 19207
rect 31496 18834 31524 26794
rect 31772 25362 31800 27270
rect 31864 27130 31892 33050
rect 32140 32910 32168 37062
rect 32232 36786 32260 38150
rect 32324 37874 32352 39918
rect 32404 38752 32456 38758
rect 32404 38694 32456 38700
rect 32312 37868 32364 37874
rect 32312 37810 32364 37816
rect 32416 36922 32444 38694
rect 32508 37262 32536 41386
rect 32588 40928 32640 40934
rect 32588 40870 32640 40876
rect 32600 40474 32628 40870
rect 32692 40594 32720 45222
rect 32876 43858 32904 45358
rect 32950 45180 33258 45189
rect 32950 45178 32956 45180
rect 33012 45178 33036 45180
rect 33092 45178 33116 45180
rect 33172 45178 33196 45180
rect 33252 45178 33258 45180
rect 33012 45126 33014 45178
rect 33194 45126 33196 45178
rect 32950 45124 32956 45126
rect 33012 45124 33036 45126
rect 33092 45124 33116 45126
rect 33172 45124 33196 45126
rect 33252 45124 33258 45126
rect 32950 45115 33258 45124
rect 32950 44092 33258 44101
rect 32950 44090 32956 44092
rect 33012 44090 33036 44092
rect 33092 44090 33116 44092
rect 33172 44090 33196 44092
rect 33252 44090 33258 44092
rect 33012 44038 33014 44090
rect 33194 44038 33196 44090
rect 32950 44036 32956 44038
rect 33012 44036 33036 44038
rect 33092 44036 33116 44038
rect 33172 44036 33196 44038
rect 33252 44036 33258 44038
rect 32950 44027 33258 44036
rect 32864 43852 32916 43858
rect 32864 43794 32916 43800
rect 33232 43716 33284 43722
rect 33232 43658 33284 43664
rect 33244 43382 33272 43658
rect 33324 43648 33376 43654
rect 33324 43590 33376 43596
rect 33232 43376 33284 43382
rect 33232 43318 33284 43324
rect 33244 43246 33272 43318
rect 33232 43240 33284 43246
rect 33232 43182 33284 43188
rect 32950 43004 33258 43013
rect 32950 43002 32956 43004
rect 33012 43002 33036 43004
rect 33092 43002 33116 43004
rect 33172 43002 33196 43004
rect 33252 43002 33258 43004
rect 33012 42950 33014 43002
rect 33194 42950 33196 43002
rect 32950 42948 32956 42950
rect 33012 42948 33036 42950
rect 33092 42948 33116 42950
rect 33172 42948 33196 42950
rect 33252 42948 33258 42950
rect 32950 42939 33258 42948
rect 32772 42356 32824 42362
rect 32772 42298 32824 42304
rect 32784 40594 32812 42298
rect 32950 41916 33258 41925
rect 32950 41914 32956 41916
rect 33012 41914 33036 41916
rect 33092 41914 33116 41916
rect 33172 41914 33196 41916
rect 33252 41914 33258 41916
rect 33012 41862 33014 41914
rect 33194 41862 33196 41914
rect 32950 41860 32956 41862
rect 33012 41860 33036 41862
rect 33092 41860 33116 41862
rect 33172 41860 33196 41862
rect 33252 41860 33258 41862
rect 32950 41851 33258 41860
rect 32864 41812 32916 41818
rect 32864 41754 32916 41760
rect 32876 41290 32904 41754
rect 32956 41540 33008 41546
rect 32956 41482 33008 41488
rect 32968 41414 32996 41482
rect 33336 41478 33364 43590
rect 33324 41472 33376 41478
rect 33324 41414 33376 41420
rect 32968 41386 33088 41414
rect 32876 41262 32996 41290
rect 32864 41200 32916 41206
rect 32864 41142 32916 41148
rect 32680 40588 32732 40594
rect 32680 40530 32732 40536
rect 32772 40588 32824 40594
rect 32772 40530 32824 40536
rect 32600 40446 32812 40474
rect 32588 39500 32640 39506
rect 32588 39442 32640 39448
rect 32600 38418 32628 39442
rect 32784 38418 32812 40446
rect 32588 38412 32640 38418
rect 32588 38354 32640 38360
rect 32772 38412 32824 38418
rect 32772 38354 32824 38360
rect 32496 37256 32548 37262
rect 32496 37198 32548 37204
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32404 36916 32456 36922
rect 32404 36858 32456 36864
rect 32220 36780 32272 36786
rect 32220 36722 32272 36728
rect 32312 36712 32364 36718
rect 32312 36654 32364 36660
rect 32220 35828 32272 35834
rect 32220 35770 32272 35776
rect 32232 35154 32260 35770
rect 32324 35630 32352 36654
rect 32508 36145 32536 37062
rect 32494 36136 32550 36145
rect 32494 36071 32550 36080
rect 32312 35624 32364 35630
rect 32312 35566 32364 35572
rect 32220 35148 32272 35154
rect 32220 35090 32272 35096
rect 32128 32904 32180 32910
rect 32128 32846 32180 32852
rect 32128 32360 32180 32366
rect 32128 32302 32180 32308
rect 32140 30802 32168 32302
rect 32220 32224 32272 32230
rect 32220 32166 32272 32172
rect 32232 31958 32260 32166
rect 32220 31952 32272 31958
rect 32220 31894 32272 31900
rect 32128 30796 32180 30802
rect 32128 30738 32180 30744
rect 32312 30796 32364 30802
rect 32312 30738 32364 30744
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 31944 29504 31996 29510
rect 31944 29446 31996 29452
rect 31852 27124 31904 27130
rect 31852 27066 31904 27072
rect 31852 26444 31904 26450
rect 31852 26386 31904 26392
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31668 24880 31720 24886
rect 31668 24822 31720 24828
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 31484 18828 31536 18834
rect 31484 18770 31536 18776
rect 31300 18760 31352 18766
rect 31300 18702 31352 18708
rect 30840 18352 30892 18358
rect 30840 18294 30892 18300
rect 30380 18216 30432 18222
rect 30380 18158 30432 18164
rect 30288 17604 30340 17610
rect 30288 17546 30340 17552
rect 30392 17490 30420 18158
rect 31024 17740 31076 17746
rect 31024 17682 31076 17688
rect 30932 17604 30984 17610
rect 30932 17546 30984 17552
rect 30300 17462 30420 17490
rect 30564 17536 30616 17542
rect 30564 17478 30616 17484
rect 30300 17134 30328 17462
rect 30576 17270 30604 17478
rect 30564 17264 30616 17270
rect 30484 17212 30564 17218
rect 30484 17206 30616 17212
rect 30484 17190 30604 17206
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30300 15994 30328 17070
rect 30484 16182 30512 17190
rect 30944 17134 30972 17546
rect 31036 17338 31064 17682
rect 31024 17332 31076 17338
rect 31024 17274 31076 17280
rect 31116 17332 31168 17338
rect 31116 17274 31168 17280
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 31128 16794 31156 17274
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30208 15966 30328 15994
rect 30208 15706 30236 15966
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 30484 15434 30512 16118
rect 30564 15904 30616 15910
rect 30564 15846 30616 15852
rect 30576 15570 30604 15846
rect 30564 15564 30616 15570
rect 30564 15506 30616 15512
rect 30472 15428 30524 15434
rect 30472 15370 30524 15376
rect 30104 15088 30156 15094
rect 30104 15030 30156 15036
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 30208 14414 30236 14758
rect 30300 14550 30328 14826
rect 30564 14612 30616 14618
rect 30564 14554 30616 14560
rect 30288 14544 30340 14550
rect 30288 14486 30340 14492
rect 30196 14408 30248 14414
rect 30196 14350 30248 14356
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29368 7404 29420 7410
rect 29368 7346 29420 7352
rect 29460 3596 29512 3602
rect 29460 3538 29512 3544
rect 29276 1828 29328 1834
rect 29276 1770 29328 1776
rect 29472 800 29500 3538
rect 29748 3534 29776 13806
rect 30300 12986 30328 14350
rect 30576 13938 30604 14554
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 30104 9988 30156 9994
rect 30104 9930 30156 9936
rect 29920 9920 29972 9926
rect 29920 9862 29972 9868
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29932 2446 29960 9862
rect 30116 3534 30144 9930
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30484 2922 30512 12922
rect 30576 12782 30604 13330
rect 30668 12986 30696 16526
rect 31588 15094 31616 23666
rect 31680 23050 31708 24822
rect 31864 23508 31892 26386
rect 31956 25294 31984 29446
rect 32140 29034 32168 30194
rect 32220 29844 32272 29850
rect 32220 29786 32272 29792
rect 32128 29028 32180 29034
rect 32128 28970 32180 28976
rect 32036 28960 32088 28966
rect 32036 28902 32088 28908
rect 32048 28150 32076 28902
rect 32128 28212 32180 28218
rect 32128 28154 32180 28160
rect 32036 28144 32088 28150
rect 32036 28086 32088 28092
rect 32036 27532 32088 27538
rect 32036 27474 32088 27480
rect 32048 26450 32076 27474
rect 32036 26444 32088 26450
rect 32036 26386 32088 26392
rect 32140 26330 32168 28154
rect 32232 27538 32260 29786
rect 32324 28014 32352 30738
rect 32402 30696 32458 30705
rect 32402 30631 32458 30640
rect 32416 30598 32444 30631
rect 32404 30592 32456 30598
rect 32404 30534 32456 30540
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 32416 29170 32444 29446
rect 32404 29164 32456 29170
rect 32404 29106 32456 29112
rect 32312 28008 32364 28014
rect 32508 27962 32536 36071
rect 32600 35834 32628 38354
rect 32680 37868 32732 37874
rect 32680 37810 32732 37816
rect 32692 36174 32720 37810
rect 32784 36242 32812 38354
rect 32772 36236 32824 36242
rect 32772 36178 32824 36184
rect 32680 36168 32732 36174
rect 32680 36110 32732 36116
rect 32784 35986 32812 36178
rect 32692 35958 32812 35986
rect 32588 35828 32640 35834
rect 32588 35770 32640 35776
rect 32692 34610 32720 35958
rect 32772 35760 32824 35766
rect 32770 35728 32772 35737
rect 32824 35728 32826 35737
rect 32770 35663 32826 35672
rect 32876 35630 32904 41142
rect 32968 40934 32996 41262
rect 33060 41002 33088 41386
rect 33048 40996 33100 41002
rect 33048 40938 33100 40944
rect 32956 40928 33008 40934
rect 32956 40870 33008 40876
rect 32950 40828 33258 40837
rect 32950 40826 32956 40828
rect 33012 40826 33036 40828
rect 33092 40826 33116 40828
rect 33172 40826 33196 40828
rect 33252 40826 33258 40828
rect 33012 40774 33014 40826
rect 33194 40774 33196 40826
rect 32950 40772 32956 40774
rect 33012 40772 33036 40774
rect 33092 40772 33116 40774
rect 33172 40772 33196 40774
rect 33252 40772 33258 40774
rect 32950 40763 33258 40772
rect 32950 39740 33258 39749
rect 32950 39738 32956 39740
rect 33012 39738 33036 39740
rect 33092 39738 33116 39740
rect 33172 39738 33196 39740
rect 33252 39738 33258 39740
rect 33012 39686 33014 39738
rect 33194 39686 33196 39738
rect 32950 39684 32956 39686
rect 33012 39684 33036 39686
rect 33092 39684 33116 39686
rect 33172 39684 33196 39686
rect 33252 39684 33258 39686
rect 32950 39675 33258 39684
rect 33324 38956 33376 38962
rect 33324 38898 33376 38904
rect 32950 38652 33258 38661
rect 32950 38650 32956 38652
rect 33012 38650 33036 38652
rect 33092 38650 33116 38652
rect 33172 38650 33196 38652
rect 33252 38650 33258 38652
rect 33012 38598 33014 38650
rect 33194 38598 33196 38650
rect 32950 38596 32956 38598
rect 33012 38596 33036 38598
rect 33092 38596 33116 38598
rect 33172 38596 33196 38598
rect 33252 38596 33258 38598
rect 32950 38587 33258 38596
rect 32950 37564 33258 37573
rect 32950 37562 32956 37564
rect 33012 37562 33036 37564
rect 33092 37562 33116 37564
rect 33172 37562 33196 37564
rect 33252 37562 33258 37564
rect 33012 37510 33014 37562
rect 33194 37510 33196 37562
rect 32950 37508 32956 37510
rect 33012 37508 33036 37510
rect 33092 37508 33116 37510
rect 33172 37508 33196 37510
rect 33252 37508 33258 37510
rect 32950 37499 33258 37508
rect 33336 37194 33364 38898
rect 33428 37806 33456 45426
rect 33980 45422 34008 53994
rect 34992 53582 35020 56200
rect 35728 54194 35756 56200
rect 36464 54194 36492 56200
rect 37200 54262 37228 56200
rect 37936 55214 37964 56200
rect 37844 55186 37964 55214
rect 37740 54324 37792 54330
rect 37740 54266 37792 54272
rect 37188 54256 37240 54262
rect 37188 54198 37240 54204
rect 35716 54188 35768 54194
rect 35716 54130 35768 54136
rect 36452 54188 36504 54194
rect 36452 54130 36504 54136
rect 35256 53984 35308 53990
rect 35256 53926 35308 53932
rect 36544 53984 36596 53990
rect 36544 53926 36596 53932
rect 37188 53984 37240 53990
rect 37188 53926 37240 53932
rect 37648 53984 37700 53990
rect 37648 53926 37700 53932
rect 34980 53576 35032 53582
rect 34980 53518 35032 53524
rect 33968 45416 34020 45422
rect 33968 45358 34020 45364
rect 34152 45416 34204 45422
rect 34152 45358 34204 45364
rect 33508 45280 33560 45286
rect 33508 45222 33560 45228
rect 33520 40594 33548 45222
rect 33876 41064 33928 41070
rect 33876 41006 33928 41012
rect 33508 40588 33560 40594
rect 33508 40530 33560 40536
rect 33600 40384 33652 40390
rect 33600 40326 33652 40332
rect 33692 40384 33744 40390
rect 33692 40326 33744 40332
rect 33508 39500 33560 39506
rect 33508 39442 33560 39448
rect 33520 39098 33548 39442
rect 33612 39098 33640 40326
rect 33508 39092 33560 39098
rect 33508 39034 33560 39040
rect 33600 39092 33652 39098
rect 33600 39034 33652 39040
rect 33508 38004 33560 38010
rect 33508 37946 33560 37952
rect 33520 37913 33548 37946
rect 33506 37904 33562 37913
rect 33506 37839 33562 37848
rect 33416 37800 33468 37806
rect 33416 37742 33468 37748
rect 33324 37188 33376 37194
rect 33324 37130 33376 37136
rect 33428 36938 33456 37742
rect 33704 37233 33732 40326
rect 33888 40118 33916 41006
rect 33876 40112 33928 40118
rect 33876 40054 33928 40060
rect 33784 39976 33836 39982
rect 33784 39918 33836 39924
rect 33796 38826 33824 39918
rect 33784 38820 33836 38826
rect 33784 38762 33836 38768
rect 33690 37224 33746 37233
rect 33690 37159 33746 37168
rect 33336 36910 33456 36938
rect 32950 36476 33258 36485
rect 32950 36474 32956 36476
rect 33012 36474 33036 36476
rect 33092 36474 33116 36476
rect 33172 36474 33196 36476
rect 33252 36474 33258 36476
rect 33012 36422 33014 36474
rect 33194 36422 33196 36474
rect 32950 36420 32956 36422
rect 33012 36420 33036 36422
rect 33092 36420 33116 36422
rect 33172 36420 33196 36422
rect 33252 36420 33258 36422
rect 32950 36411 33258 36420
rect 33048 36100 33100 36106
rect 33048 36042 33100 36048
rect 33140 36100 33192 36106
rect 33140 36042 33192 36048
rect 33060 35834 33088 36042
rect 33048 35828 33100 35834
rect 33048 35770 33100 35776
rect 32864 35624 32916 35630
rect 32864 35566 32916 35572
rect 33152 35494 33180 36042
rect 33140 35488 33192 35494
rect 33140 35430 33192 35436
rect 32950 35388 33258 35397
rect 32950 35386 32956 35388
rect 33012 35386 33036 35388
rect 33092 35386 33116 35388
rect 33172 35386 33196 35388
rect 33252 35386 33258 35388
rect 33012 35334 33014 35386
rect 33194 35334 33196 35386
rect 32950 35332 32956 35334
rect 33012 35332 33036 35334
rect 33092 35332 33116 35334
rect 33172 35332 33196 35334
rect 33252 35332 33258 35334
rect 32950 35323 33258 35332
rect 32772 34944 32824 34950
rect 32772 34886 32824 34892
rect 32784 34746 32812 34886
rect 32772 34740 32824 34746
rect 32772 34682 32824 34688
rect 32588 34604 32640 34610
rect 32588 34546 32640 34552
rect 32680 34604 32732 34610
rect 32680 34546 32732 34552
rect 32600 33930 32628 34546
rect 32950 34300 33258 34309
rect 32950 34298 32956 34300
rect 33012 34298 33036 34300
rect 33092 34298 33116 34300
rect 33172 34298 33196 34300
rect 33252 34298 33258 34300
rect 33012 34246 33014 34298
rect 33194 34246 33196 34298
rect 32950 34244 32956 34246
rect 33012 34244 33036 34246
rect 33092 34244 33116 34246
rect 33172 34244 33196 34246
rect 33252 34244 33258 34246
rect 32950 34235 33258 34244
rect 32588 33924 32640 33930
rect 32588 33866 32640 33872
rect 32950 33212 33258 33221
rect 32950 33210 32956 33212
rect 33012 33210 33036 33212
rect 33092 33210 33116 33212
rect 33172 33210 33196 33212
rect 33252 33210 33258 33212
rect 33012 33158 33014 33210
rect 33194 33158 33196 33210
rect 32950 33156 32956 33158
rect 33012 33156 33036 33158
rect 33092 33156 33116 33158
rect 33172 33156 33196 33158
rect 33252 33156 33258 33158
rect 32950 33147 33258 33156
rect 32588 33108 32640 33114
rect 32588 33050 32640 33056
rect 32600 30598 32628 33050
rect 32770 33008 32826 33017
rect 32770 32943 32826 32952
rect 32784 31890 32812 32943
rect 32950 32124 33258 32133
rect 32950 32122 32956 32124
rect 33012 32122 33036 32124
rect 33092 32122 33116 32124
rect 33172 32122 33196 32124
rect 33252 32122 33258 32124
rect 33012 32070 33014 32122
rect 33194 32070 33196 32122
rect 32950 32068 32956 32070
rect 33012 32068 33036 32070
rect 33092 32068 33116 32070
rect 33172 32068 33196 32070
rect 33252 32068 33258 32070
rect 32950 32059 33258 32068
rect 32772 31884 32824 31890
rect 32772 31826 32824 31832
rect 32784 31754 32812 31826
rect 32692 31726 32812 31754
rect 32588 30592 32640 30598
rect 32588 30534 32640 30540
rect 32600 28966 32628 30534
rect 32588 28960 32640 28966
rect 32588 28902 32640 28908
rect 32312 27950 32364 27956
rect 32220 27532 32272 27538
rect 32220 27474 32272 27480
rect 32324 27402 32352 27950
rect 32416 27934 32536 27962
rect 32312 27396 32364 27402
rect 32232 27356 32312 27384
rect 32232 26450 32260 27356
rect 32312 27338 32364 27344
rect 32220 26444 32272 26450
rect 32220 26386 32272 26392
rect 32036 26308 32088 26314
rect 32140 26302 32260 26330
rect 32416 26314 32444 27934
rect 32588 27872 32640 27878
rect 32508 27820 32588 27826
rect 32508 27814 32640 27820
rect 32508 27798 32628 27814
rect 32508 26314 32536 27798
rect 32586 27432 32642 27441
rect 32586 27367 32642 27376
rect 32600 27334 32628 27367
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32600 26314 32628 27270
rect 32036 26250 32088 26256
rect 31944 25288 31996 25294
rect 31944 25230 31996 25236
rect 31772 23480 31892 23508
rect 31668 23044 31720 23050
rect 31668 22986 31720 22992
rect 31680 22166 31708 22986
rect 31772 22982 31800 23480
rect 31852 23316 31904 23322
rect 31852 23258 31904 23264
rect 31760 22976 31812 22982
rect 31760 22918 31812 22924
rect 31772 22234 31800 22918
rect 31760 22228 31812 22234
rect 31760 22170 31812 22176
rect 31668 22160 31720 22166
rect 31668 22102 31720 22108
rect 31680 21554 31708 22102
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31668 21548 31720 21554
rect 31668 21490 31720 21496
rect 31772 21010 31800 21626
rect 31864 21486 31892 23258
rect 31942 21992 31998 22001
rect 31942 21927 31998 21936
rect 31852 21480 31904 21486
rect 31852 21422 31904 21428
rect 31760 21004 31812 21010
rect 31760 20946 31812 20952
rect 31760 20052 31812 20058
rect 31760 19994 31812 20000
rect 31772 16130 31800 19994
rect 31956 19854 31984 21927
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31944 19712 31996 19718
rect 31944 19654 31996 19660
rect 31956 18290 31984 19654
rect 31944 18284 31996 18290
rect 31944 18226 31996 18232
rect 31772 16102 31892 16130
rect 31576 15088 31628 15094
rect 31576 15030 31628 15036
rect 31024 14952 31076 14958
rect 31024 14894 31076 14900
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30564 12776 30616 12782
rect 30564 12718 30616 12724
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30472 2916 30524 2922
rect 30472 2858 30524 2864
rect 30288 2508 30340 2514
rect 30208 2468 30288 2496
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 30208 800 30236 2468
rect 30288 2450 30340 2456
rect 30944 800 30972 3538
rect 31036 2446 31064 14894
rect 31760 13184 31812 13190
rect 31760 13126 31812 13132
rect 31772 7478 31800 13126
rect 31864 10062 31892 16102
rect 31956 12986 31984 18226
rect 32048 16658 32076 26250
rect 32128 26240 32180 26246
rect 32128 26182 32180 26188
rect 32140 22001 32168 26182
rect 32232 25770 32260 26302
rect 32404 26308 32456 26314
rect 32404 26250 32456 26256
rect 32496 26308 32548 26314
rect 32496 26250 32548 26256
rect 32588 26308 32640 26314
rect 32588 26250 32640 26256
rect 32508 25838 32536 26250
rect 32692 26194 32720 31726
rect 32864 31136 32916 31142
rect 32864 31078 32916 31084
rect 32772 30048 32824 30054
rect 32772 29990 32824 29996
rect 32784 27606 32812 29990
rect 32876 28626 32904 31078
rect 32950 31036 33258 31045
rect 32950 31034 32956 31036
rect 33012 31034 33036 31036
rect 33092 31034 33116 31036
rect 33172 31034 33196 31036
rect 33252 31034 33258 31036
rect 33012 30982 33014 31034
rect 33194 30982 33196 31034
rect 32950 30980 32956 30982
rect 33012 30980 33036 30982
rect 33092 30980 33116 30982
rect 33172 30980 33196 30982
rect 33252 30980 33258 30982
rect 32950 30971 33258 30980
rect 32950 29948 33258 29957
rect 32950 29946 32956 29948
rect 33012 29946 33036 29948
rect 33092 29946 33116 29948
rect 33172 29946 33196 29948
rect 33252 29946 33258 29948
rect 33012 29894 33014 29946
rect 33194 29894 33196 29946
rect 32950 29892 32956 29894
rect 33012 29892 33036 29894
rect 33092 29892 33116 29894
rect 33172 29892 33196 29894
rect 33252 29892 33258 29894
rect 32950 29883 33258 29892
rect 32950 28860 33258 28869
rect 32950 28858 32956 28860
rect 33012 28858 33036 28860
rect 33092 28858 33116 28860
rect 33172 28858 33196 28860
rect 33252 28858 33258 28860
rect 33012 28806 33014 28858
rect 33194 28806 33196 28858
rect 32950 28804 32956 28806
rect 33012 28804 33036 28806
rect 33092 28804 33116 28806
rect 33172 28804 33196 28806
rect 33252 28804 33258 28806
rect 32950 28795 33258 28804
rect 33336 28642 33364 36910
rect 33508 36372 33560 36378
rect 33508 36314 33560 36320
rect 33416 34944 33468 34950
rect 33414 34912 33416 34921
rect 33468 34912 33470 34921
rect 33414 34847 33470 34856
rect 33520 33402 33548 36314
rect 33704 34218 33732 37159
rect 33796 34474 33824 38762
rect 33980 38298 34008 45358
rect 34164 43178 34192 45358
rect 35268 44742 35296 53926
rect 35348 53440 35400 53446
rect 35348 53382 35400 53388
rect 35360 44946 35388 53382
rect 35992 45008 36044 45014
rect 35992 44950 36044 44956
rect 35348 44940 35400 44946
rect 35348 44882 35400 44888
rect 35532 44940 35584 44946
rect 35532 44882 35584 44888
rect 35256 44736 35308 44742
rect 35254 44704 35256 44713
rect 35308 44704 35310 44713
rect 35254 44639 35310 44648
rect 34796 43376 34848 43382
rect 34796 43318 34848 43324
rect 34520 43308 34572 43314
rect 34520 43250 34572 43256
rect 34152 43172 34204 43178
rect 34152 43114 34204 43120
rect 34060 43104 34112 43110
rect 34060 43046 34112 43052
rect 34072 42344 34100 43046
rect 34532 42702 34560 43250
rect 34520 42696 34572 42702
rect 34520 42638 34572 42644
rect 34532 42362 34560 42638
rect 34520 42356 34572 42362
rect 34072 42316 34192 42344
rect 34164 41682 34192 42316
rect 34520 42298 34572 42304
rect 34532 41682 34560 42298
rect 34152 41676 34204 41682
rect 34152 41618 34204 41624
rect 34520 41676 34572 41682
rect 34520 41618 34572 41624
rect 34704 41676 34756 41682
rect 34704 41618 34756 41624
rect 34164 40594 34192 41618
rect 34428 41540 34480 41546
rect 34428 41482 34480 41488
rect 34244 41472 34296 41478
rect 34244 41414 34296 41420
rect 34152 40588 34204 40594
rect 34152 40530 34204 40536
rect 34152 40452 34204 40458
rect 34152 40394 34204 40400
rect 34060 39840 34112 39846
rect 34060 39782 34112 39788
rect 34072 39574 34100 39782
rect 34060 39568 34112 39574
rect 34060 39510 34112 39516
rect 34164 38418 34192 40394
rect 34256 38894 34284 41414
rect 34440 40662 34468 41482
rect 34428 40656 34480 40662
rect 34428 40598 34480 40604
rect 34716 40050 34744 41618
rect 34808 40934 34836 43318
rect 35544 42158 35572 44882
rect 35900 43172 35952 43178
rect 35900 43114 35952 43120
rect 35912 42294 35940 43114
rect 35900 42288 35952 42294
rect 35900 42230 35952 42236
rect 35532 42152 35584 42158
rect 35532 42094 35584 42100
rect 34888 42016 34940 42022
rect 34888 41958 34940 41964
rect 34900 41274 34928 41958
rect 35544 41818 35572 42094
rect 35532 41812 35584 41818
rect 35532 41754 35584 41760
rect 35808 41472 35860 41478
rect 35808 41414 35860 41420
rect 35820 41386 35940 41414
rect 34888 41268 34940 41274
rect 34888 41210 34940 41216
rect 34796 40928 34848 40934
rect 34796 40870 34848 40876
rect 34704 40044 34756 40050
rect 34704 39986 34756 39992
rect 34336 39840 34388 39846
rect 34336 39782 34388 39788
rect 34348 39030 34376 39782
rect 34716 39438 34744 39986
rect 34520 39432 34572 39438
rect 34520 39374 34572 39380
rect 34704 39432 34756 39438
rect 34704 39374 34756 39380
rect 34428 39092 34480 39098
rect 34428 39034 34480 39040
rect 34336 39024 34388 39030
rect 34336 38966 34388 38972
rect 34244 38888 34296 38894
rect 34440 38842 34468 39034
rect 34244 38830 34296 38836
rect 34348 38814 34468 38842
rect 34152 38412 34204 38418
rect 34152 38354 34204 38360
rect 33980 38270 34192 38298
rect 33968 38208 34020 38214
rect 33968 38150 34020 38156
rect 34060 38208 34112 38214
rect 34060 38150 34112 38156
rect 33980 38010 34008 38150
rect 33968 38004 34020 38010
rect 33968 37946 34020 37952
rect 33876 37868 33928 37874
rect 33876 37810 33928 37816
rect 33888 37466 33916 37810
rect 33876 37460 33928 37466
rect 33876 37402 33928 37408
rect 33968 36712 34020 36718
rect 33968 36654 34020 36660
rect 33876 36644 33928 36650
rect 33876 36586 33928 36592
rect 33888 35290 33916 36586
rect 33876 35284 33928 35290
rect 33876 35226 33928 35232
rect 33784 34468 33836 34474
rect 33784 34410 33836 34416
rect 33704 34190 33824 34218
rect 33692 33856 33744 33862
rect 33692 33798 33744 33804
rect 33520 33374 33640 33402
rect 33416 31204 33468 31210
rect 33416 31146 33468 31152
rect 32864 28620 32916 28626
rect 32864 28562 32916 28568
rect 33244 28614 33364 28642
rect 32864 28416 32916 28422
rect 32864 28358 32916 28364
rect 32772 27600 32824 27606
rect 32772 27542 32824 27548
rect 32600 26166 32720 26194
rect 32496 25832 32548 25838
rect 32496 25774 32548 25780
rect 32220 25764 32272 25770
rect 32220 25706 32272 25712
rect 32232 24614 32260 25706
rect 32600 25514 32628 26166
rect 32680 26036 32732 26042
rect 32680 25978 32732 25984
rect 32508 25486 32628 25514
rect 32312 24676 32364 24682
rect 32312 24618 32364 24624
rect 32220 24608 32272 24614
rect 32220 24550 32272 24556
rect 32324 23730 32352 24618
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32312 22432 32364 22438
rect 32312 22374 32364 22380
rect 32126 21992 32182 22001
rect 32126 21927 32182 21936
rect 32128 21888 32180 21894
rect 32128 21830 32180 21836
rect 32140 21350 32168 21830
rect 32220 21480 32272 21486
rect 32220 21422 32272 21428
rect 32128 21344 32180 21350
rect 32128 21286 32180 21292
rect 32128 20800 32180 20806
rect 32128 20742 32180 20748
rect 32140 16998 32168 20742
rect 32232 20398 32260 21422
rect 32220 20392 32272 20398
rect 32220 20334 32272 20340
rect 32324 19854 32352 22374
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32232 17746 32260 19790
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 32416 17202 32444 24550
rect 32508 23798 32536 25486
rect 32588 25356 32640 25362
rect 32588 25298 32640 25304
rect 32496 23792 32548 23798
rect 32496 23734 32548 23740
rect 32600 23322 32628 25298
rect 32692 25265 32720 25978
rect 32784 25974 32812 27542
rect 32772 25968 32824 25974
rect 32772 25910 32824 25916
rect 32678 25256 32734 25265
rect 32678 25191 32734 25200
rect 32772 25152 32824 25158
rect 32772 25094 32824 25100
rect 32680 24744 32732 24750
rect 32680 24686 32732 24692
rect 32692 24206 32720 24686
rect 32680 24200 32732 24206
rect 32680 24142 32732 24148
rect 32680 23656 32732 23662
rect 32680 23598 32732 23604
rect 32588 23316 32640 23322
rect 32588 23258 32640 23264
rect 32496 23044 32548 23050
rect 32496 22986 32548 22992
rect 32588 23044 32640 23050
rect 32588 22986 32640 22992
rect 32508 21554 32536 22986
rect 32600 21690 32628 22986
rect 32692 22778 32720 23598
rect 32680 22772 32732 22778
rect 32680 22714 32732 22720
rect 32680 22228 32732 22234
rect 32680 22170 32732 22176
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32496 21548 32548 21554
rect 32496 21490 32548 21496
rect 32508 21146 32536 21490
rect 32496 21140 32548 21146
rect 32496 21082 32548 21088
rect 32588 20256 32640 20262
rect 32588 20198 32640 20204
rect 32496 18828 32548 18834
rect 32496 18770 32548 18776
rect 32508 18358 32536 18770
rect 32496 18352 32548 18358
rect 32496 18294 32548 18300
rect 32508 17882 32536 18294
rect 32496 17876 32548 17882
rect 32496 17818 32548 17824
rect 32404 17196 32456 17202
rect 32404 17138 32456 17144
rect 32128 16992 32180 16998
rect 32128 16934 32180 16940
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 32036 16652 32088 16658
rect 32036 16594 32088 16600
rect 31944 12980 31996 12986
rect 31944 12922 31996 12928
rect 32140 12434 32168 16934
rect 32220 15020 32272 15026
rect 32220 14962 32272 14968
rect 32232 14618 32260 14962
rect 32220 14612 32272 14618
rect 32220 14554 32272 14560
rect 32324 13190 32352 16934
rect 32496 16040 32548 16046
rect 32496 15982 32548 15988
rect 32404 15360 32456 15366
rect 32404 15302 32456 15308
rect 32312 13184 32364 13190
rect 32312 13126 32364 13132
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32048 12406 32168 12434
rect 31852 10056 31904 10062
rect 31852 9998 31904 10004
rect 32048 9654 32076 12406
rect 32036 9648 32088 9654
rect 32036 9590 32088 9596
rect 32324 8566 32352 12922
rect 32416 12918 32444 15302
rect 32508 14482 32536 15982
rect 32600 15502 32628 20198
rect 32692 19922 32720 22170
rect 32784 20584 32812 25094
rect 32876 24818 32904 28358
rect 33244 27928 33272 28614
rect 33324 28552 33376 28558
rect 33324 28494 33376 28500
rect 33336 28098 33364 28494
rect 33428 28218 33456 31146
rect 33508 29232 33560 29238
rect 33508 29174 33560 29180
rect 33416 28212 33468 28218
rect 33416 28154 33468 28160
rect 33336 28070 33456 28098
rect 33244 27900 33364 27928
rect 32950 27772 33258 27781
rect 32950 27770 32956 27772
rect 33012 27770 33036 27772
rect 33092 27770 33116 27772
rect 33172 27770 33196 27772
rect 33252 27770 33258 27772
rect 33012 27718 33014 27770
rect 33194 27718 33196 27770
rect 32950 27716 32956 27718
rect 33012 27716 33036 27718
rect 33092 27716 33116 27718
rect 33172 27716 33196 27718
rect 33252 27716 33258 27718
rect 32950 27707 33258 27716
rect 33230 27024 33286 27033
rect 33230 26959 33286 26968
rect 33244 26926 33272 26959
rect 33232 26920 33284 26926
rect 33232 26862 33284 26868
rect 32950 26684 33258 26693
rect 32950 26682 32956 26684
rect 33012 26682 33036 26684
rect 33092 26682 33116 26684
rect 33172 26682 33196 26684
rect 33252 26682 33258 26684
rect 33012 26630 33014 26682
rect 33194 26630 33196 26682
rect 32950 26628 32956 26630
rect 33012 26628 33036 26630
rect 33092 26628 33116 26630
rect 33172 26628 33196 26630
rect 33252 26628 33258 26630
rect 32950 26619 33258 26628
rect 32950 25596 33258 25605
rect 32950 25594 32956 25596
rect 33012 25594 33036 25596
rect 33092 25594 33116 25596
rect 33172 25594 33196 25596
rect 33252 25594 33258 25596
rect 33012 25542 33014 25594
rect 33194 25542 33196 25594
rect 32950 25540 32956 25542
rect 33012 25540 33036 25542
rect 33092 25540 33116 25542
rect 33172 25540 33196 25542
rect 33252 25540 33258 25542
rect 32950 25531 33258 25540
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32864 24268 32916 24274
rect 32864 24210 32916 24216
rect 32876 22574 32904 24210
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32864 22568 32916 22574
rect 32864 22510 32916 22516
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 32876 21146 32904 21966
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32864 21140 32916 21146
rect 32864 21082 32916 21088
rect 32864 20596 32916 20602
rect 32784 20556 32864 20584
rect 32864 20538 32916 20544
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32680 19916 32732 19922
rect 32680 19858 32732 19864
rect 33336 19854 33364 27900
rect 33428 24290 33456 28070
rect 33520 24426 33548 29174
rect 33612 24562 33640 33374
rect 33704 30326 33732 33798
rect 33692 30320 33744 30326
rect 33692 30262 33744 30268
rect 33796 29238 33824 34190
rect 33888 33590 33916 35226
rect 33980 34542 34008 36654
rect 34072 36310 34100 38150
rect 34164 36378 34192 38270
rect 34244 37120 34296 37126
rect 34244 37062 34296 37068
rect 34152 36372 34204 36378
rect 34152 36314 34204 36320
rect 34060 36304 34112 36310
rect 34060 36246 34112 36252
rect 34060 36032 34112 36038
rect 34060 35974 34112 35980
rect 33968 34536 34020 34542
rect 33968 34478 34020 34484
rect 33876 33584 33928 33590
rect 33876 33526 33928 33532
rect 33980 33522 34008 34478
rect 34072 33658 34100 35974
rect 34256 35442 34284 37062
rect 34164 35414 34284 35442
rect 34060 33652 34112 33658
rect 34060 33594 34112 33600
rect 33968 33516 34020 33522
rect 33968 33458 34020 33464
rect 34060 32768 34112 32774
rect 34060 32710 34112 32716
rect 34072 32502 34100 32710
rect 34060 32496 34112 32502
rect 34060 32438 34112 32444
rect 34164 31754 34192 35414
rect 34244 33448 34296 33454
rect 34244 33390 34296 33396
rect 33980 31726 34192 31754
rect 33876 31340 33928 31346
rect 33876 31282 33928 31288
rect 33888 30433 33916 31282
rect 33874 30424 33930 30433
rect 33874 30359 33930 30368
rect 33980 30190 34008 31726
rect 34058 31376 34114 31385
rect 34058 31311 34114 31320
rect 34072 31278 34100 31311
rect 34060 31272 34112 31278
rect 34060 31214 34112 31220
rect 34150 30288 34206 30297
rect 34150 30223 34152 30232
rect 34204 30223 34206 30232
rect 34152 30194 34204 30200
rect 33968 30184 34020 30190
rect 33968 30126 34020 30132
rect 33876 30116 33928 30122
rect 33876 30058 33928 30064
rect 34060 30116 34112 30122
rect 34060 30058 34112 30064
rect 33888 29714 33916 30058
rect 33876 29708 33928 29714
rect 33876 29650 33928 29656
rect 33784 29232 33836 29238
rect 33784 29174 33836 29180
rect 33968 29096 34020 29102
rect 33968 29038 34020 29044
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33796 27946 33824 28494
rect 33876 28144 33928 28150
rect 33876 28086 33928 28092
rect 33784 27940 33836 27946
rect 33784 27882 33836 27888
rect 33888 27146 33916 28086
rect 33980 27402 34008 29038
rect 33968 27396 34020 27402
rect 33968 27338 34020 27344
rect 33796 27118 33916 27146
rect 33690 27024 33746 27033
rect 33690 26959 33746 26968
rect 33704 24818 33732 26959
rect 33796 26314 33824 27118
rect 33876 27056 33928 27062
rect 33876 26998 33928 27004
rect 33888 26450 33916 26998
rect 34072 26926 34100 30058
rect 34164 29306 34192 30194
rect 34256 29646 34284 33390
rect 34244 29640 34296 29646
rect 34244 29582 34296 29588
rect 34152 29300 34204 29306
rect 34152 29242 34204 29248
rect 34152 28620 34204 28626
rect 34152 28562 34204 28568
rect 34164 27878 34192 28562
rect 34152 27872 34204 27878
rect 34152 27814 34204 27820
rect 34060 26920 34112 26926
rect 34060 26862 34112 26868
rect 33968 26784 34020 26790
rect 33968 26726 34020 26732
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 33784 26308 33836 26314
rect 33784 26250 33836 26256
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33888 24750 33916 26386
rect 33980 25362 34008 26726
rect 34072 25514 34100 26862
rect 34152 26852 34204 26858
rect 34348 26840 34376 38814
rect 34428 38548 34480 38554
rect 34428 38490 34480 38496
rect 34440 37126 34468 38490
rect 34428 37120 34480 37126
rect 34428 37062 34480 37068
rect 34532 35018 34560 39374
rect 34716 38418 34744 39374
rect 34900 38894 34928 41210
rect 35716 40928 35768 40934
rect 35716 40870 35768 40876
rect 35072 40180 35124 40186
rect 35072 40122 35124 40128
rect 34980 39296 35032 39302
rect 34980 39238 35032 39244
rect 34888 38888 34940 38894
rect 34888 38830 34940 38836
rect 34992 38758 35020 39238
rect 34980 38752 35032 38758
rect 34980 38694 35032 38700
rect 34796 38480 34848 38486
rect 34796 38422 34848 38428
rect 34704 38412 34756 38418
rect 34704 38354 34756 38360
rect 34716 37874 34744 38354
rect 34704 37868 34756 37874
rect 34704 37810 34756 37816
rect 34612 36168 34664 36174
rect 34612 36110 34664 36116
rect 34520 35012 34572 35018
rect 34520 34954 34572 34960
rect 34624 34678 34652 36110
rect 34704 35624 34756 35630
rect 34704 35566 34756 35572
rect 34612 34672 34664 34678
rect 34612 34614 34664 34620
rect 34716 33454 34744 35566
rect 34704 33448 34756 33454
rect 34704 33390 34756 33396
rect 34612 32836 34664 32842
rect 34612 32778 34664 32784
rect 34520 32224 34572 32230
rect 34520 32166 34572 32172
rect 34428 30252 34480 30258
rect 34428 30194 34480 30200
rect 34440 29850 34468 30194
rect 34428 29844 34480 29850
rect 34428 29786 34480 29792
rect 34428 29300 34480 29306
rect 34428 29242 34480 29248
rect 34204 26812 34376 26840
rect 34152 26794 34204 26800
rect 34072 25486 34376 25514
rect 33968 25356 34020 25362
rect 33968 25298 34020 25304
rect 34060 25356 34112 25362
rect 34060 25298 34112 25304
rect 33876 24744 33928 24750
rect 33876 24686 33928 24692
rect 33612 24534 34008 24562
rect 33520 24398 33824 24426
rect 33428 24262 33548 24290
rect 33416 24200 33468 24206
rect 33416 24142 33468 24148
rect 33428 24070 33456 24142
rect 33416 24064 33468 24070
rect 33416 24006 33468 24012
rect 33520 22166 33548 24262
rect 33692 23724 33744 23730
rect 33692 23666 33744 23672
rect 33704 23118 33732 23666
rect 33692 23112 33744 23118
rect 33692 23054 33744 23060
rect 33600 22976 33652 22982
rect 33600 22918 33652 22924
rect 33508 22160 33560 22166
rect 33508 22102 33560 22108
rect 33612 21842 33640 22918
rect 33520 21814 33640 21842
rect 33520 21622 33548 21814
rect 33508 21616 33560 21622
rect 33508 21558 33560 21564
rect 33324 19848 33376 19854
rect 33324 19790 33376 19796
rect 33324 19712 33376 19718
rect 33324 19654 33376 19660
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32864 18896 32916 18902
rect 32864 18838 32916 18844
rect 32876 16998 32904 18838
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32864 16992 32916 16998
rect 32864 16934 32916 16940
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32864 15904 32916 15910
rect 32864 15846 32916 15852
rect 32588 15496 32640 15502
rect 32588 15438 32640 15444
rect 32876 14958 32904 15846
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32864 14952 32916 14958
rect 32864 14894 32916 14900
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32496 14476 32548 14482
rect 32496 14418 32548 14424
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32404 12912 32456 12918
rect 32404 12854 32456 12860
rect 32312 8560 32364 8566
rect 32312 8502 32364 8508
rect 31760 7472 31812 7478
rect 31760 7414 31812 7420
rect 32416 6730 32444 12854
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32404 6724 32456 6730
rect 32404 6666 32456 6672
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 33336 3058 33364 19654
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 33508 17128 33560 17134
rect 33508 17070 33560 17076
rect 33416 15904 33468 15910
rect 33416 15846 33468 15852
rect 33428 15502 33456 15846
rect 33520 15570 33548 17070
rect 33508 15564 33560 15570
rect 33508 15506 33560 15512
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 33612 15434 33640 18362
rect 33796 17746 33824 24398
rect 33876 24064 33928 24070
rect 33876 24006 33928 24012
rect 33888 23798 33916 24006
rect 33876 23792 33928 23798
rect 33876 23734 33928 23740
rect 33980 19854 34008 24534
rect 34072 23866 34100 25298
rect 34152 25152 34204 25158
rect 34152 25094 34204 25100
rect 34060 23860 34112 23866
rect 34060 23802 34112 23808
rect 34072 21486 34100 23802
rect 34164 22710 34192 25094
rect 34244 24744 34296 24750
rect 34244 24686 34296 24692
rect 34256 23322 34284 24686
rect 34348 23526 34376 25486
rect 34440 24410 34468 29242
rect 34532 28014 34560 32166
rect 34624 30666 34652 32778
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34612 30660 34664 30666
rect 34612 30602 34664 30608
rect 34612 30116 34664 30122
rect 34612 30058 34664 30064
rect 34520 28008 34572 28014
rect 34520 27950 34572 27956
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 34428 24404 34480 24410
rect 34428 24346 34480 24352
rect 34532 24290 34560 25842
rect 34624 25294 34652 30058
rect 34716 29850 34744 31758
rect 34808 31521 34836 38422
rect 35084 38214 35112 40122
rect 35624 39976 35676 39982
rect 35624 39918 35676 39924
rect 35256 39296 35308 39302
rect 35256 39238 35308 39244
rect 35268 38282 35296 39238
rect 35636 39114 35664 39918
rect 35360 39098 35664 39114
rect 35348 39092 35676 39098
rect 35400 39086 35624 39092
rect 35348 39034 35400 39040
rect 35624 39034 35676 39040
rect 35440 39024 35492 39030
rect 35440 38966 35492 38972
rect 35256 38276 35308 38282
rect 35308 38236 35388 38264
rect 35256 38218 35308 38224
rect 35072 38208 35124 38214
rect 35072 38150 35124 38156
rect 34888 36916 34940 36922
rect 34888 36858 34940 36864
rect 34900 33658 34928 36858
rect 35084 36718 35112 38150
rect 35072 36712 35124 36718
rect 35072 36654 35124 36660
rect 35072 36576 35124 36582
rect 35072 36518 35124 36524
rect 35164 36576 35216 36582
rect 35164 36518 35216 36524
rect 35084 35290 35112 36518
rect 35072 35284 35124 35290
rect 35072 35226 35124 35232
rect 34980 35080 35032 35086
rect 34980 35022 35032 35028
rect 34992 34678 35020 35022
rect 34980 34672 35032 34678
rect 34980 34614 35032 34620
rect 34888 33652 34940 33658
rect 34888 33594 34940 33600
rect 34992 33590 35020 34614
rect 34980 33584 35032 33590
rect 34980 33526 35032 33532
rect 34992 32774 35020 33526
rect 34980 32768 35032 32774
rect 34980 32710 35032 32716
rect 34992 31822 35020 32710
rect 35176 32434 35204 36518
rect 35256 35692 35308 35698
rect 35256 35634 35308 35640
rect 35072 32428 35124 32434
rect 35072 32370 35124 32376
rect 35164 32428 35216 32434
rect 35164 32370 35216 32376
rect 35084 31958 35112 32370
rect 35072 31952 35124 31958
rect 35072 31894 35124 31900
rect 34980 31816 35032 31822
rect 34980 31758 35032 31764
rect 34794 31512 34850 31521
rect 34794 31447 34850 31456
rect 34992 30734 35020 31758
rect 34796 30728 34848 30734
rect 34796 30670 34848 30676
rect 34980 30728 35032 30734
rect 34980 30670 35032 30676
rect 34808 30598 34836 30670
rect 34796 30592 34848 30598
rect 34992 30569 35020 30670
rect 34796 30534 34848 30540
rect 34978 30560 35034 30569
rect 34704 29844 34756 29850
rect 34704 29786 34756 29792
rect 34704 29708 34756 29714
rect 34704 29650 34756 29656
rect 34716 25974 34744 29650
rect 34808 29238 34836 30534
rect 34978 30495 35034 30504
rect 35164 30048 35216 30054
rect 35164 29990 35216 29996
rect 34796 29232 34848 29238
rect 34796 29174 34848 29180
rect 34808 28150 34836 29174
rect 35176 28490 35204 29990
rect 35268 29782 35296 35634
rect 35360 34066 35388 38236
rect 35452 37346 35480 38966
rect 35452 37318 35572 37346
rect 35544 36242 35572 37318
rect 35728 36242 35756 40870
rect 35912 40186 35940 41386
rect 35900 40180 35952 40186
rect 35900 40122 35952 40128
rect 35900 39568 35952 39574
rect 35898 39536 35900 39545
rect 35952 39536 35954 39545
rect 35898 39471 35954 39480
rect 36004 39098 36032 44950
rect 36556 44402 36584 53926
rect 36544 44396 36596 44402
rect 36544 44338 36596 44344
rect 36556 44305 36584 44338
rect 36912 44328 36964 44334
rect 36542 44296 36598 44305
rect 36912 44270 36964 44276
rect 36542 44231 36598 44240
rect 36176 44192 36228 44198
rect 36176 44134 36228 44140
rect 35992 39092 36044 39098
rect 35992 39034 36044 39040
rect 36084 39024 36136 39030
rect 36084 38966 36136 38972
rect 35808 38412 35860 38418
rect 35808 38354 35860 38360
rect 35820 36786 35848 38354
rect 35808 36780 35860 36786
rect 35808 36722 35860 36728
rect 35532 36236 35584 36242
rect 35532 36178 35584 36184
rect 35716 36236 35768 36242
rect 35716 36178 35768 36184
rect 35820 35086 35848 36722
rect 35808 35080 35860 35086
rect 35808 35022 35860 35028
rect 35992 34196 36044 34202
rect 35992 34138 36044 34144
rect 35348 34060 35400 34066
rect 35348 34002 35400 34008
rect 35900 33312 35952 33318
rect 35900 33254 35952 33260
rect 35912 32774 35940 33254
rect 35900 32768 35952 32774
rect 35900 32710 35952 32716
rect 35912 32026 35940 32710
rect 35900 32020 35952 32026
rect 35900 31962 35952 31968
rect 36004 31929 36032 34138
rect 36096 32366 36124 38966
rect 36188 38962 36216 44134
rect 36924 42770 36952 44270
rect 37200 43722 37228 53926
rect 37660 44402 37688 53926
rect 37648 44396 37700 44402
rect 37648 44338 37700 44344
rect 37660 44305 37688 44338
rect 37646 44296 37702 44305
rect 37646 44231 37702 44240
rect 37752 43858 37780 54266
rect 37844 53582 37872 55186
rect 37950 54428 38258 54437
rect 37950 54426 37956 54428
rect 38012 54426 38036 54428
rect 38092 54426 38116 54428
rect 38172 54426 38196 54428
rect 38252 54426 38258 54428
rect 38012 54374 38014 54426
rect 38194 54374 38196 54426
rect 37950 54372 37956 54374
rect 38012 54372 38036 54374
rect 38092 54372 38116 54374
rect 38172 54372 38196 54374
rect 38252 54372 38258 54374
rect 37950 54363 38258 54372
rect 38672 54194 38700 56200
rect 39408 54194 39436 56200
rect 40144 54194 40172 56200
rect 40880 54194 40908 56200
rect 38660 54188 38712 54194
rect 38660 54130 38712 54136
rect 39396 54188 39448 54194
rect 39396 54130 39448 54136
rect 40132 54188 40184 54194
rect 40132 54130 40184 54136
rect 40868 54188 40920 54194
rect 40868 54130 40920 54136
rect 40316 54052 40368 54058
rect 40316 53994 40368 54000
rect 38936 53984 38988 53990
rect 38936 53926 38988 53932
rect 37832 53576 37884 53582
rect 37832 53518 37884 53524
rect 37832 53440 37884 53446
rect 37832 53382 37884 53388
rect 37844 44538 37872 53382
rect 37950 53340 38258 53349
rect 37950 53338 37956 53340
rect 38012 53338 38036 53340
rect 38092 53338 38116 53340
rect 38172 53338 38196 53340
rect 38252 53338 38258 53340
rect 38012 53286 38014 53338
rect 38194 53286 38196 53338
rect 37950 53284 37956 53286
rect 38012 53284 38036 53286
rect 38092 53284 38116 53286
rect 38172 53284 38196 53286
rect 38252 53284 38258 53286
rect 37950 53275 38258 53284
rect 37950 52252 38258 52261
rect 37950 52250 37956 52252
rect 38012 52250 38036 52252
rect 38092 52250 38116 52252
rect 38172 52250 38196 52252
rect 38252 52250 38258 52252
rect 38012 52198 38014 52250
rect 38194 52198 38196 52250
rect 37950 52196 37956 52198
rect 38012 52196 38036 52198
rect 38092 52196 38116 52198
rect 38172 52196 38196 52198
rect 38252 52196 38258 52198
rect 37950 52187 38258 52196
rect 37950 51164 38258 51173
rect 37950 51162 37956 51164
rect 38012 51162 38036 51164
rect 38092 51162 38116 51164
rect 38172 51162 38196 51164
rect 38252 51162 38258 51164
rect 38012 51110 38014 51162
rect 38194 51110 38196 51162
rect 37950 51108 37956 51110
rect 38012 51108 38036 51110
rect 38092 51108 38116 51110
rect 38172 51108 38196 51110
rect 38252 51108 38258 51110
rect 37950 51099 38258 51108
rect 37950 50076 38258 50085
rect 37950 50074 37956 50076
rect 38012 50074 38036 50076
rect 38092 50074 38116 50076
rect 38172 50074 38196 50076
rect 38252 50074 38258 50076
rect 38012 50022 38014 50074
rect 38194 50022 38196 50074
rect 37950 50020 37956 50022
rect 38012 50020 38036 50022
rect 38092 50020 38116 50022
rect 38172 50020 38196 50022
rect 38252 50020 38258 50022
rect 37950 50011 38258 50020
rect 37950 48988 38258 48997
rect 37950 48986 37956 48988
rect 38012 48986 38036 48988
rect 38092 48986 38116 48988
rect 38172 48986 38196 48988
rect 38252 48986 38258 48988
rect 38012 48934 38014 48986
rect 38194 48934 38196 48986
rect 37950 48932 37956 48934
rect 38012 48932 38036 48934
rect 38092 48932 38116 48934
rect 38172 48932 38196 48934
rect 38252 48932 38258 48934
rect 37950 48923 38258 48932
rect 37950 47900 38258 47909
rect 37950 47898 37956 47900
rect 38012 47898 38036 47900
rect 38092 47898 38116 47900
rect 38172 47898 38196 47900
rect 38252 47898 38258 47900
rect 38012 47846 38014 47898
rect 38194 47846 38196 47898
rect 37950 47844 37956 47846
rect 38012 47844 38036 47846
rect 38092 47844 38116 47846
rect 38172 47844 38196 47846
rect 38252 47844 38258 47846
rect 37950 47835 38258 47844
rect 37950 46812 38258 46821
rect 37950 46810 37956 46812
rect 38012 46810 38036 46812
rect 38092 46810 38116 46812
rect 38172 46810 38196 46812
rect 38252 46810 38258 46812
rect 38012 46758 38014 46810
rect 38194 46758 38196 46810
rect 37950 46756 37956 46758
rect 38012 46756 38036 46758
rect 38092 46756 38116 46758
rect 38172 46756 38196 46758
rect 38252 46756 38258 46758
rect 37950 46747 38258 46756
rect 37950 45724 38258 45733
rect 37950 45722 37956 45724
rect 38012 45722 38036 45724
rect 38092 45722 38116 45724
rect 38172 45722 38196 45724
rect 38252 45722 38258 45724
rect 38012 45670 38014 45722
rect 38194 45670 38196 45722
rect 37950 45668 37956 45670
rect 38012 45668 38036 45670
rect 38092 45668 38116 45670
rect 38172 45668 38196 45670
rect 38252 45668 38258 45670
rect 37950 45659 38258 45668
rect 38384 44872 38436 44878
rect 38384 44814 38436 44820
rect 37950 44636 38258 44645
rect 37950 44634 37956 44636
rect 38012 44634 38036 44636
rect 38092 44634 38116 44636
rect 38172 44634 38196 44636
rect 38252 44634 38258 44636
rect 38012 44582 38014 44634
rect 38194 44582 38196 44634
rect 37950 44580 37956 44582
rect 38012 44580 38036 44582
rect 38092 44580 38116 44582
rect 38172 44580 38196 44582
rect 38252 44580 38258 44582
rect 37950 44571 38258 44580
rect 37832 44532 37884 44538
rect 37832 44474 37884 44480
rect 37740 43852 37792 43858
rect 37740 43794 37792 43800
rect 38292 43852 38344 43858
rect 38292 43794 38344 43800
rect 37188 43716 37240 43722
rect 37188 43658 37240 43664
rect 37200 43489 37228 43658
rect 37280 43648 37332 43654
rect 37280 43590 37332 43596
rect 37186 43480 37242 43489
rect 37186 43415 37242 43424
rect 36912 42764 36964 42770
rect 36912 42706 36964 42712
rect 36924 41818 36952 42706
rect 37004 42696 37056 42702
rect 37004 42638 37056 42644
rect 37016 42294 37044 42638
rect 37188 42560 37240 42566
rect 37188 42502 37240 42508
rect 37004 42288 37056 42294
rect 37004 42230 37056 42236
rect 36912 41812 36964 41818
rect 36912 41754 36964 41760
rect 36636 41540 36688 41546
rect 36636 41482 36688 41488
rect 36452 39024 36504 39030
rect 36452 38966 36504 38972
rect 36176 38956 36228 38962
rect 36176 38898 36228 38904
rect 36464 36242 36492 38966
rect 36648 38554 36676 41482
rect 37016 41478 37044 42230
rect 37004 41472 37056 41478
rect 37004 41414 37056 41420
rect 37016 41138 37044 41414
rect 37004 41132 37056 41138
rect 37004 41074 37056 41080
rect 36820 40180 36872 40186
rect 36820 40122 36872 40128
rect 36636 38548 36688 38554
rect 36636 38490 36688 38496
rect 36544 36304 36596 36310
rect 36544 36246 36596 36252
rect 36452 36236 36504 36242
rect 36452 36178 36504 36184
rect 36452 36032 36504 36038
rect 36452 35974 36504 35980
rect 36176 34944 36228 34950
rect 36176 34886 36228 34892
rect 36360 34944 36412 34950
rect 36360 34886 36412 34892
rect 36084 32360 36136 32366
rect 36084 32302 36136 32308
rect 36082 32056 36138 32065
rect 36082 31991 36138 32000
rect 35990 31920 36046 31929
rect 36096 31890 36124 31991
rect 35990 31855 36046 31864
rect 36084 31884 36136 31890
rect 35716 31816 35768 31822
rect 35716 31758 35768 31764
rect 36004 31770 36032 31855
rect 36084 31826 36136 31832
rect 35624 31748 35676 31754
rect 35624 31690 35676 31696
rect 35440 31680 35492 31686
rect 35440 31622 35492 31628
rect 35256 29776 35308 29782
rect 35256 29718 35308 29724
rect 35452 29050 35480 31622
rect 35532 31272 35584 31278
rect 35532 31214 35584 31220
rect 35544 29306 35572 31214
rect 35636 30954 35664 31690
rect 35728 31668 35756 31758
rect 36004 31742 36124 31770
rect 35728 31640 35848 31668
rect 35820 31414 35848 31640
rect 35808 31408 35860 31414
rect 35808 31350 35860 31356
rect 35990 31240 36046 31249
rect 35990 31175 36046 31184
rect 35898 30968 35954 30977
rect 35636 30926 35756 30954
rect 35728 30802 35756 30926
rect 35898 30903 35954 30912
rect 35912 30870 35940 30903
rect 36004 30870 36032 31175
rect 35900 30864 35952 30870
rect 35900 30806 35952 30812
rect 35992 30864 36044 30870
rect 35992 30806 36044 30812
rect 35716 30796 35768 30802
rect 35716 30738 35768 30744
rect 35912 30410 35940 30806
rect 35636 30382 35940 30410
rect 35532 29300 35584 29306
rect 35532 29242 35584 29248
rect 35360 29022 35480 29050
rect 35164 28484 35216 28490
rect 35164 28426 35216 28432
rect 35072 28416 35124 28422
rect 35072 28358 35124 28364
rect 35256 28416 35308 28422
rect 35256 28358 35308 28364
rect 34796 28144 34848 28150
rect 34796 28086 34848 28092
rect 34808 27554 34836 28086
rect 34808 27526 35020 27554
rect 34888 27464 34940 27470
rect 34888 27406 34940 27412
rect 34796 27328 34848 27334
rect 34796 27270 34848 27276
rect 34704 25968 34756 25974
rect 34704 25910 34756 25916
rect 34704 25832 34756 25838
rect 34704 25774 34756 25780
rect 34612 25288 34664 25294
rect 34612 25230 34664 25236
rect 34716 24750 34744 25774
rect 34704 24744 34756 24750
rect 34704 24686 34756 24692
rect 34612 24404 34664 24410
rect 34612 24346 34664 24352
rect 34440 24262 34560 24290
rect 34440 24206 34468 24262
rect 34428 24200 34480 24206
rect 34428 24142 34480 24148
rect 34518 24168 34574 24177
rect 34518 24103 34574 24112
rect 34532 24070 34560 24103
rect 34428 24064 34480 24070
rect 34428 24006 34480 24012
rect 34520 24064 34572 24070
rect 34520 24006 34572 24012
rect 34440 23866 34468 24006
rect 34428 23860 34480 23866
rect 34428 23802 34480 23808
rect 34532 23730 34560 24006
rect 34520 23724 34572 23730
rect 34520 23666 34572 23672
rect 34336 23520 34388 23526
rect 34336 23462 34388 23468
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34244 23316 34296 23322
rect 34244 23258 34296 23264
rect 34152 22704 34204 22710
rect 34152 22646 34204 22652
rect 34256 22574 34284 23258
rect 34348 23254 34376 23462
rect 34336 23248 34388 23254
rect 34336 23190 34388 23196
rect 34532 22778 34560 23462
rect 34520 22772 34572 22778
rect 34520 22714 34572 22720
rect 34244 22568 34296 22574
rect 34244 22510 34296 22516
rect 34244 22228 34296 22234
rect 34244 22170 34296 22176
rect 34060 21480 34112 21486
rect 34060 21422 34112 21428
rect 34256 21350 34284 22170
rect 34428 22160 34480 22166
rect 34428 22102 34480 22108
rect 34244 21344 34296 21350
rect 34244 21286 34296 21292
rect 34256 20398 34284 21286
rect 34244 20392 34296 20398
rect 34244 20334 34296 20340
rect 33968 19848 34020 19854
rect 33968 19790 34020 19796
rect 34336 19780 34388 19786
rect 34336 19722 34388 19728
rect 34244 18760 34296 18766
rect 34244 18702 34296 18708
rect 34152 18624 34204 18630
rect 34152 18566 34204 18572
rect 33876 18352 33928 18358
rect 33876 18294 33928 18300
rect 33784 17740 33836 17746
rect 33784 17682 33836 17688
rect 33888 17678 33916 18294
rect 33876 17672 33928 17678
rect 33876 17614 33928 17620
rect 33692 17536 33744 17542
rect 33692 17478 33744 17484
rect 33600 15428 33652 15434
rect 33600 15370 33652 15376
rect 33704 13326 33732 17478
rect 33784 14884 33836 14890
rect 33784 14826 33836 14832
rect 33692 13320 33744 13326
rect 33692 13262 33744 13268
rect 33324 3052 33376 3058
rect 33324 2994 33376 3000
rect 31668 2984 31720 2990
rect 31668 2926 31720 2932
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 31680 800 31708 2926
rect 32404 2916 32456 2922
rect 32404 2858 32456 2864
rect 32416 800 32444 2858
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33796 2446 33824 14826
rect 33968 14476 34020 14482
rect 33968 14418 34020 14424
rect 33980 13530 34008 14418
rect 33968 13524 34020 13530
rect 33968 13466 34020 13472
rect 33980 12918 34008 13466
rect 34164 13326 34192 18566
rect 34256 18358 34284 18702
rect 34244 18352 34296 18358
rect 34244 18294 34296 18300
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 34244 13184 34296 13190
rect 34244 13126 34296 13132
rect 33968 12912 34020 12918
rect 33968 12854 34020 12860
rect 33968 9444 34020 9450
rect 33968 9386 34020 9392
rect 33980 4146 34008 9386
rect 33968 4140 34020 4146
rect 33968 4082 34020 4088
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 33152 800 33180 2246
rect 33888 800 33916 4014
rect 34256 3534 34284 13126
rect 34244 3528 34296 3534
rect 34244 3470 34296 3476
rect 34348 3058 34376 19722
rect 34440 17338 34468 22102
rect 34428 17332 34480 17338
rect 34428 17274 34480 17280
rect 34440 15366 34468 17274
rect 34428 15360 34480 15366
rect 34428 15302 34480 15308
rect 34428 14544 34480 14550
rect 34428 14486 34480 14492
rect 34440 12782 34468 14486
rect 34624 14414 34652 24346
rect 34704 24132 34756 24138
rect 34704 24074 34756 24080
rect 34716 20942 34744 24074
rect 34808 21010 34836 27270
rect 34900 26382 34928 27406
rect 34992 27062 35020 27526
rect 34980 27056 35032 27062
rect 34980 26998 35032 27004
rect 34980 26784 35032 26790
rect 34980 26726 35032 26732
rect 34888 26376 34940 26382
rect 34888 26318 34940 26324
rect 34992 26314 35020 26726
rect 34980 26308 35032 26314
rect 34980 26250 35032 26256
rect 34888 26240 34940 26246
rect 34888 26182 34940 26188
rect 34900 24886 34928 26182
rect 34992 25294 35020 26250
rect 34980 25288 35032 25294
rect 34980 25230 35032 25236
rect 34888 24880 34940 24886
rect 34888 24822 34940 24828
rect 34900 24313 34928 24822
rect 34992 24614 35020 25230
rect 35084 25226 35112 28358
rect 35164 27872 35216 27878
rect 35164 27814 35216 27820
rect 35072 25220 35124 25226
rect 35072 25162 35124 25168
rect 34980 24608 35032 24614
rect 34980 24550 35032 24556
rect 34886 24304 34942 24313
rect 34992 24274 35020 24550
rect 34886 24239 34942 24248
rect 34980 24268 35032 24274
rect 34980 24210 35032 24216
rect 34992 24154 35020 24210
rect 35176 24154 35204 27814
rect 35268 27577 35296 28358
rect 35254 27568 35310 27577
rect 35360 27538 35388 29022
rect 35440 28756 35492 28762
rect 35440 28698 35492 28704
rect 35452 28422 35480 28698
rect 35440 28416 35492 28422
rect 35440 28358 35492 28364
rect 35452 27878 35480 28358
rect 35440 27872 35492 27878
rect 35440 27814 35492 27820
rect 35544 27538 35572 29242
rect 35254 27503 35310 27512
rect 35348 27532 35400 27538
rect 35348 27474 35400 27480
rect 35532 27532 35584 27538
rect 35532 27474 35584 27480
rect 35636 27418 35664 30382
rect 36096 30326 36124 31742
rect 36188 30938 36216 34886
rect 36372 34134 36400 34886
rect 36360 34128 36412 34134
rect 36360 34070 36412 34076
rect 36268 32904 36320 32910
rect 36268 32846 36320 32852
rect 36280 32434 36308 32846
rect 36268 32428 36320 32434
rect 36268 32370 36320 32376
rect 36280 31482 36308 32370
rect 36360 31952 36412 31958
rect 36360 31894 36412 31900
rect 36268 31476 36320 31482
rect 36268 31418 36320 31424
rect 36176 30932 36228 30938
rect 36176 30874 36228 30880
rect 35808 30320 35860 30326
rect 36084 30320 36136 30326
rect 35860 30268 35940 30274
rect 35808 30262 35940 30268
rect 36084 30262 36136 30268
rect 35820 30246 35940 30262
rect 35912 30138 35940 30246
rect 35912 30110 36032 30138
rect 36280 30122 36308 31418
rect 36372 31278 36400 31894
rect 36464 31278 36492 35974
rect 36556 31414 36584 36246
rect 36648 35154 36676 38490
rect 36728 36576 36780 36582
rect 36728 36518 36780 36524
rect 36740 35154 36768 36518
rect 36832 36242 36860 40122
rect 37016 39370 37044 41074
rect 37094 39536 37150 39545
rect 37094 39471 37150 39480
rect 37004 39364 37056 39370
rect 37004 39306 37056 39312
rect 37016 38282 37044 39306
rect 37108 38434 37136 39471
rect 37200 38894 37228 42502
rect 37292 39098 37320 43590
rect 37950 43548 38258 43557
rect 37950 43546 37956 43548
rect 38012 43546 38036 43548
rect 38092 43546 38116 43548
rect 38172 43546 38196 43548
rect 38252 43546 38258 43548
rect 38012 43494 38014 43546
rect 38194 43494 38196 43546
rect 37950 43492 37956 43494
rect 38012 43492 38036 43494
rect 38092 43492 38116 43494
rect 38172 43492 38196 43494
rect 38252 43492 38258 43494
rect 37950 43483 38258 43492
rect 37950 42460 38258 42469
rect 37950 42458 37956 42460
rect 38012 42458 38036 42460
rect 38092 42458 38116 42460
rect 38172 42458 38196 42460
rect 38252 42458 38258 42460
rect 38012 42406 38014 42458
rect 38194 42406 38196 42458
rect 37950 42404 37956 42406
rect 38012 42404 38036 42406
rect 38092 42404 38116 42406
rect 38172 42404 38196 42406
rect 38252 42404 38258 42406
rect 37950 42395 38258 42404
rect 38304 42362 38332 43794
rect 38292 42356 38344 42362
rect 38292 42298 38344 42304
rect 37832 42152 37884 42158
rect 37832 42094 37884 42100
rect 37844 41682 37872 42094
rect 37832 41676 37884 41682
rect 37832 41618 37884 41624
rect 37844 41138 37872 41618
rect 37950 41372 38258 41381
rect 37950 41370 37956 41372
rect 38012 41370 38036 41372
rect 38092 41370 38116 41372
rect 38172 41370 38196 41372
rect 38252 41370 38258 41372
rect 38012 41318 38014 41370
rect 38194 41318 38196 41370
rect 37950 41316 37956 41318
rect 38012 41316 38036 41318
rect 38092 41316 38116 41318
rect 38172 41316 38196 41318
rect 38252 41316 38258 41318
rect 37950 41307 38258 41316
rect 37832 41132 37884 41138
rect 37832 41074 37884 41080
rect 37648 40452 37700 40458
rect 37648 40394 37700 40400
rect 37372 40384 37424 40390
rect 37372 40326 37424 40332
rect 37280 39092 37332 39098
rect 37280 39034 37332 39040
rect 37280 38956 37332 38962
rect 37280 38898 37332 38904
rect 37188 38888 37240 38894
rect 37188 38830 37240 38836
rect 37108 38406 37228 38434
rect 37004 38276 37056 38282
rect 37004 38218 37056 38224
rect 37096 38276 37148 38282
rect 37096 38218 37148 38224
rect 37108 37942 37136 38218
rect 37096 37936 37148 37942
rect 37096 37878 37148 37884
rect 37096 37256 37148 37262
rect 37096 37198 37148 37204
rect 36912 37120 36964 37126
rect 36912 37062 36964 37068
rect 36924 36582 36952 37062
rect 36912 36576 36964 36582
rect 36912 36518 36964 36524
rect 36820 36236 36872 36242
rect 36820 36178 36872 36184
rect 37108 36106 37136 37198
rect 37096 36100 37148 36106
rect 37096 36042 37148 36048
rect 36820 35692 36872 35698
rect 36820 35634 36872 35640
rect 36832 35222 36860 35634
rect 36820 35216 36872 35222
rect 36820 35158 36872 35164
rect 36636 35148 36688 35154
rect 36636 35090 36688 35096
rect 36728 35148 36780 35154
rect 36728 35090 36780 35096
rect 37096 34536 37148 34542
rect 37096 34478 37148 34484
rect 36912 33448 36964 33454
rect 36912 33390 36964 33396
rect 37002 33416 37058 33425
rect 36924 33289 36952 33390
rect 37002 33351 37004 33360
rect 37056 33351 37058 33360
rect 37004 33322 37056 33328
rect 36910 33280 36966 33289
rect 36910 33215 36966 33224
rect 36912 33108 36964 33114
rect 36912 33050 36964 33056
rect 36634 32056 36690 32065
rect 36634 31991 36690 32000
rect 36544 31408 36596 31414
rect 36544 31350 36596 31356
rect 36360 31272 36412 31278
rect 36360 31214 36412 31220
rect 36452 31272 36504 31278
rect 36452 31214 36504 31220
rect 36544 30864 36596 30870
rect 36544 30806 36596 30812
rect 36556 30598 36584 30806
rect 36544 30592 36596 30598
rect 36544 30534 36596 30540
rect 35900 29504 35952 29510
rect 35900 29446 35952 29452
rect 35808 29028 35860 29034
rect 35808 28970 35860 28976
rect 35820 28626 35848 28970
rect 35808 28620 35860 28626
rect 35808 28562 35860 28568
rect 34900 24126 35020 24154
rect 35084 24126 35204 24154
rect 35360 27390 35664 27418
rect 34796 21004 34848 21010
rect 34796 20946 34848 20952
rect 34704 20936 34756 20942
rect 34704 20878 34756 20884
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34808 18222 34836 18362
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34900 18086 34928 24126
rect 35084 22094 35112 24126
rect 35164 24064 35216 24070
rect 35164 24006 35216 24012
rect 35176 23662 35204 24006
rect 35164 23656 35216 23662
rect 35164 23598 35216 23604
rect 35176 23050 35204 23598
rect 35164 23044 35216 23050
rect 35164 22986 35216 22992
rect 35360 22094 35388 27390
rect 35820 27010 35848 28562
rect 35912 28218 35940 29446
rect 35900 28212 35952 28218
rect 35900 28154 35952 28160
rect 36004 28098 36032 30110
rect 36268 30116 36320 30122
rect 36268 30058 36320 30064
rect 36176 30048 36228 30054
rect 36176 29990 36228 29996
rect 36084 28416 36136 28422
rect 36084 28358 36136 28364
rect 35912 28070 36032 28098
rect 35912 27334 35940 28070
rect 35992 27872 36044 27878
rect 35992 27814 36044 27820
rect 35900 27328 35952 27334
rect 35900 27270 35952 27276
rect 35728 26982 35848 27010
rect 35532 26580 35584 26586
rect 35532 26522 35584 26528
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 34992 22066 35112 22094
rect 35176 22066 35388 22094
rect 34992 20330 35020 22066
rect 35072 21344 35124 21350
rect 35072 21286 35124 21292
rect 35084 21146 35112 21286
rect 35072 21140 35124 21146
rect 35072 21082 35124 21088
rect 34980 20324 35032 20330
rect 34980 20266 35032 20272
rect 34980 19712 35032 19718
rect 34980 19654 35032 19660
rect 34992 18970 35020 19654
rect 34980 18964 35032 18970
rect 34980 18906 35032 18912
rect 34888 18080 34940 18086
rect 34888 18022 34940 18028
rect 34900 16658 34928 18022
rect 34888 16652 34940 16658
rect 34888 16594 34940 16600
rect 34612 14408 34664 14414
rect 34612 14350 34664 14356
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34808 13394 34836 14010
rect 34796 13388 34848 13394
rect 34796 13330 34848 13336
rect 34900 12986 34928 16594
rect 34888 12980 34940 12986
rect 34888 12922 34940 12928
rect 34428 12776 34480 12782
rect 34428 12718 34480 12724
rect 34992 9654 35020 18906
rect 35176 18630 35204 22066
rect 35256 21956 35308 21962
rect 35256 21898 35308 21904
rect 35268 21554 35296 21898
rect 35256 21548 35308 21554
rect 35256 21490 35308 21496
rect 35348 19916 35400 19922
rect 35348 19858 35400 19864
rect 35360 19378 35388 19858
rect 35452 19854 35480 24550
rect 35544 22982 35572 26522
rect 35624 25356 35676 25362
rect 35624 25298 35676 25304
rect 35636 24070 35664 25298
rect 35728 24274 35756 26982
rect 35808 26852 35860 26858
rect 35808 26794 35860 26800
rect 35820 25974 35848 26794
rect 36004 26450 36032 27814
rect 36096 27470 36124 28358
rect 36084 27464 36136 27470
rect 36084 27406 36136 27412
rect 36084 27328 36136 27334
rect 36084 27270 36136 27276
rect 36096 26790 36124 27270
rect 36084 26784 36136 26790
rect 36084 26726 36136 26732
rect 35992 26444 36044 26450
rect 35992 26386 36044 26392
rect 35808 25968 35860 25974
rect 35808 25910 35860 25916
rect 36096 25838 36124 26726
rect 36084 25832 36136 25838
rect 36084 25774 36136 25780
rect 36188 25430 36216 29990
rect 36280 29714 36308 30058
rect 36648 30002 36676 31991
rect 36924 31754 36952 33050
rect 36832 31726 36952 31754
rect 36726 30424 36782 30433
rect 36726 30359 36782 30368
rect 36372 29974 36676 30002
rect 36268 29708 36320 29714
rect 36268 29650 36320 29656
rect 36372 29594 36400 29974
rect 36452 29844 36504 29850
rect 36452 29786 36504 29792
rect 36280 29566 36400 29594
rect 36280 29510 36308 29566
rect 36268 29504 36320 29510
rect 36268 29446 36320 29452
rect 36280 28966 36308 29446
rect 36268 28960 36320 28966
rect 36268 28902 36320 28908
rect 36360 28960 36412 28966
rect 36360 28902 36412 28908
rect 36280 28626 36308 28902
rect 36268 28620 36320 28626
rect 36268 28562 36320 28568
rect 36372 28558 36400 28902
rect 36360 28552 36412 28558
rect 36360 28494 36412 28500
rect 36176 25424 36228 25430
rect 36176 25366 36228 25372
rect 36176 24880 36228 24886
rect 36176 24822 36228 24828
rect 35716 24268 35768 24274
rect 35716 24210 35768 24216
rect 35716 24132 35768 24138
rect 35716 24074 35768 24080
rect 35624 24064 35676 24070
rect 35624 24006 35676 24012
rect 35728 24018 35756 24074
rect 35728 23990 35940 24018
rect 35912 23050 35940 23990
rect 35900 23044 35952 23050
rect 35900 22986 35952 22992
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35912 22094 35940 22986
rect 35912 22066 36124 22094
rect 36096 21962 36124 22066
rect 36084 21956 36136 21962
rect 36084 21898 36136 21904
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 36096 19446 36124 21898
rect 36084 19440 36136 19446
rect 36084 19382 36136 19388
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 36096 18766 36124 19382
rect 36188 18766 36216 24822
rect 36464 22094 36492 29786
rect 36636 29572 36688 29578
rect 36636 29514 36688 29520
rect 36544 28416 36596 28422
rect 36544 28358 36596 28364
rect 36556 28218 36584 28358
rect 36544 28212 36596 28218
rect 36544 28154 36596 28160
rect 36544 25152 36596 25158
rect 36544 25094 36596 25100
rect 36556 24954 36584 25094
rect 36544 24948 36596 24954
rect 36544 24890 36596 24896
rect 36648 24818 36676 29514
rect 36740 24886 36768 30359
rect 36832 28694 36860 31726
rect 37108 31686 37136 34478
rect 37096 31680 37148 31686
rect 37096 31622 37148 31628
rect 37004 31136 37056 31142
rect 37004 31078 37056 31084
rect 37016 30802 37044 31078
rect 36912 30796 36964 30802
rect 36912 30738 36964 30744
rect 37004 30796 37056 30802
rect 37004 30738 37056 30744
rect 36924 30394 36952 30738
rect 37096 30592 37148 30598
rect 37096 30534 37148 30540
rect 36912 30388 36964 30394
rect 36912 30330 36964 30336
rect 36820 28688 36872 28694
rect 36820 28630 36872 28636
rect 36818 28520 36874 28529
rect 36818 28455 36874 28464
rect 36832 28150 36860 28455
rect 36820 28144 36872 28150
rect 36820 28086 36872 28092
rect 36832 25786 36860 28086
rect 37108 27130 37136 30534
rect 37200 30258 37228 38406
rect 37292 37126 37320 38898
rect 37280 37120 37332 37126
rect 37280 37062 37332 37068
rect 37384 36922 37412 40326
rect 37556 39500 37608 39506
rect 37556 39442 37608 39448
rect 37464 38752 37516 38758
rect 37464 38694 37516 38700
rect 37372 36916 37424 36922
rect 37372 36858 37424 36864
rect 37372 36712 37424 36718
rect 37372 36654 37424 36660
rect 37384 36378 37412 36654
rect 37372 36372 37424 36378
rect 37372 36314 37424 36320
rect 37476 35086 37504 38694
rect 37568 37330 37596 39442
rect 37660 37754 37688 40394
rect 37844 40050 37872 41074
rect 37950 40284 38258 40293
rect 37950 40282 37956 40284
rect 38012 40282 38036 40284
rect 38092 40282 38116 40284
rect 38172 40282 38196 40284
rect 38252 40282 38258 40284
rect 38012 40230 38014 40282
rect 38194 40230 38196 40282
rect 37950 40228 37956 40230
rect 38012 40228 38036 40230
rect 38092 40228 38116 40230
rect 38172 40228 38196 40230
rect 38252 40228 38258 40230
rect 37950 40219 38258 40228
rect 37832 40044 37884 40050
rect 37832 39986 37884 39992
rect 38304 39506 38332 42298
rect 38396 40390 38424 44814
rect 38660 44328 38712 44334
rect 38660 44270 38712 44276
rect 38672 41414 38700 44270
rect 38752 44192 38804 44198
rect 38752 44134 38804 44140
rect 38488 41386 38700 41414
rect 38488 41070 38516 41386
rect 38476 41064 38528 41070
rect 38476 41006 38528 41012
rect 38384 40384 38436 40390
rect 38384 40326 38436 40332
rect 38384 39568 38436 39574
rect 38384 39510 38436 39516
rect 38292 39500 38344 39506
rect 38292 39442 38344 39448
rect 37740 39296 37792 39302
rect 37740 39238 37792 39244
rect 37752 38894 37780 39238
rect 37950 39196 38258 39205
rect 37950 39194 37956 39196
rect 38012 39194 38036 39196
rect 38092 39194 38116 39196
rect 38172 39194 38196 39196
rect 38252 39194 38258 39196
rect 38012 39142 38014 39194
rect 38194 39142 38196 39194
rect 37950 39140 37956 39142
rect 38012 39140 38036 39142
rect 38092 39140 38116 39142
rect 38172 39140 38196 39142
rect 38252 39140 38258 39142
rect 37950 39131 38258 39140
rect 38292 39024 38344 39030
rect 38292 38966 38344 38972
rect 37740 38888 37792 38894
rect 37740 38830 37792 38836
rect 37832 38820 37884 38826
rect 37832 38762 37884 38768
rect 37660 37726 37780 37754
rect 37648 37664 37700 37670
rect 37648 37606 37700 37612
rect 37556 37324 37608 37330
rect 37556 37266 37608 37272
rect 37556 37188 37608 37194
rect 37556 37130 37608 37136
rect 37568 36106 37596 37130
rect 37660 36378 37688 37606
rect 37648 36372 37700 36378
rect 37648 36314 37700 36320
rect 37752 36174 37780 37726
rect 37740 36168 37792 36174
rect 37740 36110 37792 36116
rect 37556 36100 37608 36106
rect 37556 36042 37608 36048
rect 37648 35692 37700 35698
rect 37648 35634 37700 35640
rect 37464 35080 37516 35086
rect 37464 35022 37516 35028
rect 37660 34678 37688 35634
rect 37648 34672 37700 34678
rect 37648 34614 37700 34620
rect 37280 34604 37332 34610
rect 37280 34546 37332 34552
rect 37292 32978 37320 34546
rect 37752 34474 37780 36110
rect 37844 35630 37872 38762
rect 38304 38418 38332 38966
rect 38292 38412 38344 38418
rect 38292 38354 38344 38360
rect 37950 38108 38258 38117
rect 37950 38106 37956 38108
rect 38012 38106 38036 38108
rect 38092 38106 38116 38108
rect 38172 38106 38196 38108
rect 38252 38106 38258 38108
rect 38012 38054 38014 38106
rect 38194 38054 38196 38106
rect 37950 38052 37956 38054
rect 38012 38052 38036 38054
rect 38092 38052 38116 38054
rect 38172 38052 38196 38054
rect 38252 38052 38258 38054
rect 37950 38043 38258 38052
rect 38108 37392 38160 37398
rect 38108 37334 38160 37340
rect 38120 37233 38148 37334
rect 38106 37224 38162 37233
rect 38106 37159 38162 37168
rect 38120 37126 38148 37159
rect 38108 37120 38160 37126
rect 38108 37062 38160 37068
rect 37950 37020 38258 37029
rect 37950 37018 37956 37020
rect 38012 37018 38036 37020
rect 38092 37018 38116 37020
rect 38172 37018 38196 37020
rect 38252 37018 38258 37020
rect 38012 36966 38014 37018
rect 38194 36966 38196 37018
rect 37950 36964 37956 36966
rect 38012 36964 38036 36966
rect 38092 36964 38116 36966
rect 38172 36964 38196 36966
rect 38252 36964 38258 36966
rect 37950 36955 38258 36964
rect 38016 36576 38068 36582
rect 38016 36518 38068 36524
rect 38028 36242 38056 36518
rect 38016 36236 38068 36242
rect 38016 36178 38068 36184
rect 37950 35932 38258 35941
rect 37950 35930 37956 35932
rect 38012 35930 38036 35932
rect 38092 35930 38116 35932
rect 38172 35930 38196 35932
rect 38252 35930 38258 35932
rect 38012 35878 38014 35930
rect 38194 35878 38196 35930
rect 37950 35876 37956 35878
rect 38012 35876 38036 35878
rect 38092 35876 38116 35878
rect 38172 35876 38196 35878
rect 38252 35876 38258 35878
rect 37950 35867 38258 35876
rect 38304 35714 38332 38354
rect 38396 36281 38424 39510
rect 38488 38826 38516 41006
rect 38764 40594 38792 44134
rect 38948 43314 38976 53926
rect 40132 48000 40184 48006
rect 40132 47942 40184 47948
rect 38936 43308 38988 43314
rect 38936 43250 38988 43256
rect 39764 43308 39816 43314
rect 39764 43250 39816 43256
rect 39580 42288 39632 42294
rect 39580 42230 39632 42236
rect 39304 42152 39356 42158
rect 39304 42094 39356 42100
rect 38752 40588 38804 40594
rect 38752 40530 38804 40536
rect 38844 40520 38896 40526
rect 38844 40462 38896 40468
rect 38752 40384 38804 40390
rect 38752 40326 38804 40332
rect 38568 40044 38620 40050
rect 38568 39986 38620 39992
rect 38580 39030 38608 39986
rect 38660 39636 38712 39642
rect 38660 39578 38712 39584
rect 38568 39024 38620 39030
rect 38568 38966 38620 38972
rect 38476 38820 38528 38826
rect 38476 38762 38528 38768
rect 38476 38276 38528 38282
rect 38476 38218 38528 38224
rect 38488 37806 38516 38218
rect 38476 37800 38528 37806
rect 38476 37742 38528 37748
rect 38488 36718 38516 37742
rect 38568 37392 38620 37398
rect 38568 37334 38620 37340
rect 38580 37194 38608 37334
rect 38568 37188 38620 37194
rect 38568 37130 38620 37136
rect 38476 36712 38528 36718
rect 38476 36654 38528 36660
rect 38382 36272 38438 36281
rect 38382 36207 38438 36216
rect 38396 35737 38424 36207
rect 38488 35766 38516 36654
rect 38568 36644 38620 36650
rect 38568 36586 38620 36592
rect 38476 35760 38528 35766
rect 38212 35686 38332 35714
rect 38382 35728 38438 35737
rect 37832 35624 37884 35630
rect 37832 35566 37884 35572
rect 38212 35442 38240 35686
rect 38476 35702 38528 35708
rect 38382 35663 38438 35672
rect 38384 35624 38436 35630
rect 37844 35414 38240 35442
rect 38304 35572 38384 35578
rect 38580 35578 38608 36586
rect 38304 35566 38436 35572
rect 38304 35550 38424 35566
rect 38488 35550 38608 35578
rect 37740 34468 37792 34474
rect 37740 34410 37792 34416
rect 37844 34354 37872 35414
rect 37950 34844 38258 34853
rect 37950 34842 37956 34844
rect 38012 34842 38036 34844
rect 38092 34842 38116 34844
rect 38172 34842 38196 34844
rect 38252 34842 38258 34844
rect 38012 34790 38014 34842
rect 38194 34790 38196 34842
rect 37950 34788 37956 34790
rect 38012 34788 38036 34790
rect 38092 34788 38116 34790
rect 38172 34788 38196 34790
rect 38252 34788 38258 34790
rect 37950 34779 38258 34788
rect 37660 34326 37872 34354
rect 37372 34128 37424 34134
rect 37372 34070 37424 34076
rect 37280 32972 37332 32978
rect 37280 32914 37332 32920
rect 37280 32836 37332 32842
rect 37280 32778 37332 32784
rect 37292 31890 37320 32778
rect 37280 31884 37332 31890
rect 37280 31826 37332 31832
rect 37384 31754 37412 34070
rect 37464 33992 37516 33998
rect 37464 33934 37516 33940
rect 37476 33862 37504 33934
rect 37464 33856 37516 33862
rect 37464 33798 37516 33804
rect 37464 33584 37516 33590
rect 37464 33526 37516 33532
rect 37476 33386 37504 33526
rect 37464 33380 37516 33386
rect 37464 33322 37516 33328
rect 37462 33280 37518 33289
rect 37462 33215 37518 33224
rect 37476 31890 37504 33215
rect 37556 32972 37608 32978
rect 37556 32914 37608 32920
rect 37464 31884 37516 31890
rect 37464 31826 37516 31832
rect 37384 31726 37504 31754
rect 37372 31680 37424 31686
rect 37372 31622 37424 31628
rect 37278 30560 37334 30569
rect 37278 30495 37334 30504
rect 37188 30252 37240 30258
rect 37188 30194 37240 30200
rect 37292 29578 37320 30495
rect 37280 29572 37332 29578
rect 37280 29514 37332 29520
rect 37292 29102 37320 29514
rect 37280 29096 37332 29102
rect 37280 29038 37332 29044
rect 37280 28416 37332 28422
rect 37280 28358 37332 28364
rect 37188 27872 37240 27878
rect 37188 27814 37240 27820
rect 37200 27402 37228 27814
rect 37188 27396 37240 27402
rect 37188 27338 37240 27344
rect 37096 27124 37148 27130
rect 37096 27066 37148 27072
rect 36832 25758 37044 25786
rect 36820 25696 36872 25702
rect 36820 25638 36872 25644
rect 36912 25696 36964 25702
rect 36912 25638 36964 25644
rect 36832 25362 36860 25638
rect 36820 25356 36872 25362
rect 36820 25298 36872 25304
rect 36924 25226 36952 25638
rect 36912 25220 36964 25226
rect 36912 25162 36964 25168
rect 37016 25106 37044 25758
rect 36832 25078 37044 25106
rect 36728 24880 36780 24886
rect 36728 24822 36780 24828
rect 36636 24812 36688 24818
rect 36636 24754 36688 24760
rect 36372 22066 36492 22094
rect 36372 19854 36400 22066
rect 36832 21418 36860 25078
rect 37108 23866 37136 27066
rect 37292 24818 37320 28358
rect 37384 27169 37412 31622
rect 37476 30394 37504 31726
rect 37568 31385 37596 32914
rect 37660 32502 37688 34326
rect 37740 33856 37792 33862
rect 37740 33798 37792 33804
rect 37752 32570 37780 33798
rect 37950 33756 38258 33765
rect 37950 33754 37956 33756
rect 38012 33754 38036 33756
rect 38092 33754 38116 33756
rect 38172 33754 38196 33756
rect 38252 33754 38258 33756
rect 38012 33702 38014 33754
rect 38194 33702 38196 33754
rect 37950 33700 37956 33702
rect 38012 33700 38036 33702
rect 38092 33700 38116 33702
rect 38172 33700 38196 33702
rect 38252 33700 38258 33702
rect 37950 33691 38258 33700
rect 37830 33552 37886 33561
rect 37830 33487 37832 33496
rect 37884 33487 37886 33496
rect 37832 33458 37884 33464
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 37832 32836 37884 32842
rect 37832 32778 37884 32784
rect 37740 32564 37792 32570
rect 37740 32506 37792 32512
rect 37648 32496 37700 32502
rect 37648 32438 37700 32444
rect 37844 32230 37872 32778
rect 38304 32774 38332 35550
rect 38488 34066 38516 35550
rect 38672 35154 38700 39578
rect 38764 39506 38792 40326
rect 38856 40118 38884 40462
rect 39212 40452 39264 40458
rect 39212 40394 39264 40400
rect 39120 40384 39172 40390
rect 39120 40326 39172 40332
rect 38844 40112 38896 40118
rect 38896 40060 39068 40066
rect 38844 40054 39068 40060
rect 38856 40038 39068 40054
rect 38752 39500 38804 39506
rect 38752 39442 38804 39448
rect 38844 39296 38896 39302
rect 38844 39238 38896 39244
rect 38856 39098 38884 39238
rect 38844 39092 38896 39098
rect 38844 39034 38896 39040
rect 38844 38956 38896 38962
rect 38844 38898 38896 38904
rect 38856 36786 38884 38898
rect 39040 38894 39068 40038
rect 39132 39098 39160 40326
rect 39120 39092 39172 39098
rect 39120 39034 39172 39040
rect 38936 38888 38988 38894
rect 38936 38830 38988 38836
rect 39028 38888 39080 38894
rect 39028 38830 39080 38836
rect 38844 36780 38896 36786
rect 38844 36722 38896 36728
rect 38752 35828 38804 35834
rect 38752 35770 38804 35776
rect 38764 35290 38792 35770
rect 38948 35494 38976 38830
rect 39224 38554 39252 40394
rect 39316 40202 39344 42094
rect 39592 41546 39620 42230
rect 39580 41540 39632 41546
rect 39580 41482 39632 41488
rect 39592 41138 39620 41482
rect 39776 41414 39804 43250
rect 40040 42560 40092 42566
rect 40040 42502 40092 42508
rect 39856 42084 39908 42090
rect 39856 42026 39908 42032
rect 39684 41386 39804 41414
rect 39580 41132 39632 41138
rect 39580 41074 39632 41080
rect 39316 40186 39528 40202
rect 39316 40180 39540 40186
rect 39316 40174 39488 40180
rect 39316 39506 39344 40174
rect 39488 40122 39540 40128
rect 39592 40118 39620 41074
rect 39580 40112 39632 40118
rect 39580 40054 39632 40060
rect 39304 39500 39356 39506
rect 39304 39442 39356 39448
rect 39396 39364 39448 39370
rect 39396 39306 39448 39312
rect 39408 38962 39436 39306
rect 39396 38956 39448 38962
rect 39396 38898 39448 38904
rect 39212 38548 39264 38554
rect 39212 38490 39264 38496
rect 39028 38208 39080 38214
rect 39028 38150 39080 38156
rect 38936 35488 38988 35494
rect 38936 35430 38988 35436
rect 38752 35284 38804 35290
rect 38752 35226 38804 35232
rect 38660 35148 38712 35154
rect 38660 35090 38712 35096
rect 38568 34468 38620 34474
rect 38568 34410 38620 34416
rect 38580 34082 38608 34410
rect 38476 34060 38528 34066
rect 38580 34054 38700 34082
rect 38476 34002 38528 34008
rect 38292 32768 38344 32774
rect 38292 32710 38344 32716
rect 37950 32668 38258 32677
rect 37950 32666 37956 32668
rect 38012 32666 38036 32668
rect 38092 32666 38116 32668
rect 38172 32666 38196 32668
rect 38252 32666 38258 32668
rect 38012 32614 38014 32666
rect 38194 32614 38196 32666
rect 37950 32612 37956 32614
rect 38012 32612 38036 32614
rect 38092 32612 38116 32614
rect 38172 32612 38196 32614
rect 38252 32612 38258 32614
rect 37950 32603 38258 32612
rect 37924 32496 37976 32502
rect 37924 32438 37976 32444
rect 38290 32464 38346 32473
rect 37832 32224 37884 32230
rect 37832 32166 37884 32172
rect 37738 31512 37794 31521
rect 37738 31447 37794 31456
rect 37554 31376 37610 31385
rect 37752 31346 37780 31447
rect 37554 31311 37610 31320
rect 37740 31340 37792 31346
rect 37740 31282 37792 31288
rect 37556 31136 37608 31142
rect 37556 31078 37608 31084
rect 37464 30388 37516 30394
rect 37464 30330 37516 30336
rect 37464 29708 37516 29714
rect 37464 29650 37516 29656
rect 37476 28082 37504 29650
rect 37464 28076 37516 28082
rect 37464 28018 37516 28024
rect 37370 27160 37426 27169
rect 37370 27095 37426 27104
rect 37462 27024 37518 27033
rect 37462 26959 37518 26968
rect 37476 25838 37504 26959
rect 37464 25832 37516 25838
rect 37464 25774 37516 25780
rect 37464 25696 37516 25702
rect 37464 25638 37516 25644
rect 37476 25362 37504 25638
rect 37568 25498 37596 31078
rect 37740 30592 37792 30598
rect 37740 30534 37792 30540
rect 37648 29232 37700 29238
rect 37648 29174 37700 29180
rect 37660 28014 37688 29174
rect 37648 28008 37700 28014
rect 37648 27950 37700 27956
rect 37660 26234 37688 27950
rect 37752 27554 37780 30534
rect 37844 30326 37872 32166
rect 37936 31686 37964 32438
rect 38290 32399 38346 32408
rect 37924 31680 37976 31686
rect 37924 31622 37976 31628
rect 37950 31580 38258 31589
rect 37950 31578 37956 31580
rect 38012 31578 38036 31580
rect 38092 31578 38116 31580
rect 38172 31578 38196 31580
rect 38252 31578 38258 31580
rect 38012 31526 38014 31578
rect 38194 31526 38196 31578
rect 37950 31524 37956 31526
rect 38012 31524 38036 31526
rect 38092 31524 38116 31526
rect 38172 31524 38196 31526
rect 38252 31524 38258 31526
rect 37950 31515 38258 31524
rect 38200 31408 38252 31414
rect 38198 31376 38200 31385
rect 38252 31376 38254 31385
rect 38198 31311 38254 31320
rect 37950 30492 38258 30501
rect 37950 30490 37956 30492
rect 38012 30490 38036 30492
rect 38092 30490 38116 30492
rect 38172 30490 38196 30492
rect 38252 30490 38258 30492
rect 38012 30438 38014 30490
rect 38194 30438 38196 30490
rect 37950 30436 37956 30438
rect 38012 30436 38036 30438
rect 38092 30436 38116 30438
rect 38172 30436 38196 30438
rect 38252 30436 38258 30438
rect 37950 30427 38258 30436
rect 38304 30326 38332 32399
rect 38488 32026 38516 34002
rect 38672 33998 38700 34054
rect 38568 33992 38620 33998
rect 38568 33934 38620 33940
rect 38660 33992 38712 33998
rect 38660 33934 38712 33940
rect 38476 32020 38528 32026
rect 38476 31962 38528 31968
rect 38476 31884 38528 31890
rect 38476 31826 38528 31832
rect 38384 31340 38436 31346
rect 38384 31282 38436 31288
rect 38396 30394 38424 31282
rect 38488 31210 38516 31826
rect 38476 31204 38528 31210
rect 38476 31146 38528 31152
rect 38384 30388 38436 30394
rect 38384 30330 38436 30336
rect 37832 30320 37884 30326
rect 37832 30262 37884 30268
rect 38292 30320 38344 30326
rect 38292 30262 38344 30268
rect 37950 29404 38258 29413
rect 37950 29402 37956 29404
rect 38012 29402 38036 29404
rect 38092 29402 38116 29404
rect 38172 29402 38196 29404
rect 38252 29402 38258 29404
rect 38012 29350 38014 29402
rect 38194 29350 38196 29402
rect 37950 29348 37956 29350
rect 38012 29348 38036 29350
rect 38092 29348 38116 29350
rect 38172 29348 38196 29350
rect 38252 29348 38258 29350
rect 37950 29339 38258 29348
rect 37832 29096 37884 29102
rect 37832 29038 37884 29044
rect 37844 27690 37872 29038
rect 38292 28620 38344 28626
rect 38292 28562 38344 28568
rect 37950 28316 38258 28325
rect 37950 28314 37956 28316
rect 38012 28314 38036 28316
rect 38092 28314 38116 28316
rect 38172 28314 38196 28316
rect 38252 28314 38258 28316
rect 38012 28262 38014 28314
rect 38194 28262 38196 28314
rect 37950 28260 37956 28262
rect 38012 28260 38036 28262
rect 38092 28260 38116 28262
rect 38172 28260 38196 28262
rect 38252 28260 38258 28262
rect 37950 28251 38258 28260
rect 37844 27662 37964 27690
rect 37752 27526 37872 27554
rect 37740 26988 37792 26994
rect 37740 26930 37792 26936
rect 37752 26382 37780 26930
rect 37740 26376 37792 26382
rect 37740 26318 37792 26324
rect 37660 26206 37780 26234
rect 37648 25832 37700 25838
rect 37648 25774 37700 25780
rect 37556 25492 37608 25498
rect 37556 25434 37608 25440
rect 37372 25356 37424 25362
rect 37372 25298 37424 25304
rect 37464 25356 37516 25362
rect 37464 25298 37516 25304
rect 37384 25226 37412 25298
rect 37372 25220 37424 25226
rect 37372 25162 37424 25168
rect 37280 24812 37332 24818
rect 37280 24754 37332 24760
rect 37372 24132 37424 24138
rect 37372 24074 37424 24080
rect 37096 23860 37148 23866
rect 37096 23802 37148 23808
rect 37384 22642 37412 24074
rect 37660 24070 37688 25774
rect 37752 24274 37780 26206
rect 37844 25770 37872 27526
rect 37936 27402 37964 27662
rect 37924 27396 37976 27402
rect 37924 27338 37976 27344
rect 38304 27334 38332 28562
rect 38396 27946 38424 30330
rect 38488 30326 38516 31146
rect 38476 30320 38528 30326
rect 38476 30262 38528 30268
rect 38580 29782 38608 33934
rect 38764 32910 38792 35226
rect 39040 35222 39068 38150
rect 39212 37800 39264 37806
rect 39212 37742 39264 37748
rect 39224 37330 39252 37742
rect 39212 37324 39264 37330
rect 39212 37266 39264 37272
rect 39120 37256 39172 37262
rect 39118 37224 39120 37233
rect 39172 37224 39174 37233
rect 39118 37159 39174 37168
rect 39120 36848 39172 36854
rect 39120 36790 39172 36796
rect 39028 35216 39080 35222
rect 39028 35158 39080 35164
rect 38936 34944 38988 34950
rect 38936 34886 38988 34892
rect 38844 33856 38896 33862
rect 38844 33798 38896 33804
rect 38856 33318 38884 33798
rect 38844 33312 38896 33318
rect 38844 33254 38896 33260
rect 38752 32904 38804 32910
rect 38752 32846 38804 32852
rect 38752 32768 38804 32774
rect 38752 32710 38804 32716
rect 38658 31784 38714 31793
rect 38658 31719 38660 31728
rect 38712 31719 38714 31728
rect 38660 31690 38712 31696
rect 38764 30802 38792 32710
rect 38752 30796 38804 30802
rect 38752 30738 38804 30744
rect 38752 30592 38804 30598
rect 38752 30534 38804 30540
rect 38568 29776 38620 29782
rect 38568 29718 38620 29724
rect 38660 29096 38712 29102
rect 38660 29038 38712 29044
rect 38672 28218 38700 29038
rect 38660 28212 38712 28218
rect 38660 28154 38712 28160
rect 38476 28076 38528 28082
rect 38476 28018 38528 28024
rect 38660 28076 38712 28082
rect 38660 28018 38712 28024
rect 38384 27940 38436 27946
rect 38384 27882 38436 27888
rect 38292 27328 38344 27334
rect 38292 27270 38344 27276
rect 37950 27228 38258 27237
rect 37950 27226 37956 27228
rect 38012 27226 38036 27228
rect 38092 27226 38116 27228
rect 38172 27226 38196 27228
rect 38252 27226 38258 27228
rect 38012 27174 38014 27226
rect 38194 27174 38196 27226
rect 37950 27172 37956 27174
rect 38012 27172 38036 27174
rect 38092 27172 38116 27174
rect 38172 27172 38196 27174
rect 38252 27172 38258 27174
rect 37950 27163 38258 27172
rect 37950 26140 38258 26149
rect 37950 26138 37956 26140
rect 38012 26138 38036 26140
rect 38092 26138 38116 26140
rect 38172 26138 38196 26140
rect 38252 26138 38258 26140
rect 38012 26086 38014 26138
rect 38194 26086 38196 26138
rect 37950 26084 37956 26086
rect 38012 26084 38036 26086
rect 38092 26084 38116 26086
rect 38172 26084 38196 26086
rect 38252 26084 38258 26086
rect 37950 26075 38258 26084
rect 37832 25764 37884 25770
rect 37832 25706 37884 25712
rect 37740 24268 37792 24274
rect 37740 24210 37792 24216
rect 37464 24064 37516 24070
rect 37464 24006 37516 24012
rect 37648 24064 37700 24070
rect 37648 24006 37700 24012
rect 37476 23050 37504 24006
rect 37752 23798 37780 24210
rect 37844 24206 37872 25706
rect 38304 25226 38332 27270
rect 38384 26512 38436 26518
rect 38384 26454 38436 26460
rect 38292 25220 38344 25226
rect 38292 25162 38344 25168
rect 37950 25052 38258 25061
rect 37950 25050 37956 25052
rect 38012 25050 38036 25052
rect 38092 25050 38116 25052
rect 38172 25050 38196 25052
rect 38252 25050 38258 25052
rect 38012 24998 38014 25050
rect 38194 24998 38196 25050
rect 37950 24996 37956 24998
rect 38012 24996 38036 24998
rect 38092 24996 38116 24998
rect 38172 24996 38196 24998
rect 38252 24996 38258 24998
rect 37950 24987 38258 24996
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37832 24064 37884 24070
rect 37832 24006 37884 24012
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37752 23202 37780 23734
rect 37556 23180 37608 23186
rect 37556 23122 37608 23128
rect 37660 23174 37780 23202
rect 37464 23044 37516 23050
rect 37464 22986 37516 22992
rect 37568 22778 37596 23122
rect 37556 22772 37608 22778
rect 37556 22714 37608 22720
rect 37372 22636 37424 22642
rect 37372 22578 37424 22584
rect 37660 22522 37688 23174
rect 37844 22658 37872 24006
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38292 22976 38344 22982
rect 38292 22918 38344 22924
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 36912 22500 36964 22506
rect 36912 22442 36964 22448
rect 37476 22494 37688 22522
rect 37752 22630 37872 22658
rect 36820 21412 36872 21418
rect 36820 21354 36872 21360
rect 36452 20800 36504 20806
rect 36452 20742 36504 20748
rect 36360 19848 36412 19854
rect 36360 19790 36412 19796
rect 36084 18760 36136 18766
rect 36084 18702 36136 18708
rect 36176 18760 36228 18766
rect 36176 18702 36228 18708
rect 35164 18624 35216 18630
rect 35164 18566 35216 18572
rect 35072 18420 35124 18426
rect 35072 18362 35124 18368
rect 35084 15978 35112 18362
rect 36096 18358 36124 18702
rect 36084 18352 36136 18358
rect 36084 18294 36136 18300
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 35360 17134 35388 18158
rect 35900 18080 35952 18086
rect 35900 18022 35952 18028
rect 35808 17740 35860 17746
rect 35808 17682 35860 17688
rect 35348 17128 35400 17134
rect 35348 17070 35400 17076
rect 35532 17060 35584 17066
rect 35532 17002 35584 17008
rect 35544 16658 35572 17002
rect 35532 16652 35584 16658
rect 35532 16594 35584 16600
rect 35440 16516 35492 16522
rect 35440 16458 35492 16464
rect 35072 15972 35124 15978
rect 35072 15914 35124 15920
rect 35452 14482 35480 16458
rect 35440 14476 35492 14482
rect 35440 14418 35492 14424
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 34980 9648 35032 9654
rect 34980 9590 35032 9596
rect 35176 6914 35204 14282
rect 35256 13932 35308 13938
rect 35256 13874 35308 13880
rect 35268 12850 35296 13874
rect 35544 13870 35572 16594
rect 35820 15570 35848 17682
rect 35912 17610 35940 18022
rect 35900 17604 35952 17610
rect 35900 17546 35952 17552
rect 36464 16114 36492 20742
rect 36636 19236 36688 19242
rect 36636 19178 36688 19184
rect 36544 18352 36596 18358
rect 36544 18294 36596 18300
rect 36556 17610 36584 18294
rect 36544 17604 36596 17610
rect 36544 17546 36596 17552
rect 36556 17338 36584 17546
rect 36544 17332 36596 17338
rect 36544 17274 36596 17280
rect 36556 16522 36584 17274
rect 36544 16516 36596 16522
rect 36544 16458 36596 16464
rect 36452 16108 36504 16114
rect 36452 16050 36504 16056
rect 36452 15904 36504 15910
rect 36452 15846 36504 15852
rect 35808 15564 35860 15570
rect 35808 15506 35860 15512
rect 35820 14074 35848 15506
rect 35808 14068 35860 14074
rect 35808 14010 35860 14016
rect 35532 13864 35584 13870
rect 35532 13806 35584 13812
rect 35440 13728 35492 13734
rect 35440 13670 35492 13676
rect 35452 12986 35480 13670
rect 35440 12980 35492 12986
rect 35440 12922 35492 12928
rect 36176 12980 36228 12986
rect 36176 12922 36228 12928
rect 36188 12850 36216 12922
rect 35256 12844 35308 12850
rect 35256 12786 35308 12792
rect 36176 12844 36228 12850
rect 36176 12786 36228 12792
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 36280 12442 36308 12786
rect 36268 12436 36320 12442
rect 36464 12434 36492 15846
rect 36556 15434 36584 16458
rect 36648 16454 36676 19178
rect 36728 18692 36780 18698
rect 36728 18634 36780 18640
rect 36636 16448 36688 16454
rect 36636 16390 36688 16396
rect 36544 15428 36596 15434
rect 36544 15370 36596 15376
rect 36556 13258 36584 15370
rect 36648 14958 36676 16390
rect 36636 14952 36688 14958
rect 36636 14894 36688 14900
rect 36544 13252 36596 13258
rect 36544 13194 36596 13200
rect 36556 12986 36584 13194
rect 36544 12980 36596 12986
rect 36544 12922 36596 12928
rect 36544 12708 36596 12714
rect 36544 12650 36596 12656
rect 36556 12434 36584 12650
rect 36464 12406 36584 12434
rect 36268 12378 36320 12384
rect 35176 6886 35296 6914
rect 34612 3596 34664 3602
rect 34612 3538 34664 3544
rect 34336 3052 34388 3058
rect 34336 2994 34388 3000
rect 34624 800 34652 3538
rect 35268 2446 35296 6886
rect 36556 6798 36584 12406
rect 36544 6792 36596 6798
rect 36544 6734 36596 6740
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 35348 2508 35400 2514
rect 35348 2450 35400 2456
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 35360 800 35388 2450
rect 36096 800 36124 3538
rect 36740 3534 36768 18634
rect 36832 14006 36860 21354
rect 36924 20466 36952 22442
rect 37476 22098 37504 22494
rect 37464 22092 37516 22098
rect 37752 22094 37780 22630
rect 37832 22568 37884 22574
rect 37832 22510 37884 22516
rect 37464 22034 37516 22040
rect 37660 22066 37780 22094
rect 36912 20460 36964 20466
rect 36912 20402 36964 20408
rect 37188 20324 37240 20330
rect 37188 20266 37240 20272
rect 37096 17604 37148 17610
rect 37096 17546 37148 17552
rect 37108 16794 37136 17546
rect 37096 16788 37148 16794
rect 37096 16730 37148 16736
rect 37108 15570 37136 16730
rect 37096 15564 37148 15570
rect 37096 15506 37148 15512
rect 36912 14272 36964 14278
rect 36912 14214 36964 14220
rect 36820 14000 36872 14006
rect 36820 13942 36872 13948
rect 36924 13938 36952 14214
rect 36912 13932 36964 13938
rect 36912 13874 36964 13880
rect 37200 13326 37228 20266
rect 37280 19372 37332 19378
rect 37280 19314 37332 19320
rect 37292 18834 37320 19314
rect 37464 19236 37516 19242
rect 37464 19178 37516 19184
rect 37280 18828 37332 18834
rect 37280 18770 37332 18776
rect 37292 17746 37320 18770
rect 37476 18630 37504 19178
rect 37660 18816 37688 22066
rect 37844 21486 37872 22510
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37832 21480 37884 21486
rect 37832 21422 37884 21428
rect 37844 21010 37872 21422
rect 37832 21004 37884 21010
rect 37832 20946 37884 20952
rect 38304 20942 38332 22918
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38396 20806 38424 26454
rect 38488 24138 38516 28018
rect 38568 26308 38620 26314
rect 38568 26250 38620 26256
rect 38580 25974 38608 26250
rect 38672 26042 38700 28018
rect 38660 26036 38712 26042
rect 38660 25978 38712 25984
rect 38568 25968 38620 25974
rect 38568 25910 38620 25916
rect 38476 24132 38528 24138
rect 38476 24074 38528 24080
rect 38580 23730 38608 25910
rect 38660 25696 38712 25702
rect 38660 25638 38712 25644
rect 38568 23724 38620 23730
rect 38568 23666 38620 23672
rect 38580 22778 38608 23666
rect 38568 22772 38620 22778
rect 38568 22714 38620 22720
rect 38476 21548 38528 21554
rect 38580 21536 38608 22714
rect 38528 21508 38608 21536
rect 38476 21490 38528 21496
rect 38384 20800 38436 20806
rect 38384 20742 38436 20748
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 38488 19514 38516 21490
rect 38476 19508 38528 19514
rect 38476 19450 38528 19456
rect 38568 19508 38620 19514
rect 38568 19450 38620 19456
rect 37660 18788 37872 18816
rect 37372 18624 37424 18630
rect 37372 18566 37424 18572
rect 37464 18624 37516 18630
rect 37464 18566 37516 18572
rect 37384 17882 37412 18566
rect 37372 17876 37424 17882
rect 37372 17818 37424 17824
rect 37280 17740 37332 17746
rect 37280 17682 37332 17688
rect 37384 16658 37412 17818
rect 37372 16652 37424 16658
rect 37372 16594 37424 16600
rect 37476 16046 37504 18566
rect 37740 17536 37792 17542
rect 37740 17478 37792 17484
rect 37556 17264 37608 17270
rect 37556 17206 37608 17212
rect 37464 16040 37516 16046
rect 37464 15982 37516 15988
rect 37568 15094 37596 17206
rect 37752 16522 37780 17478
rect 37740 16516 37792 16522
rect 37740 16458 37792 16464
rect 37648 15904 37700 15910
rect 37648 15846 37700 15852
rect 37660 15162 37688 15846
rect 37740 15360 37792 15366
rect 37740 15302 37792 15308
rect 37648 15156 37700 15162
rect 37648 15098 37700 15104
rect 37556 15088 37608 15094
rect 37556 15030 37608 15036
rect 37372 14816 37424 14822
rect 37372 14758 37424 14764
rect 37384 13326 37412 14758
rect 37752 14482 37780 15302
rect 37740 14476 37792 14482
rect 37740 14418 37792 14424
rect 37752 13394 37780 14418
rect 37844 13938 37872 18788
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 38580 18222 38608 19450
rect 38672 18426 38700 25638
rect 38764 25158 38792 30534
rect 38856 26042 38884 33254
rect 38948 30954 38976 34886
rect 39040 32910 39068 35158
rect 39028 32904 39080 32910
rect 39028 32846 39080 32852
rect 39026 31376 39082 31385
rect 39026 31311 39028 31320
rect 39080 31311 39082 31320
rect 39028 31282 39080 31288
rect 38948 30926 39068 30954
rect 38936 30864 38988 30870
rect 38936 30806 38988 30812
rect 38948 28490 38976 30806
rect 39040 29102 39068 30926
rect 39028 29096 39080 29102
rect 39028 29038 39080 29044
rect 39132 28762 39160 36790
rect 39408 36145 39436 38898
rect 39488 38480 39540 38486
rect 39488 38422 39540 38428
rect 39394 36136 39450 36145
rect 39394 36071 39450 36080
rect 39408 35834 39436 36071
rect 39396 35828 39448 35834
rect 39396 35770 39448 35776
rect 39302 35592 39358 35601
rect 39302 35527 39358 35536
rect 39212 33516 39264 33522
rect 39212 33458 39264 33464
rect 39120 28756 39172 28762
rect 39120 28698 39172 28704
rect 39224 28694 39252 33458
rect 39316 32774 39344 35527
rect 39304 32768 39356 32774
rect 39304 32710 39356 32716
rect 39304 32292 39356 32298
rect 39304 32234 39356 32240
rect 39316 31822 39344 32234
rect 39304 31816 39356 31822
rect 39304 31758 39356 31764
rect 39500 31482 39528 38422
rect 39592 37942 39620 40054
rect 39580 37936 39632 37942
rect 39580 37878 39632 37884
rect 39592 36530 39620 37878
rect 39684 36854 39712 41386
rect 39868 38214 39896 42026
rect 39948 40928 40000 40934
rect 39948 40870 40000 40876
rect 39960 40594 39988 40870
rect 39948 40588 40000 40594
rect 39948 40530 40000 40536
rect 39948 39840 40000 39846
rect 39948 39782 40000 39788
rect 39960 39574 39988 39782
rect 39948 39568 40000 39574
rect 39948 39510 40000 39516
rect 39948 39296 40000 39302
rect 39948 39238 40000 39244
rect 39960 38894 39988 39238
rect 39948 38888 40000 38894
rect 39948 38830 40000 38836
rect 40052 38434 40080 42502
rect 40144 39982 40172 47942
rect 40328 43450 40356 53994
rect 40408 53984 40460 53990
rect 40408 53926 40460 53932
rect 41052 53984 41104 53990
rect 41052 53926 41104 53932
rect 40316 43444 40368 43450
rect 40316 43386 40368 43392
rect 40420 42566 40448 53926
rect 40684 53440 40736 53446
rect 40684 53382 40736 53388
rect 40696 44538 40724 53382
rect 40684 44532 40736 44538
rect 40684 44474 40736 44480
rect 40776 43784 40828 43790
rect 40776 43726 40828 43732
rect 40500 43240 40552 43246
rect 40500 43182 40552 43188
rect 40408 42560 40460 42566
rect 40408 42502 40460 42508
rect 40420 41721 40448 42502
rect 40406 41712 40462 41721
rect 40406 41647 40462 41656
rect 40132 39976 40184 39982
rect 40132 39918 40184 39924
rect 40144 39098 40172 39918
rect 40316 39432 40368 39438
rect 40316 39374 40368 39380
rect 40132 39092 40184 39098
rect 40132 39034 40184 39040
rect 40328 38894 40356 39374
rect 40408 39092 40460 39098
rect 40408 39034 40460 39040
rect 40316 38888 40368 38894
rect 40316 38830 40368 38836
rect 40052 38406 40264 38434
rect 40132 38276 40184 38282
rect 40132 38218 40184 38224
rect 39856 38208 39908 38214
rect 39856 38150 39908 38156
rect 40144 37942 40172 38218
rect 40132 37936 40184 37942
rect 40132 37878 40184 37884
rect 39868 37738 40172 37754
rect 39868 37732 40184 37738
rect 39868 37726 40132 37732
rect 39764 37392 39816 37398
rect 39764 37334 39816 37340
rect 39672 36848 39724 36854
rect 39672 36790 39724 36796
rect 39672 36644 39724 36650
rect 39672 36586 39724 36592
rect 39684 36530 39712 36586
rect 39592 36502 39712 36530
rect 39684 35766 39712 36502
rect 39672 35760 39724 35766
rect 39672 35702 39724 35708
rect 39684 32502 39712 35702
rect 39776 35630 39804 37334
rect 39764 35624 39816 35630
rect 39764 35566 39816 35572
rect 39868 35086 39896 37726
rect 40132 37674 40184 37680
rect 39948 37664 40000 37670
rect 39948 37606 40000 37612
rect 39960 37398 39988 37606
rect 39948 37392 40000 37398
rect 39948 37334 40000 37340
rect 40040 37392 40092 37398
rect 40092 37340 40172 37346
rect 40040 37334 40172 37340
rect 40052 37318 40172 37334
rect 39948 36848 40000 36854
rect 39948 36790 40000 36796
rect 39960 35834 39988 36790
rect 40144 36224 40172 37318
rect 40236 37262 40264 38406
rect 40316 37664 40368 37670
rect 40316 37606 40368 37612
rect 40328 37330 40356 37606
rect 40316 37324 40368 37330
rect 40316 37266 40368 37272
rect 40224 37256 40276 37262
rect 40224 37198 40276 37204
rect 40052 36196 40172 36224
rect 39948 35828 40000 35834
rect 39948 35770 40000 35776
rect 39856 35080 39908 35086
rect 39856 35022 39908 35028
rect 39960 34542 39988 35770
rect 40052 34746 40080 36196
rect 40132 36100 40184 36106
rect 40132 36042 40184 36048
rect 40144 35834 40172 36042
rect 40132 35828 40184 35834
rect 40132 35770 40184 35776
rect 40224 35760 40276 35766
rect 40224 35702 40276 35708
rect 40040 34740 40092 34746
rect 40040 34682 40092 34688
rect 39948 34536 40000 34542
rect 39948 34478 40000 34484
rect 39764 34400 39816 34406
rect 39764 34342 39816 34348
rect 39672 32496 39724 32502
rect 39672 32438 39724 32444
rect 39672 32224 39724 32230
rect 39672 32166 39724 32172
rect 39684 31686 39712 32166
rect 39776 32026 39804 34342
rect 40236 33522 40264 35702
rect 40420 35630 40448 39034
rect 40512 38418 40540 43182
rect 40684 42764 40736 42770
rect 40684 42706 40736 42712
rect 40592 42560 40644 42566
rect 40592 42502 40644 42508
rect 40500 38412 40552 38418
rect 40500 38354 40552 38360
rect 40604 36310 40632 42502
rect 40696 37398 40724 42706
rect 40788 41414 40816 43726
rect 41064 42226 41092 53926
rect 41616 53582 41644 56200
rect 42352 54262 42380 56200
rect 42340 54256 42392 54262
rect 42340 54198 42392 54204
rect 43088 54194 43116 56200
rect 43824 56114 43852 56200
rect 43916 56114 43944 56222
rect 43824 56086 43944 56114
rect 44100 54194 44128 56222
rect 44546 56200 44602 57000
rect 46754 56200 46810 57000
rect 47490 56200 47546 57000
rect 48226 56200 48282 57000
rect 48962 56200 49018 57000
rect 49698 56200 49754 57000
rect 50434 56200 50490 57000
rect 44560 54194 44588 56200
rect 43076 54188 43128 54194
rect 43076 54130 43128 54136
rect 44088 54188 44140 54194
rect 44088 54130 44140 54136
rect 44548 54188 44600 54194
rect 44548 54130 44600 54136
rect 43996 54120 44048 54126
rect 43996 54062 44048 54068
rect 43444 54052 43496 54058
rect 43444 53994 43496 54000
rect 42950 53884 43258 53893
rect 42950 53882 42956 53884
rect 43012 53882 43036 53884
rect 43092 53882 43116 53884
rect 43172 53882 43196 53884
rect 43252 53882 43258 53884
rect 43012 53830 43014 53882
rect 43194 53830 43196 53882
rect 42950 53828 42956 53830
rect 43012 53828 43036 53830
rect 43092 53828 43116 53830
rect 43172 53828 43196 53830
rect 43252 53828 43258 53830
rect 42950 53819 43258 53828
rect 41604 53576 41656 53582
rect 41604 53518 41656 53524
rect 42950 52796 43258 52805
rect 42950 52794 42956 52796
rect 43012 52794 43036 52796
rect 43092 52794 43116 52796
rect 43172 52794 43196 52796
rect 43252 52794 43258 52796
rect 43012 52742 43014 52794
rect 43194 52742 43196 52794
rect 42950 52740 42956 52742
rect 43012 52740 43036 52742
rect 43092 52740 43116 52742
rect 43172 52740 43196 52742
rect 43252 52740 43258 52742
rect 42950 52731 43258 52740
rect 42950 51708 43258 51717
rect 42950 51706 42956 51708
rect 43012 51706 43036 51708
rect 43092 51706 43116 51708
rect 43172 51706 43196 51708
rect 43252 51706 43258 51708
rect 43012 51654 43014 51706
rect 43194 51654 43196 51706
rect 42950 51652 42956 51654
rect 43012 51652 43036 51654
rect 43092 51652 43116 51654
rect 43172 51652 43196 51654
rect 43252 51652 43258 51654
rect 42950 51643 43258 51652
rect 42950 50620 43258 50629
rect 42950 50618 42956 50620
rect 43012 50618 43036 50620
rect 43092 50618 43116 50620
rect 43172 50618 43196 50620
rect 43252 50618 43258 50620
rect 43012 50566 43014 50618
rect 43194 50566 43196 50618
rect 42950 50564 42956 50566
rect 43012 50564 43036 50566
rect 43092 50564 43116 50566
rect 43172 50564 43196 50566
rect 43252 50564 43258 50566
rect 42950 50555 43258 50564
rect 42950 49532 43258 49541
rect 42950 49530 42956 49532
rect 43012 49530 43036 49532
rect 43092 49530 43116 49532
rect 43172 49530 43196 49532
rect 43252 49530 43258 49532
rect 43012 49478 43014 49530
rect 43194 49478 43196 49530
rect 42950 49476 42956 49478
rect 43012 49476 43036 49478
rect 43092 49476 43116 49478
rect 43172 49476 43196 49478
rect 43252 49476 43258 49478
rect 42950 49467 43258 49476
rect 42950 48444 43258 48453
rect 42950 48442 42956 48444
rect 43012 48442 43036 48444
rect 43092 48442 43116 48444
rect 43172 48442 43196 48444
rect 43252 48442 43258 48444
rect 43012 48390 43014 48442
rect 43194 48390 43196 48442
rect 42950 48388 42956 48390
rect 43012 48388 43036 48390
rect 43092 48388 43116 48390
rect 43172 48388 43196 48390
rect 43252 48388 43258 48390
rect 42950 48379 43258 48388
rect 42950 47356 43258 47365
rect 42950 47354 42956 47356
rect 43012 47354 43036 47356
rect 43092 47354 43116 47356
rect 43172 47354 43196 47356
rect 43252 47354 43258 47356
rect 43012 47302 43014 47354
rect 43194 47302 43196 47354
rect 42950 47300 42956 47302
rect 43012 47300 43036 47302
rect 43092 47300 43116 47302
rect 43172 47300 43196 47302
rect 43252 47300 43258 47302
rect 42950 47291 43258 47300
rect 42950 46268 43258 46277
rect 42950 46266 42956 46268
rect 43012 46266 43036 46268
rect 43092 46266 43116 46268
rect 43172 46266 43196 46268
rect 43252 46266 43258 46268
rect 43012 46214 43014 46266
rect 43194 46214 43196 46266
rect 42950 46212 42956 46214
rect 43012 46212 43036 46214
rect 43092 46212 43116 46214
rect 43172 46212 43196 46214
rect 43252 46212 43258 46214
rect 42950 46203 43258 46212
rect 42950 45180 43258 45189
rect 42950 45178 42956 45180
rect 43012 45178 43036 45180
rect 43092 45178 43116 45180
rect 43172 45178 43196 45180
rect 43252 45178 43258 45180
rect 43012 45126 43014 45178
rect 43194 45126 43196 45178
rect 42950 45124 42956 45126
rect 43012 45124 43036 45126
rect 43092 45124 43116 45126
rect 43172 45124 43196 45126
rect 43252 45124 43258 45126
rect 42950 45115 43258 45124
rect 42950 44092 43258 44101
rect 42950 44090 42956 44092
rect 43012 44090 43036 44092
rect 43092 44090 43116 44092
rect 43172 44090 43196 44092
rect 43252 44090 43258 44092
rect 43012 44038 43014 44090
rect 43194 44038 43196 44090
rect 42950 44036 42956 44038
rect 43012 44036 43036 44038
rect 43092 44036 43116 44038
rect 43172 44036 43196 44038
rect 43252 44036 43258 44038
rect 42950 44027 43258 44036
rect 41604 43240 41656 43246
rect 41604 43182 41656 43188
rect 41236 43104 41288 43110
rect 41236 43046 41288 43052
rect 41052 42220 41104 42226
rect 41052 42162 41104 42168
rect 40788 41386 41000 41414
rect 40972 38758 41000 41386
rect 41144 40112 41196 40118
rect 41144 40054 41196 40060
rect 41052 38888 41104 38894
rect 41052 38830 41104 38836
rect 40960 38752 41012 38758
rect 40960 38694 41012 38700
rect 40684 37392 40736 37398
rect 40684 37334 40736 37340
rect 40696 37194 40724 37334
rect 40684 37188 40736 37194
rect 40684 37130 40736 37136
rect 40592 36304 40644 36310
rect 40592 36246 40644 36252
rect 40604 36122 40632 36246
rect 40604 36094 40724 36122
rect 40592 36032 40644 36038
rect 40592 35974 40644 35980
rect 40408 35624 40460 35630
rect 40408 35566 40460 35572
rect 40500 34944 40552 34950
rect 40500 34886 40552 34892
rect 40512 34746 40540 34886
rect 40500 34740 40552 34746
rect 40500 34682 40552 34688
rect 40512 34610 40540 34682
rect 40500 34604 40552 34610
rect 40500 34546 40552 34552
rect 40604 34202 40632 35974
rect 40592 34196 40644 34202
rect 40592 34138 40644 34144
rect 40224 33516 40276 33522
rect 40224 33458 40276 33464
rect 40316 33448 40368 33454
rect 40316 33390 40368 33396
rect 40592 33448 40644 33454
rect 40592 33390 40644 33396
rect 40224 32768 40276 32774
rect 40224 32710 40276 32716
rect 39764 32020 39816 32026
rect 39764 31962 39816 31968
rect 39672 31680 39724 31686
rect 39672 31622 39724 31628
rect 39304 31476 39356 31482
rect 39304 31418 39356 31424
rect 39488 31476 39540 31482
rect 39488 31418 39540 31424
rect 39316 30705 39344 31418
rect 39488 30932 39540 30938
rect 39488 30874 39540 30880
rect 39396 30796 39448 30802
rect 39396 30738 39448 30744
rect 39302 30696 39358 30705
rect 39302 30631 39358 30640
rect 39212 28688 39264 28694
rect 39212 28630 39264 28636
rect 39028 28552 39080 28558
rect 39028 28494 39080 28500
rect 38936 28484 38988 28490
rect 38936 28426 38988 28432
rect 39040 28218 39068 28494
rect 39028 28212 39080 28218
rect 39028 28154 39080 28160
rect 39120 28008 39172 28014
rect 39120 27950 39172 27956
rect 39132 27674 39160 27950
rect 39120 27668 39172 27674
rect 39120 27610 39172 27616
rect 39028 26784 39080 26790
rect 39028 26726 39080 26732
rect 39040 26518 39068 26726
rect 39028 26512 39080 26518
rect 39028 26454 39080 26460
rect 39316 26042 39344 30631
rect 39408 29034 39436 30738
rect 39500 30734 39528 30874
rect 39488 30728 39540 30734
rect 39488 30670 39540 30676
rect 39776 29714 39804 31962
rect 40040 30592 40092 30598
rect 40040 30534 40092 30540
rect 39764 29708 39816 29714
rect 39764 29650 39816 29656
rect 40052 29306 40080 30534
rect 40132 30116 40184 30122
rect 40132 30058 40184 30064
rect 40040 29300 40092 29306
rect 40040 29242 40092 29248
rect 39396 29028 39448 29034
rect 39396 28970 39448 28976
rect 39488 28688 39540 28694
rect 39488 28630 39540 28636
rect 39500 28082 39528 28630
rect 39488 28076 39540 28082
rect 39488 28018 39540 28024
rect 40144 27010 40172 30058
rect 40236 28626 40264 32710
rect 40328 32570 40356 33390
rect 40604 33046 40632 33390
rect 40592 33040 40644 33046
rect 40592 32982 40644 32988
rect 40696 32978 40724 36094
rect 40776 35828 40828 35834
rect 40776 35770 40828 35776
rect 40684 32972 40736 32978
rect 40684 32914 40736 32920
rect 40788 32910 40816 35770
rect 40866 35048 40922 35057
rect 40866 34983 40922 34992
rect 40880 34950 40908 34983
rect 40868 34944 40920 34950
rect 40868 34886 40920 34892
rect 40880 34626 40908 34886
rect 40972 34746 41000 38694
rect 41064 38418 41092 38830
rect 41156 38554 41184 40054
rect 41248 40050 41276 43046
rect 41328 42220 41380 42226
rect 41328 42162 41380 42168
rect 41340 42129 41368 42162
rect 41326 42120 41382 42129
rect 41326 42055 41382 42064
rect 41236 40044 41288 40050
rect 41236 39986 41288 39992
rect 41616 39914 41644 43182
rect 42950 43004 43258 43013
rect 42950 43002 42956 43004
rect 43012 43002 43036 43004
rect 43092 43002 43116 43004
rect 43172 43002 43196 43004
rect 43252 43002 43258 43004
rect 43012 42950 43014 43002
rect 43194 42950 43196 43002
rect 42950 42948 42956 42950
rect 43012 42948 43036 42950
rect 43092 42948 43116 42950
rect 43172 42948 43196 42950
rect 43252 42948 43258 42950
rect 42950 42939 43258 42948
rect 43456 42702 43484 53994
rect 43444 42696 43496 42702
rect 43444 42638 43496 42644
rect 41880 42152 41932 42158
rect 41880 42094 41932 42100
rect 41788 39976 41840 39982
rect 41788 39918 41840 39924
rect 41604 39908 41656 39914
rect 41604 39850 41656 39856
rect 41236 39364 41288 39370
rect 41236 39306 41288 39312
rect 41248 38894 41276 39306
rect 41236 38888 41288 38894
rect 41236 38830 41288 38836
rect 41144 38548 41196 38554
rect 41144 38490 41196 38496
rect 41236 38548 41288 38554
rect 41236 38490 41288 38496
rect 41052 38412 41104 38418
rect 41052 38354 41104 38360
rect 41064 36582 41092 38354
rect 41248 38010 41276 38490
rect 41328 38480 41380 38486
rect 41328 38422 41380 38428
rect 41340 38214 41368 38422
rect 41512 38344 41564 38350
rect 41512 38286 41564 38292
rect 41328 38208 41380 38214
rect 41328 38150 41380 38156
rect 41236 38004 41288 38010
rect 41236 37946 41288 37952
rect 41328 37800 41380 37806
rect 41328 37742 41380 37748
rect 41340 36904 41368 37742
rect 41524 37330 41552 38286
rect 41512 37324 41564 37330
rect 41512 37266 41564 37272
rect 41420 37256 41472 37262
rect 41420 37198 41472 37204
rect 41248 36876 41368 36904
rect 41052 36576 41104 36582
rect 41052 36518 41104 36524
rect 40960 34740 41012 34746
rect 40960 34682 41012 34688
rect 40880 34598 41000 34626
rect 40868 34536 40920 34542
rect 40868 34478 40920 34484
rect 40880 33590 40908 34478
rect 40868 33584 40920 33590
rect 40868 33526 40920 33532
rect 40776 32904 40828 32910
rect 40776 32846 40828 32852
rect 40316 32564 40368 32570
rect 40316 32506 40368 32512
rect 40328 31890 40356 32506
rect 40972 32314 41000 34598
rect 41064 33998 41092 36518
rect 41248 34762 41276 36876
rect 41328 36780 41380 36786
rect 41328 36722 41380 36728
rect 41340 36378 41368 36722
rect 41328 36372 41380 36378
rect 41328 36314 41380 36320
rect 41432 36174 41460 37198
rect 41524 36922 41552 37266
rect 41616 37210 41644 39850
rect 41800 38758 41828 39918
rect 41788 38752 41840 38758
rect 41788 38694 41840 38700
rect 41800 38282 41828 38694
rect 41788 38276 41840 38282
rect 41788 38218 41840 38224
rect 41616 37182 41736 37210
rect 41604 37120 41656 37126
rect 41604 37062 41656 37068
rect 41616 36922 41644 37062
rect 41512 36916 41564 36922
rect 41512 36858 41564 36864
rect 41604 36916 41656 36922
rect 41604 36858 41656 36864
rect 41420 36168 41472 36174
rect 41420 36110 41472 36116
rect 41708 35894 41736 37182
rect 41800 36242 41828 38218
rect 41788 36236 41840 36242
rect 41788 36178 41840 36184
rect 41708 35866 41828 35894
rect 41696 35080 41748 35086
rect 41696 35022 41748 35028
rect 41156 34734 41276 34762
rect 41708 34746 41736 35022
rect 41696 34740 41748 34746
rect 41052 33992 41104 33998
rect 41052 33934 41104 33940
rect 41156 33454 41184 34734
rect 41696 34682 41748 34688
rect 41236 34672 41288 34678
rect 41288 34632 41552 34660
rect 41236 34614 41288 34620
rect 41420 33856 41472 33862
rect 41420 33798 41472 33804
rect 41144 33448 41196 33454
rect 41144 33390 41196 33396
rect 41236 32972 41288 32978
rect 41236 32914 41288 32920
rect 41052 32768 41104 32774
rect 41052 32710 41104 32716
rect 40880 32286 41000 32314
rect 40500 31952 40552 31958
rect 40592 31952 40644 31958
rect 40500 31894 40552 31900
rect 40590 31920 40592 31929
rect 40644 31920 40646 31929
rect 40316 31884 40368 31890
rect 40316 31826 40368 31832
rect 40408 31136 40460 31142
rect 40408 31078 40460 31084
rect 40420 30734 40448 31078
rect 40512 30802 40540 31894
rect 40590 31855 40646 31864
rect 40776 31136 40828 31142
rect 40776 31078 40828 31084
rect 40500 30796 40552 30802
rect 40500 30738 40552 30744
rect 40592 30796 40644 30802
rect 40592 30738 40644 30744
rect 40408 30728 40460 30734
rect 40408 30670 40460 30676
rect 40604 30138 40632 30738
rect 40512 30110 40632 30138
rect 40684 30184 40736 30190
rect 40684 30126 40736 30132
rect 40512 30054 40540 30110
rect 40500 30048 40552 30054
rect 40500 29990 40552 29996
rect 40316 29708 40368 29714
rect 40316 29650 40368 29656
rect 40224 28620 40276 28626
rect 40224 28562 40276 28568
rect 40224 28416 40276 28422
rect 40224 28358 40276 28364
rect 39856 26988 39908 26994
rect 39856 26930 39908 26936
rect 40052 26982 40172 27010
rect 39868 26450 39896 26930
rect 39396 26444 39448 26450
rect 39396 26386 39448 26392
rect 39856 26444 39908 26450
rect 39856 26386 39908 26392
rect 38844 26036 38896 26042
rect 38844 25978 38896 25984
rect 39304 26036 39356 26042
rect 39304 25978 39356 25984
rect 39212 25832 39264 25838
rect 39212 25774 39264 25780
rect 38752 25152 38804 25158
rect 38752 25094 38804 25100
rect 38752 23180 38804 23186
rect 38752 23122 38804 23128
rect 38764 21622 38792 23122
rect 39028 22568 39080 22574
rect 39028 22510 39080 22516
rect 39040 21622 39068 22510
rect 38752 21616 38804 21622
rect 38752 21558 38804 21564
rect 38844 21616 38896 21622
rect 38844 21558 38896 21564
rect 39028 21616 39080 21622
rect 39028 21558 39080 21564
rect 38856 21434 38884 21558
rect 38764 21406 38884 21434
rect 38764 19446 38792 21406
rect 38752 19440 38804 19446
rect 38752 19382 38804 19388
rect 38764 18698 38792 19382
rect 38752 18692 38804 18698
rect 38752 18634 38804 18640
rect 38660 18420 38712 18426
rect 38660 18362 38712 18368
rect 38764 18306 38792 18634
rect 39224 18630 39252 25774
rect 39408 23866 39436 26386
rect 39948 26376 40000 26382
rect 40052 26364 40080 26982
rect 40132 26920 40184 26926
rect 40132 26862 40184 26868
rect 40144 26586 40172 26862
rect 40132 26580 40184 26586
rect 40132 26522 40184 26528
rect 40000 26336 40080 26364
rect 39948 26318 40000 26324
rect 39488 26308 39540 26314
rect 39488 26250 39540 26256
rect 39500 25498 39528 26250
rect 40144 25906 40172 26522
rect 40132 25900 40184 25906
rect 40132 25842 40184 25848
rect 39672 25764 39724 25770
rect 39672 25706 39724 25712
rect 39580 25696 39632 25702
rect 39580 25638 39632 25644
rect 39488 25492 39540 25498
rect 39488 25434 39540 25440
rect 39500 24750 39528 25434
rect 39592 25226 39620 25638
rect 39684 25498 39712 25706
rect 39672 25492 39724 25498
rect 39672 25434 39724 25440
rect 39580 25220 39632 25226
rect 39580 25162 39632 25168
rect 39488 24744 39540 24750
rect 39488 24686 39540 24692
rect 39488 24336 39540 24342
rect 39488 24278 39540 24284
rect 39396 23860 39448 23866
rect 39396 23802 39448 23808
rect 39408 23186 39436 23802
rect 39396 23180 39448 23186
rect 39396 23122 39448 23128
rect 39500 22574 39528 24278
rect 39592 23798 39620 25162
rect 40040 25152 40092 25158
rect 40040 25094 40092 25100
rect 40052 24206 40080 25094
rect 40236 24274 40264 28358
rect 40328 27538 40356 29650
rect 40512 29578 40540 29990
rect 40696 29714 40724 30126
rect 40684 29708 40736 29714
rect 40684 29650 40736 29656
rect 40788 29646 40816 31078
rect 40880 30190 40908 32286
rect 40960 32224 41012 32230
rect 40960 32166 41012 32172
rect 40972 32026 41000 32166
rect 40960 32020 41012 32026
rect 40960 31962 41012 31968
rect 40868 30184 40920 30190
rect 40868 30126 40920 30132
rect 40776 29640 40828 29646
rect 40776 29582 40828 29588
rect 40500 29572 40552 29578
rect 40500 29514 40552 29520
rect 40512 28014 40540 29514
rect 40684 28620 40736 28626
rect 40684 28562 40736 28568
rect 40500 28008 40552 28014
rect 40500 27950 40552 27956
rect 40316 27532 40368 27538
rect 40316 27474 40368 27480
rect 40328 26994 40356 27474
rect 40590 27160 40646 27169
rect 40696 27130 40724 28562
rect 41064 28558 41092 32710
rect 41248 31754 41276 32914
rect 41328 32564 41380 32570
rect 41328 32506 41380 32512
rect 41156 31726 41276 31754
rect 41156 29322 41184 31726
rect 41236 30660 41288 30666
rect 41340 30648 41368 32506
rect 41288 30620 41368 30648
rect 41236 30602 41288 30608
rect 41248 30394 41276 30602
rect 41236 30388 41288 30394
rect 41236 30330 41288 30336
rect 41328 30116 41380 30122
rect 41328 30058 41380 30064
rect 41156 29294 41276 29322
rect 41144 29164 41196 29170
rect 41144 29106 41196 29112
rect 41052 28552 41104 28558
rect 41052 28494 41104 28500
rect 41156 27946 41184 29106
rect 41144 27940 41196 27946
rect 41144 27882 41196 27888
rect 41248 27878 41276 29294
rect 41340 29238 41368 30058
rect 41432 29510 41460 33798
rect 41524 30870 41552 34632
rect 41604 34468 41656 34474
rect 41604 34410 41656 34416
rect 41512 30864 41564 30870
rect 41512 30806 41564 30812
rect 41420 29504 41472 29510
rect 41420 29446 41472 29452
rect 41328 29232 41380 29238
rect 41328 29174 41380 29180
rect 41616 28082 41644 34410
rect 41800 32978 41828 35866
rect 41892 35766 41920 42094
rect 42340 42016 42392 42022
rect 42340 41958 42392 41964
rect 41972 37936 42024 37942
rect 41972 37878 42024 37884
rect 41880 35760 41932 35766
rect 41880 35702 41932 35708
rect 41984 33998 42012 37878
rect 42156 37664 42208 37670
rect 42156 37606 42208 37612
rect 42248 37664 42300 37670
rect 42248 37606 42300 37612
rect 42064 34128 42116 34134
rect 42064 34070 42116 34076
rect 41972 33992 42024 33998
rect 41972 33934 42024 33940
rect 41880 33856 41932 33862
rect 41880 33798 41932 33804
rect 41788 32972 41840 32978
rect 41788 32914 41840 32920
rect 41788 31680 41840 31686
rect 41788 31622 41840 31628
rect 41696 30252 41748 30258
rect 41696 30194 41748 30200
rect 41708 29578 41736 30194
rect 41696 29572 41748 29578
rect 41696 29514 41748 29520
rect 41604 28076 41656 28082
rect 41604 28018 41656 28024
rect 41236 27872 41288 27878
rect 41236 27814 41288 27820
rect 40776 27668 40828 27674
rect 40776 27610 40828 27616
rect 40590 27095 40592 27104
rect 40644 27095 40646 27104
rect 40684 27124 40736 27130
rect 40592 27066 40644 27072
rect 40684 27066 40736 27072
rect 40316 26988 40368 26994
rect 40316 26930 40368 26936
rect 40696 25974 40724 27066
rect 40788 26042 40816 27610
rect 41616 27606 41644 28018
rect 41604 27600 41656 27606
rect 41604 27542 41656 27548
rect 41420 27464 41472 27470
rect 41420 27406 41472 27412
rect 41432 27044 41460 27406
rect 41604 27056 41656 27062
rect 41432 27016 41604 27044
rect 41432 26382 41460 27016
rect 41604 26998 41656 27004
rect 41800 26586 41828 31622
rect 41892 30938 41920 33798
rect 42076 33318 42104 34070
rect 42168 34066 42196 37606
rect 42260 37466 42288 37606
rect 42248 37460 42300 37466
rect 42248 37402 42300 37408
rect 42352 36242 42380 41958
rect 42950 41916 43258 41925
rect 42950 41914 42956 41916
rect 43012 41914 43036 41916
rect 43092 41914 43116 41916
rect 43172 41914 43196 41916
rect 43252 41914 43258 41916
rect 43012 41862 43014 41914
rect 43194 41862 43196 41914
rect 42950 41860 42956 41862
rect 43012 41860 43036 41862
rect 43092 41860 43116 41862
rect 43172 41860 43196 41862
rect 43252 41860 43258 41862
rect 42950 41851 43258 41860
rect 42950 40828 43258 40837
rect 42950 40826 42956 40828
rect 43012 40826 43036 40828
rect 43092 40826 43116 40828
rect 43172 40826 43196 40828
rect 43252 40826 43258 40828
rect 43012 40774 43014 40826
rect 43194 40774 43196 40826
rect 42950 40772 42956 40774
rect 43012 40772 43036 40774
rect 43092 40772 43116 40774
rect 43172 40772 43196 40774
rect 43252 40772 43258 40774
rect 42950 40763 43258 40772
rect 42708 40180 42760 40186
rect 42708 40122 42760 40128
rect 42524 37324 42576 37330
rect 42524 37266 42576 37272
rect 42536 37210 42564 37266
rect 42536 37182 42656 37210
rect 42524 36576 42576 36582
rect 42524 36518 42576 36524
rect 42340 36236 42392 36242
rect 42340 36178 42392 36184
rect 42248 36032 42300 36038
rect 42248 35974 42300 35980
rect 42260 35562 42288 35974
rect 42340 35624 42392 35630
rect 42340 35566 42392 35572
rect 42248 35556 42300 35562
rect 42248 35498 42300 35504
rect 42156 34060 42208 34066
rect 42156 34002 42208 34008
rect 42352 33658 42380 35566
rect 42432 35012 42484 35018
rect 42432 34954 42484 34960
rect 42340 33652 42392 33658
rect 42340 33594 42392 33600
rect 42064 33312 42116 33318
rect 42064 33254 42116 33260
rect 42076 32366 42104 33254
rect 42248 32972 42300 32978
rect 42248 32914 42300 32920
rect 42064 32360 42116 32366
rect 42064 32302 42116 32308
rect 42076 31346 42104 32302
rect 42260 31686 42288 32914
rect 42352 32910 42380 33594
rect 42340 32904 42392 32910
rect 42340 32846 42392 32852
rect 42248 31680 42300 31686
rect 42248 31622 42300 31628
rect 42444 31414 42472 34954
rect 42536 32434 42564 36518
rect 42628 35698 42656 37182
rect 42720 36854 42748 40122
rect 42950 39740 43258 39749
rect 42950 39738 42956 39740
rect 43012 39738 43036 39740
rect 43092 39738 43116 39740
rect 43172 39738 43196 39740
rect 43252 39738 43258 39740
rect 43012 39686 43014 39738
rect 43194 39686 43196 39738
rect 42950 39684 42956 39686
rect 43012 39684 43036 39686
rect 43092 39684 43116 39686
rect 43172 39684 43196 39686
rect 43252 39684 43258 39686
rect 42950 39675 43258 39684
rect 43812 39636 43864 39642
rect 43812 39578 43864 39584
rect 43904 39636 43956 39642
rect 43904 39578 43956 39584
rect 42800 39500 42852 39506
rect 42800 39442 42852 39448
rect 42812 38486 42840 39442
rect 43444 39364 43496 39370
rect 43444 39306 43496 39312
rect 43456 39030 43484 39306
rect 43444 39024 43496 39030
rect 43444 38966 43496 38972
rect 42950 38652 43258 38661
rect 42950 38650 42956 38652
rect 43012 38650 43036 38652
rect 43092 38650 43116 38652
rect 43172 38650 43196 38652
rect 43252 38650 43258 38652
rect 43012 38598 43014 38650
rect 43194 38598 43196 38650
rect 42950 38596 42956 38598
rect 43012 38596 43036 38598
rect 43092 38596 43116 38598
rect 43172 38596 43196 38598
rect 43252 38596 43258 38598
rect 42950 38587 43258 38596
rect 42800 38480 42852 38486
rect 42800 38422 42852 38428
rect 43352 38480 43404 38486
rect 43352 38422 43404 38428
rect 43168 38004 43220 38010
rect 43168 37946 43220 37952
rect 43180 37806 43208 37946
rect 43168 37800 43220 37806
rect 43168 37742 43220 37748
rect 42950 37564 43258 37573
rect 42950 37562 42956 37564
rect 43012 37562 43036 37564
rect 43092 37562 43116 37564
rect 43172 37562 43196 37564
rect 43252 37562 43258 37564
rect 43012 37510 43014 37562
rect 43194 37510 43196 37562
rect 42950 37508 42956 37510
rect 43012 37508 43036 37510
rect 43092 37508 43116 37510
rect 43172 37508 43196 37510
rect 43252 37508 43258 37510
rect 42950 37499 43258 37508
rect 42708 36848 42760 36854
rect 42708 36790 42760 36796
rect 43364 36718 43392 38422
rect 43456 38282 43484 38966
rect 43444 38276 43496 38282
rect 43444 38218 43496 38224
rect 43456 37194 43484 38218
rect 43536 37460 43588 37466
rect 43536 37402 43588 37408
rect 43444 37188 43496 37194
rect 43444 37130 43496 37136
rect 43352 36712 43404 36718
rect 43352 36654 43404 36660
rect 43456 36650 43484 37130
rect 43444 36644 43496 36650
rect 43444 36586 43496 36592
rect 42950 36476 43258 36485
rect 42950 36474 42956 36476
rect 43012 36474 43036 36476
rect 43092 36474 43116 36476
rect 43172 36474 43196 36476
rect 43252 36474 43258 36476
rect 43012 36422 43014 36474
rect 43194 36422 43196 36474
rect 42950 36420 42956 36422
rect 43012 36420 43036 36422
rect 43092 36420 43116 36422
rect 43172 36420 43196 36422
rect 43252 36420 43258 36422
rect 42950 36411 43258 36420
rect 42800 36304 42852 36310
rect 42800 36246 42852 36252
rect 42708 36236 42760 36242
rect 42708 36178 42760 36184
rect 42616 35692 42668 35698
rect 42616 35634 42668 35640
rect 42628 35154 42656 35634
rect 42720 35494 42748 36178
rect 42708 35488 42760 35494
rect 42708 35430 42760 35436
rect 42616 35148 42668 35154
rect 42616 35090 42668 35096
rect 42720 35018 42748 35430
rect 42708 35012 42760 35018
rect 42708 34954 42760 34960
rect 42720 34542 42748 34954
rect 42812 34746 42840 36246
rect 43456 35766 43484 36586
rect 43168 35760 43220 35766
rect 43444 35760 43496 35766
rect 43220 35708 43392 35714
rect 43168 35702 43392 35708
rect 43444 35702 43496 35708
rect 43180 35686 43392 35702
rect 42950 35388 43258 35397
rect 42950 35386 42956 35388
rect 43012 35386 43036 35388
rect 43092 35386 43116 35388
rect 43172 35386 43196 35388
rect 43252 35386 43258 35388
rect 43012 35334 43014 35386
rect 43194 35334 43196 35386
rect 42950 35332 42956 35334
rect 43012 35332 43036 35334
rect 43092 35332 43116 35334
rect 43172 35332 43196 35334
rect 43252 35332 43258 35334
rect 42950 35323 43258 35332
rect 42800 34740 42852 34746
rect 42800 34682 42852 34688
rect 42708 34536 42760 34542
rect 42708 34478 42760 34484
rect 42950 34300 43258 34309
rect 42950 34298 42956 34300
rect 43012 34298 43036 34300
rect 43092 34298 43116 34300
rect 43172 34298 43196 34300
rect 43252 34298 43258 34300
rect 43012 34246 43014 34298
rect 43194 34246 43196 34298
rect 42950 34244 42956 34246
rect 43012 34244 43036 34246
rect 43092 34244 43116 34246
rect 43172 34244 43196 34246
rect 43252 34244 43258 34246
rect 42950 34235 43258 34244
rect 42616 33584 42668 33590
rect 42616 33526 42668 33532
rect 42524 32428 42576 32434
rect 42524 32370 42576 32376
rect 42628 31754 42656 33526
rect 42950 33212 43258 33221
rect 42950 33210 42956 33212
rect 43012 33210 43036 33212
rect 43092 33210 43116 33212
rect 43172 33210 43196 33212
rect 43252 33210 43258 33212
rect 43012 33158 43014 33210
rect 43194 33158 43196 33210
rect 42950 33156 42956 33158
rect 43012 33156 43036 33158
rect 43092 33156 43116 33158
rect 43172 33156 43196 33158
rect 43252 33156 43258 33158
rect 42950 33147 43258 33156
rect 42800 32224 42852 32230
rect 42800 32166 42852 32172
rect 42708 31884 42760 31890
rect 42708 31826 42760 31832
rect 42616 31748 42668 31754
rect 42616 31690 42668 31696
rect 42432 31408 42484 31414
rect 42432 31350 42484 31356
rect 42064 31340 42116 31346
rect 42064 31282 42116 31288
rect 42156 31272 42208 31278
rect 42156 31214 42208 31220
rect 41880 30932 41932 30938
rect 41880 30874 41932 30880
rect 42168 30734 42196 31214
rect 42156 30728 42208 30734
rect 42156 30670 42208 30676
rect 41972 30592 42024 30598
rect 41972 30534 42024 30540
rect 41788 26580 41840 26586
rect 41788 26522 41840 26528
rect 41420 26376 41472 26382
rect 41420 26318 41472 26324
rect 41432 26234 41460 26318
rect 41432 26206 41644 26234
rect 40776 26036 40828 26042
rect 40776 25978 40828 25984
rect 40684 25968 40736 25974
rect 40684 25910 40736 25916
rect 40696 25362 40724 25910
rect 40684 25356 40736 25362
rect 40684 25298 40736 25304
rect 40408 25152 40460 25158
rect 40408 25094 40460 25100
rect 40420 24818 40448 25094
rect 40408 24812 40460 24818
rect 40408 24754 40460 24760
rect 40788 24274 40816 25978
rect 41616 25906 41644 26206
rect 41984 25906 42012 30534
rect 42628 30258 42656 31690
rect 42616 30252 42668 30258
rect 42616 30194 42668 30200
rect 42720 29850 42748 31826
rect 42812 31482 42840 32166
rect 42950 32124 43258 32133
rect 42950 32122 42956 32124
rect 43012 32122 43036 32124
rect 43092 32122 43116 32124
rect 43172 32122 43196 32124
rect 43252 32122 43258 32124
rect 43012 32070 43014 32122
rect 43194 32070 43196 32122
rect 42950 32068 42956 32070
rect 43012 32068 43036 32070
rect 43092 32068 43116 32070
rect 43172 32068 43196 32070
rect 43252 32068 43258 32070
rect 42950 32059 43258 32068
rect 43364 31958 43392 35686
rect 43456 35018 43484 35702
rect 43548 35154 43576 37402
rect 43536 35148 43588 35154
rect 43536 35090 43588 35096
rect 43444 35012 43496 35018
rect 43444 34954 43496 34960
rect 43456 33590 43484 34954
rect 43548 34542 43576 35090
rect 43536 34536 43588 34542
rect 43536 34478 43588 34484
rect 43444 33584 43496 33590
rect 43444 33526 43496 33532
rect 43824 32910 43852 39578
rect 43916 38894 43944 39578
rect 43904 38888 43956 38894
rect 43904 38830 43956 38836
rect 43812 32904 43864 32910
rect 43812 32846 43864 32852
rect 43352 31952 43404 31958
rect 43352 31894 43404 31900
rect 44008 31793 44036 54062
rect 45192 53984 45244 53990
rect 45192 53926 45244 53932
rect 45204 42362 45232 53926
rect 46768 53650 46796 56200
rect 48240 54618 48268 56200
rect 48240 54590 48360 54618
rect 47950 54428 48258 54437
rect 47950 54426 47956 54428
rect 48012 54426 48036 54428
rect 48092 54426 48116 54428
rect 48172 54426 48196 54428
rect 48252 54426 48258 54428
rect 48012 54374 48014 54426
rect 48194 54374 48196 54426
rect 47950 54372 47956 54374
rect 48012 54372 48036 54374
rect 48092 54372 48116 54374
rect 48172 54372 48196 54374
rect 48252 54372 48258 54374
rect 47950 54363 48258 54372
rect 48332 54210 48360 54590
rect 47860 54188 47912 54194
rect 47860 54130 47912 54136
rect 48240 54182 48360 54210
rect 46756 53644 46808 53650
rect 46756 53586 46808 53592
rect 46204 53576 46256 53582
rect 46204 53518 46256 53524
rect 46216 53242 46244 53518
rect 46204 53236 46256 53242
rect 46204 53178 46256 53184
rect 46388 53100 46440 53106
rect 46388 53042 46440 53048
rect 47676 53100 47728 53106
rect 47676 53042 47728 53048
rect 46400 45558 46428 53042
rect 46388 45552 46440 45558
rect 46388 45494 46440 45500
rect 45192 42356 45244 42362
rect 45192 42298 45244 42304
rect 46400 39370 46428 45494
rect 46940 45280 46992 45286
rect 46940 45222 46992 45228
rect 46388 39364 46440 39370
rect 46388 39306 46440 39312
rect 46952 37738 46980 45222
rect 46940 37732 46992 37738
rect 46940 37674 46992 37680
rect 44364 37664 44416 37670
rect 44364 37606 44416 37612
rect 44272 34536 44324 34542
rect 44272 34478 44324 34484
rect 43994 31784 44050 31793
rect 43994 31719 44050 31728
rect 42800 31476 42852 31482
rect 42800 31418 42852 31424
rect 44284 31346 44312 34478
rect 44272 31340 44324 31346
rect 44272 31282 44324 31288
rect 44376 31278 44404 37606
rect 46940 36576 46992 36582
rect 46940 36518 46992 36524
rect 46952 34950 46980 36518
rect 44548 34944 44600 34950
rect 44548 34886 44600 34892
rect 46940 34944 46992 34950
rect 46940 34886 46992 34892
rect 44560 34610 44588 34886
rect 44548 34604 44600 34610
rect 44548 34546 44600 34552
rect 47216 32768 47268 32774
rect 47216 32710 47268 32716
rect 45284 32292 45336 32298
rect 45284 32234 45336 32240
rect 44824 32224 44876 32230
rect 44824 32166 44876 32172
rect 44364 31272 44416 31278
rect 44364 31214 44416 31220
rect 42950 31036 43258 31045
rect 42950 31034 42956 31036
rect 43012 31034 43036 31036
rect 43092 31034 43116 31036
rect 43172 31034 43196 31036
rect 43252 31034 43258 31036
rect 43012 30982 43014 31034
rect 43194 30982 43196 31034
rect 42950 30980 42956 30982
rect 43012 30980 43036 30982
rect 43092 30980 43116 30982
rect 43172 30980 43196 30982
rect 43252 30980 43258 30982
rect 42950 30971 43258 30980
rect 42950 29948 43258 29957
rect 42950 29946 42956 29948
rect 43012 29946 43036 29948
rect 43092 29946 43116 29948
rect 43172 29946 43196 29948
rect 43252 29946 43258 29948
rect 43012 29894 43014 29946
rect 43194 29894 43196 29946
rect 42950 29892 42956 29894
rect 43012 29892 43036 29894
rect 43092 29892 43116 29894
rect 43172 29892 43196 29894
rect 43252 29892 43258 29894
rect 42950 29883 43258 29892
rect 42708 29844 42760 29850
rect 42708 29786 42760 29792
rect 42720 29102 42748 29786
rect 42708 29096 42760 29102
rect 42708 29038 42760 29044
rect 44180 29028 44232 29034
rect 44180 28970 44232 28976
rect 42950 28860 43258 28869
rect 42950 28858 42956 28860
rect 43012 28858 43036 28860
rect 43092 28858 43116 28860
rect 43172 28858 43196 28860
rect 43252 28858 43258 28860
rect 43012 28806 43014 28858
rect 43194 28806 43196 28858
rect 42950 28804 42956 28806
rect 43012 28804 43036 28806
rect 43092 28804 43116 28806
rect 43172 28804 43196 28806
rect 43252 28804 43258 28806
rect 42950 28795 43258 28804
rect 42950 27772 43258 27781
rect 42950 27770 42956 27772
rect 43012 27770 43036 27772
rect 43092 27770 43116 27772
rect 43172 27770 43196 27772
rect 43252 27770 43258 27772
rect 43012 27718 43014 27770
rect 43194 27718 43196 27770
rect 42950 27716 42956 27718
rect 43012 27716 43036 27718
rect 43092 27716 43116 27718
rect 43172 27716 43196 27718
rect 43252 27716 43258 27718
rect 42950 27707 43258 27716
rect 44192 27470 44220 28970
rect 44180 27464 44232 27470
rect 44180 27406 44232 27412
rect 43996 27328 44048 27334
rect 43996 27270 44048 27276
rect 42154 27160 42210 27169
rect 42154 27095 42156 27104
rect 42208 27095 42210 27104
rect 42156 27066 42208 27072
rect 42950 26684 43258 26693
rect 42950 26682 42956 26684
rect 43012 26682 43036 26684
rect 43092 26682 43116 26684
rect 43172 26682 43196 26684
rect 43252 26682 43258 26684
rect 43012 26630 43014 26682
rect 43194 26630 43196 26682
rect 42950 26628 42956 26630
rect 43012 26628 43036 26630
rect 43092 26628 43116 26630
rect 43172 26628 43196 26630
rect 43252 26628 43258 26630
rect 42950 26619 43258 26628
rect 44008 26382 44036 27270
rect 44836 27062 44864 32166
rect 44824 27056 44876 27062
rect 44824 26998 44876 27004
rect 42800 26376 42852 26382
rect 42800 26318 42852 26324
rect 43996 26376 44048 26382
rect 43996 26318 44048 26324
rect 41604 25900 41656 25906
rect 41604 25842 41656 25848
rect 41972 25900 42024 25906
rect 41972 25842 42024 25848
rect 40224 24268 40276 24274
rect 40224 24210 40276 24216
rect 40776 24268 40828 24274
rect 40776 24210 40828 24216
rect 40040 24200 40092 24206
rect 40040 24142 40092 24148
rect 40040 24064 40092 24070
rect 40040 24006 40092 24012
rect 39580 23792 39632 23798
rect 39580 23734 39632 23740
rect 39592 22710 39620 23734
rect 39580 22704 39632 22710
rect 39580 22646 39632 22652
rect 39488 22568 39540 22574
rect 39488 22510 39540 22516
rect 39212 18624 39264 18630
rect 39212 18566 39264 18572
rect 38672 18278 38792 18306
rect 38016 18216 38068 18222
rect 38016 18158 38068 18164
rect 38568 18216 38620 18222
rect 38568 18158 38620 18164
rect 38028 17746 38056 18158
rect 38200 17876 38252 17882
rect 38200 17818 38252 17824
rect 38212 17762 38240 17818
rect 38016 17740 38068 17746
rect 38212 17734 38332 17762
rect 38016 17682 38068 17688
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 38108 16992 38160 16998
rect 38108 16934 38160 16940
rect 38120 16590 38148 16934
rect 38108 16584 38160 16590
rect 38108 16526 38160 16532
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 37832 13932 37884 13938
rect 37832 13874 37884 13880
rect 37740 13388 37792 13394
rect 37740 13330 37792 13336
rect 37188 13320 37240 13326
rect 37188 13262 37240 13268
rect 37372 13320 37424 13326
rect 37372 13262 37424 13268
rect 37280 13184 37332 13190
rect 37280 13126 37332 13132
rect 36728 3528 36780 3534
rect 36728 3470 36780 3476
rect 37292 3126 37320 13126
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 38304 12238 38332 17734
rect 38672 17610 38700 18278
rect 39764 18080 39816 18086
rect 39764 18022 39816 18028
rect 38660 17604 38712 17610
rect 38660 17546 38712 17552
rect 38672 17338 38700 17546
rect 38660 17332 38712 17338
rect 38660 17274 38712 17280
rect 39488 16448 39540 16454
rect 39488 16390 39540 16396
rect 38476 15904 38528 15910
rect 38476 15846 38528 15852
rect 38384 13864 38436 13870
rect 38384 13806 38436 13812
rect 38292 12232 38344 12238
rect 38292 12174 38344 12180
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37372 9444 37424 9450
rect 37372 9386 37424 9392
rect 37384 3534 37412 9386
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 37648 8356 37700 8362
rect 37648 8298 37700 8304
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 37280 3120 37332 3126
rect 37280 3062 37332 3068
rect 37660 3058 37688 8298
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 38396 4146 38424 13806
rect 38488 8566 38516 15846
rect 39120 15700 39172 15706
rect 39120 15642 39172 15648
rect 38568 14068 38620 14074
rect 38568 14010 38620 14016
rect 38580 12918 38608 14010
rect 39132 13938 39160 15642
rect 39500 13938 39528 16390
rect 39776 15026 39804 18022
rect 39948 17060 40000 17066
rect 39948 17002 40000 17008
rect 39764 15020 39816 15026
rect 39764 14962 39816 14968
rect 39764 14544 39816 14550
rect 39764 14486 39816 14492
rect 39120 13932 39172 13938
rect 39120 13874 39172 13880
rect 39488 13932 39540 13938
rect 39488 13874 39540 13880
rect 38568 12912 38620 12918
rect 38568 12854 38620 12860
rect 39776 11762 39804 14486
rect 39960 14414 39988 17002
rect 40052 16114 40080 24006
rect 42812 22710 42840 26318
rect 42950 25596 43258 25605
rect 42950 25594 42956 25596
rect 43012 25594 43036 25596
rect 43092 25594 43116 25596
rect 43172 25594 43196 25596
rect 43252 25594 43258 25596
rect 43012 25542 43014 25594
rect 43194 25542 43196 25594
rect 42950 25540 42956 25542
rect 43012 25540 43036 25542
rect 43092 25540 43116 25542
rect 43172 25540 43196 25542
rect 43252 25540 43258 25542
rect 42950 25531 43258 25540
rect 45296 25294 45324 32234
rect 45744 31408 45796 31414
rect 45744 31350 45796 31356
rect 45756 30054 45784 31350
rect 46020 31204 46072 31210
rect 46020 31146 46072 31152
rect 45744 30048 45796 30054
rect 45744 29990 45796 29996
rect 46032 25294 46060 31146
rect 46940 31136 46992 31142
rect 46940 31078 46992 31084
rect 46112 30660 46164 30666
rect 46112 30602 46164 30608
rect 46124 25974 46152 30602
rect 46952 28150 46980 31078
rect 47032 30592 47084 30598
rect 47032 30534 47084 30540
rect 46940 28144 46992 28150
rect 46940 28086 46992 28092
rect 47044 26994 47072 30534
rect 47124 27532 47176 27538
rect 47124 27474 47176 27480
rect 47136 26994 47164 27474
rect 47228 27470 47256 32710
rect 47400 31340 47452 31346
rect 47400 31282 47452 31288
rect 47216 27464 47268 27470
rect 47216 27406 47268 27412
rect 47032 26988 47084 26994
rect 47032 26930 47084 26936
rect 47124 26988 47176 26994
rect 47124 26930 47176 26936
rect 46756 26784 46808 26790
rect 46756 26726 46808 26732
rect 46112 25968 46164 25974
rect 46112 25910 46164 25916
rect 46296 25764 46348 25770
rect 46296 25706 46348 25712
rect 45284 25288 45336 25294
rect 45284 25230 45336 25236
rect 46020 25288 46072 25294
rect 46020 25230 46072 25236
rect 44640 25220 44692 25226
rect 44640 25162 44692 25168
rect 45468 25220 45520 25226
rect 45468 25162 45520 25168
rect 43812 24608 43864 24614
rect 43812 24550 43864 24556
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 42800 22704 42852 22710
rect 42800 22646 42852 22652
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 43352 21344 43404 21350
rect 43352 21286 43404 21292
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42800 21140 42852 21146
rect 42800 21082 42852 21088
rect 42812 17678 42840 21082
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 43364 17678 43392 21286
rect 43720 21072 43772 21078
rect 43720 21014 43772 21020
rect 42800 17672 42852 17678
rect 42800 17614 42852 17620
rect 43352 17672 43404 17678
rect 43352 17614 43404 17620
rect 43732 17270 43760 21014
rect 43824 20942 43852 24550
rect 44088 23248 44140 23254
rect 44088 23190 44140 23196
rect 43812 20936 43864 20942
rect 43812 20878 43864 20884
rect 44100 19854 44128 23190
rect 44180 21888 44232 21894
rect 44180 21830 44232 21836
rect 44088 19848 44140 19854
rect 44088 19790 44140 19796
rect 44192 18766 44220 21830
rect 44456 20256 44508 20262
rect 44456 20198 44508 20204
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 44468 17610 44496 20198
rect 44652 18766 44680 25162
rect 45192 20868 45244 20874
rect 45192 20810 45244 20816
rect 44916 19984 44968 19990
rect 44916 19926 44968 19932
rect 44640 18760 44692 18766
rect 44640 18702 44692 18708
rect 44456 17604 44508 17610
rect 44456 17546 44508 17552
rect 44548 17536 44600 17542
rect 44548 17478 44600 17484
rect 43720 17264 43772 17270
rect 43720 17206 43772 17212
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 40040 16108 40092 16114
rect 40040 16050 40092 16056
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 41328 14816 41380 14822
rect 41328 14758 41380 14764
rect 44180 14816 44232 14822
rect 44180 14758 44232 14764
rect 39948 14408 40000 14414
rect 39948 14350 40000 14356
rect 40040 14000 40092 14006
rect 40040 13942 40092 13948
rect 39856 13184 39908 13190
rect 39856 13126 39908 13132
rect 39868 12306 39896 13126
rect 39948 12640 40000 12646
rect 39948 12582 40000 12588
rect 39856 12300 39908 12306
rect 39856 12242 39908 12248
rect 39764 11756 39816 11762
rect 39764 11698 39816 11704
rect 39960 10674 39988 12582
rect 39948 10668 40000 10674
rect 39948 10610 40000 10616
rect 38476 8560 38528 8566
rect 38476 8502 38528 8508
rect 38384 4140 38436 4146
rect 38384 4082 38436 4088
rect 39028 4072 39080 4078
rect 39028 4014 39080 4020
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 37648 3052 37700 3058
rect 37648 2994 37700 3000
rect 36820 2984 36872 2990
rect 36820 2926 36872 2932
rect 36832 800 36860 2926
rect 37556 2916 37608 2922
rect 37556 2858 37608 2864
rect 37568 800 37596 2858
rect 38292 2508 38344 2514
rect 38292 2450 38344 2456
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38304 800 38332 2450
rect 39040 800 39068 4014
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39776 800 39804 3538
rect 40052 2446 40080 13942
rect 40684 13864 40736 13870
rect 40684 13806 40736 13812
rect 40696 13326 40724 13806
rect 40684 13320 40736 13326
rect 40684 13262 40736 13268
rect 41340 12238 41368 14758
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 44088 14272 44140 14278
rect 44088 14214 44140 14220
rect 42708 14068 42760 14074
rect 42708 14010 42760 14016
rect 41328 12232 41380 12238
rect 41328 12174 41380 12180
rect 41880 12164 41932 12170
rect 41880 12106 41932 12112
rect 41420 7200 41472 7206
rect 41420 7142 41472 7148
rect 40132 6792 40184 6798
rect 40132 6734 40184 6740
rect 40144 4146 40172 6734
rect 40132 4140 40184 4146
rect 40132 4082 40184 4088
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 40592 2508 40644 2514
rect 40512 2468 40592 2496
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 40512 800 40540 2468
rect 40592 2450 40644 2456
rect 41248 800 41276 3538
rect 41432 2446 41460 7142
rect 41892 3534 41920 12106
rect 42720 11762 42748 14010
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 43352 12096 43404 12102
rect 43352 12038 43404 12044
rect 42708 11756 42760 11762
rect 42708 11698 42760 11704
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 42708 10464 42760 10470
rect 42708 10406 42760 10412
rect 42720 8566 42748 10406
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 43364 8974 43392 12038
rect 44100 11694 44128 14214
rect 44192 11830 44220 14758
rect 44364 13864 44416 13870
rect 44364 13806 44416 13812
rect 44272 12096 44324 12102
rect 44272 12038 44324 12044
rect 44180 11824 44232 11830
rect 44180 11766 44232 11772
rect 44088 11688 44140 11694
rect 44088 11630 44140 11636
rect 44180 11552 44232 11558
rect 44180 11494 44232 11500
rect 44192 9586 44220 11494
rect 44284 11150 44312 12038
rect 44272 11144 44324 11150
rect 44272 11086 44324 11092
rect 44376 11082 44404 13806
rect 44560 13326 44588 17478
rect 44548 13320 44600 13326
rect 44548 13262 44600 13268
rect 44732 12708 44784 12714
rect 44732 12650 44784 12656
rect 44744 12238 44772 12650
rect 44732 12232 44784 12238
rect 44732 12174 44784 12180
rect 44364 11076 44416 11082
rect 44364 11018 44416 11024
rect 44180 9580 44232 9586
rect 44180 9522 44232 9528
rect 43352 8968 43404 8974
rect 43352 8910 43404 8916
rect 42708 8560 42760 8566
rect 42708 8502 42760 8508
rect 42616 8424 42668 8430
rect 42616 8366 42668 8372
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42628 3058 42656 8366
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 44456 6724 44508 6730
rect 44456 6666 44508 6672
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 43444 4072 43496 4078
rect 43444 4014 43496 4020
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 41972 2984 42024 2990
rect 41972 2926 42024 2932
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 41984 800 42012 2926
rect 42708 2916 42760 2922
rect 42708 2858 42760 2864
rect 42720 800 42748 2858
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 43456 800 43484 4014
rect 44180 3596 44232 3602
rect 44180 3538 44232 3544
rect 44192 800 44220 3538
rect 44468 3058 44496 6666
rect 44456 3052 44508 3058
rect 44456 2994 44508 3000
rect 44928 800 44956 19926
rect 45204 17678 45232 20810
rect 45480 19378 45508 25162
rect 46308 21554 46336 25706
rect 46768 23730 46796 26726
rect 47216 26240 47268 26246
rect 47216 26182 47268 26188
rect 47032 25764 47084 25770
rect 47032 25706 47084 25712
rect 46756 23724 46808 23730
rect 46756 23666 46808 23672
rect 46756 22500 46808 22506
rect 46756 22442 46808 22448
rect 46296 21548 46348 21554
rect 46296 21490 46348 21496
rect 46204 19780 46256 19786
rect 46204 19722 46256 19728
rect 45468 19372 45520 19378
rect 45468 19314 45520 19320
rect 45192 17672 45244 17678
rect 45192 17614 45244 17620
rect 46216 16590 46244 19722
rect 46768 18290 46796 22442
rect 47044 20942 47072 25706
rect 47228 24818 47256 26182
rect 47216 24812 47268 24818
rect 47216 24754 47268 24760
rect 47032 20936 47084 20942
rect 47032 20878 47084 20884
rect 46756 18284 46808 18290
rect 46756 18226 46808 18232
rect 46848 17604 46900 17610
rect 46848 17546 46900 17552
rect 46664 17536 46716 17542
rect 46664 17478 46716 17484
rect 46204 16584 46256 16590
rect 46204 16526 46256 16532
rect 46676 13938 46704 17478
rect 46756 17060 46808 17066
rect 46756 17002 46808 17008
rect 46768 15026 46796 17002
rect 46860 15502 46888 17546
rect 46848 15496 46900 15502
rect 46848 15438 46900 15444
rect 46756 15020 46808 15026
rect 46756 14962 46808 14968
rect 46664 13932 46716 13938
rect 46664 13874 46716 13880
rect 46756 13184 46808 13190
rect 46756 13126 46808 13132
rect 46020 12980 46072 12986
rect 46020 12922 46072 12928
rect 45928 8356 45980 8362
rect 45928 8298 45980 8304
rect 45192 7268 45244 7274
rect 45192 7210 45244 7216
rect 45204 3534 45232 7210
rect 45940 6866 45968 8298
rect 45928 6860 45980 6866
rect 45928 6802 45980 6808
rect 46032 4146 46060 12922
rect 46768 12850 46796 13126
rect 46756 12844 46808 12850
rect 46756 12786 46808 12792
rect 46756 11688 46808 11694
rect 46756 11630 46808 11636
rect 46664 11620 46716 11626
rect 46664 11562 46716 11568
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46204 8900 46256 8906
rect 46204 8842 46256 8848
rect 46216 5710 46244 8842
rect 46308 7886 46336 11494
rect 46480 11076 46532 11082
rect 46480 11018 46532 11024
rect 46492 8498 46520 11018
rect 46676 9586 46704 11562
rect 46768 10062 46796 11630
rect 46756 10056 46808 10062
rect 46756 9998 46808 10004
rect 46664 9580 46716 9586
rect 46664 9522 46716 9528
rect 46480 8492 46532 8498
rect 46480 8434 46532 8440
rect 46296 7880 46348 7886
rect 46296 7822 46348 7828
rect 47412 6798 47440 31282
rect 47688 30938 47716 53042
rect 47872 31482 47900 54130
rect 48240 54126 48268 54182
rect 48228 54120 48280 54126
rect 48228 54062 48280 54068
rect 47950 53340 48258 53349
rect 47950 53338 47956 53340
rect 48012 53338 48036 53340
rect 48092 53338 48116 53340
rect 48172 53338 48196 53340
rect 48252 53338 48258 53340
rect 48012 53286 48014 53338
rect 48194 53286 48196 53338
rect 47950 53284 47956 53286
rect 48012 53284 48036 53286
rect 48092 53284 48116 53286
rect 48172 53284 48196 53286
rect 48252 53284 48258 53286
rect 47950 53275 48258 53284
rect 49712 53174 49740 56200
rect 49700 53168 49752 53174
rect 49700 53110 49752 53116
rect 47950 52252 48258 52261
rect 47950 52250 47956 52252
rect 48012 52250 48036 52252
rect 48092 52250 48116 52252
rect 48172 52250 48196 52252
rect 48252 52250 48258 52252
rect 48012 52198 48014 52250
rect 48194 52198 48196 52250
rect 47950 52196 47956 52198
rect 48012 52196 48036 52198
rect 48092 52196 48116 52198
rect 48172 52196 48196 52198
rect 48252 52196 48258 52198
rect 47950 52187 48258 52196
rect 49056 52012 49108 52018
rect 49056 51954 49108 51960
rect 49068 51921 49096 51954
rect 49054 51912 49110 51921
rect 49054 51847 49110 51856
rect 49240 51808 49292 51814
rect 49240 51750 49292 51756
rect 49056 51400 49108 51406
rect 49056 51342 49108 51348
rect 49068 51241 49096 51342
rect 49148 51264 49200 51270
rect 49054 51232 49110 51241
rect 49148 51206 49200 51212
rect 47950 51164 48258 51173
rect 49054 51167 49110 51176
rect 47950 51162 47956 51164
rect 48012 51162 48036 51164
rect 48092 51162 48116 51164
rect 48172 51162 48196 51164
rect 48252 51162 48258 51164
rect 48012 51110 48014 51162
rect 48194 51110 48196 51162
rect 47950 51108 47956 51110
rect 48012 51108 48036 51110
rect 48092 51108 48116 51110
rect 48172 51108 48196 51110
rect 48252 51108 48258 51110
rect 47950 51099 48258 51108
rect 48964 50924 49016 50930
rect 48964 50866 49016 50872
rect 48976 50561 49004 50866
rect 48962 50552 49018 50561
rect 48962 50487 49018 50496
rect 49056 50312 49108 50318
rect 49056 50254 49108 50260
rect 48412 50176 48464 50182
rect 48412 50118 48464 50124
rect 47950 50076 48258 50085
rect 47950 50074 47956 50076
rect 48012 50074 48036 50076
rect 48092 50074 48116 50076
rect 48172 50074 48196 50076
rect 48252 50074 48258 50076
rect 48012 50022 48014 50074
rect 48194 50022 48196 50074
rect 47950 50020 47956 50022
rect 48012 50020 48036 50022
rect 48092 50020 48116 50022
rect 48172 50020 48196 50022
rect 48252 50020 48258 50022
rect 47950 50011 48258 50020
rect 47950 48988 48258 48997
rect 47950 48986 47956 48988
rect 48012 48986 48036 48988
rect 48092 48986 48116 48988
rect 48172 48986 48196 48988
rect 48252 48986 48258 48988
rect 48012 48934 48014 48986
rect 48194 48934 48196 48986
rect 47950 48932 47956 48934
rect 48012 48932 48036 48934
rect 48092 48932 48116 48934
rect 48172 48932 48196 48934
rect 48252 48932 48258 48934
rect 47950 48923 48258 48932
rect 47950 47900 48258 47909
rect 47950 47898 47956 47900
rect 48012 47898 48036 47900
rect 48092 47898 48116 47900
rect 48172 47898 48196 47900
rect 48252 47898 48258 47900
rect 48012 47846 48014 47898
rect 48194 47846 48196 47898
rect 47950 47844 47956 47846
rect 48012 47844 48036 47846
rect 48092 47844 48116 47846
rect 48172 47844 48196 47846
rect 48252 47844 48258 47846
rect 47950 47835 48258 47844
rect 47950 46812 48258 46821
rect 47950 46810 47956 46812
rect 48012 46810 48036 46812
rect 48092 46810 48116 46812
rect 48172 46810 48196 46812
rect 48252 46810 48258 46812
rect 48012 46758 48014 46810
rect 48194 46758 48196 46810
rect 47950 46756 47956 46758
rect 48012 46756 48036 46758
rect 48092 46756 48116 46758
rect 48172 46756 48196 46758
rect 48252 46756 48258 46758
rect 47950 46747 48258 46756
rect 47950 45724 48258 45733
rect 47950 45722 47956 45724
rect 48012 45722 48036 45724
rect 48092 45722 48116 45724
rect 48172 45722 48196 45724
rect 48252 45722 48258 45724
rect 48012 45670 48014 45722
rect 48194 45670 48196 45722
rect 47950 45668 47956 45670
rect 48012 45668 48036 45670
rect 48092 45668 48116 45670
rect 48172 45668 48196 45670
rect 48252 45668 48258 45670
rect 47950 45659 48258 45668
rect 48320 45484 48372 45490
rect 48320 45426 48372 45432
rect 48332 45121 48360 45426
rect 48318 45112 48374 45121
rect 48318 45047 48374 45056
rect 47950 44636 48258 44645
rect 47950 44634 47956 44636
rect 48012 44634 48036 44636
rect 48092 44634 48116 44636
rect 48172 44634 48196 44636
rect 48252 44634 48258 44636
rect 48012 44582 48014 44634
rect 48194 44582 48196 44634
rect 47950 44580 47956 44582
rect 48012 44580 48036 44582
rect 48092 44580 48116 44582
rect 48172 44580 48196 44582
rect 48252 44580 48258 44582
rect 47950 44571 48258 44580
rect 47950 43548 48258 43557
rect 47950 43546 47956 43548
rect 48012 43546 48036 43548
rect 48092 43546 48116 43548
rect 48172 43546 48196 43548
rect 48252 43546 48258 43548
rect 48012 43494 48014 43546
rect 48194 43494 48196 43546
rect 47950 43492 47956 43494
rect 48012 43492 48036 43494
rect 48092 43492 48116 43494
rect 48172 43492 48196 43494
rect 48252 43492 48258 43494
rect 47950 43483 48258 43492
rect 47950 42460 48258 42469
rect 47950 42458 47956 42460
rect 48012 42458 48036 42460
rect 48092 42458 48116 42460
rect 48172 42458 48196 42460
rect 48252 42458 48258 42460
rect 48012 42406 48014 42458
rect 48194 42406 48196 42458
rect 47950 42404 47956 42406
rect 48012 42404 48036 42406
rect 48092 42404 48116 42406
rect 48172 42404 48196 42406
rect 48252 42404 48258 42406
rect 47950 42395 48258 42404
rect 47950 41372 48258 41381
rect 47950 41370 47956 41372
rect 48012 41370 48036 41372
rect 48092 41370 48116 41372
rect 48172 41370 48196 41372
rect 48252 41370 48258 41372
rect 48012 41318 48014 41370
rect 48194 41318 48196 41370
rect 47950 41316 47956 41318
rect 48012 41316 48036 41318
rect 48092 41316 48116 41318
rect 48172 41316 48196 41318
rect 48252 41316 48258 41318
rect 47950 41307 48258 41316
rect 48424 40746 48452 50118
rect 49068 49881 49096 50254
rect 49054 49872 49110 49881
rect 49054 49807 49110 49816
rect 49056 49224 49108 49230
rect 49054 49192 49056 49201
rect 49108 49192 49110 49201
rect 49054 49127 49110 49136
rect 48872 49088 48924 49094
rect 48872 49030 48924 49036
rect 48688 47456 48740 47462
rect 48688 47398 48740 47404
rect 48596 45960 48648 45966
rect 48596 45902 48648 45908
rect 48608 45626 48636 45902
rect 48596 45620 48648 45626
rect 48596 45562 48648 45568
rect 48504 44872 48556 44878
rect 48504 44814 48556 44820
rect 48516 44441 48544 44814
rect 48502 44432 48558 44441
rect 48502 44367 48558 44376
rect 48504 43784 48556 43790
rect 48502 43752 48504 43761
rect 48556 43752 48558 43761
rect 48502 43687 48558 43696
rect 48504 43240 48556 43246
rect 48504 43182 48556 43188
rect 48516 43081 48544 43182
rect 48502 43072 48558 43081
rect 48502 43007 48558 43016
rect 48504 42696 48556 42702
rect 48504 42638 48556 42644
rect 48516 42401 48544 42638
rect 48502 42392 48558 42401
rect 48502 42327 48558 42336
rect 48504 42152 48556 42158
rect 48504 42094 48556 42100
rect 48516 41721 48544 42094
rect 48502 41712 48558 41721
rect 48502 41647 48558 41656
rect 48504 41064 48556 41070
rect 48502 41032 48504 41041
rect 48596 41064 48648 41070
rect 48556 41032 48558 41041
rect 48596 41006 48648 41012
rect 48502 40967 48558 40976
rect 48332 40718 48452 40746
rect 47950 40284 48258 40293
rect 47950 40282 47956 40284
rect 48012 40282 48036 40284
rect 48092 40282 48116 40284
rect 48172 40282 48196 40284
rect 48252 40282 48258 40284
rect 48012 40230 48014 40282
rect 48194 40230 48196 40282
rect 47950 40228 47956 40230
rect 48012 40228 48036 40230
rect 48092 40228 48116 40230
rect 48172 40228 48196 40230
rect 48252 40228 48258 40230
rect 47950 40219 48258 40228
rect 48332 39642 48360 40718
rect 48412 40588 48464 40594
rect 48412 40530 48464 40536
rect 48320 39636 48372 39642
rect 48320 39578 48372 39584
rect 47950 39196 48258 39205
rect 47950 39194 47956 39196
rect 48012 39194 48036 39196
rect 48092 39194 48116 39196
rect 48172 39194 48196 39196
rect 48252 39194 48258 39196
rect 48012 39142 48014 39194
rect 48194 39142 48196 39194
rect 47950 39140 47956 39142
rect 48012 39140 48036 39142
rect 48092 39140 48116 39142
rect 48172 39140 48196 39142
rect 48252 39140 48258 39142
rect 47950 39131 48258 39140
rect 47950 38108 48258 38117
rect 47950 38106 47956 38108
rect 48012 38106 48036 38108
rect 48092 38106 48116 38108
rect 48172 38106 48196 38108
rect 48252 38106 48258 38108
rect 48012 38054 48014 38106
rect 48194 38054 48196 38106
rect 47950 38052 47956 38054
rect 48012 38052 48036 38054
rect 48092 38052 48116 38054
rect 48172 38052 48196 38054
rect 48252 38052 48258 38054
rect 47950 38043 48258 38052
rect 47950 37020 48258 37029
rect 47950 37018 47956 37020
rect 48012 37018 48036 37020
rect 48092 37018 48116 37020
rect 48172 37018 48196 37020
rect 48252 37018 48258 37020
rect 48012 36966 48014 37018
rect 48194 36966 48196 37018
rect 47950 36964 47956 36966
rect 48012 36964 48036 36966
rect 48092 36964 48116 36966
rect 48172 36964 48196 36966
rect 48252 36964 48258 36966
rect 47950 36955 48258 36964
rect 47950 35932 48258 35941
rect 47950 35930 47956 35932
rect 48012 35930 48036 35932
rect 48092 35930 48116 35932
rect 48172 35930 48196 35932
rect 48252 35930 48258 35932
rect 48012 35878 48014 35930
rect 48194 35878 48196 35930
rect 47950 35876 47956 35878
rect 48012 35876 48036 35878
rect 48092 35876 48116 35878
rect 48172 35876 48196 35878
rect 48252 35876 48258 35878
rect 47950 35867 48258 35876
rect 48424 35086 48452 40530
rect 48504 40520 48556 40526
rect 48504 40462 48556 40468
rect 48516 40361 48544 40462
rect 48502 40352 48558 40361
rect 48502 40287 48558 40296
rect 48504 39976 48556 39982
rect 48504 39918 48556 39924
rect 48516 39681 48544 39918
rect 48502 39672 48558 39681
rect 48502 39607 48558 39616
rect 48504 39432 48556 39438
rect 48504 39374 48556 39380
rect 48516 39001 48544 39374
rect 48502 38992 48558 39001
rect 48502 38927 48558 38936
rect 48504 37324 48556 37330
rect 48504 37266 48556 37272
rect 48516 36961 48544 37266
rect 48502 36952 48558 36961
rect 48502 36887 48558 36896
rect 48608 35601 48636 41006
rect 48700 38418 48728 47398
rect 48778 39536 48834 39545
rect 48778 39471 48780 39480
rect 48832 39471 48834 39480
rect 48780 39442 48832 39448
rect 48688 38412 48740 38418
rect 48688 38354 48740 38360
rect 48884 38214 48912 49030
rect 49056 48748 49108 48754
rect 49056 48690 49108 48696
rect 48964 48544 49016 48550
rect 49068 48521 49096 48690
rect 48964 48486 49016 48492
rect 49054 48512 49110 48521
rect 48872 38208 48924 38214
rect 48872 38150 48924 38156
rect 48780 37256 48832 37262
rect 48780 37198 48832 37204
rect 48792 36378 48820 37198
rect 48976 36922 49004 48486
rect 49054 48447 49110 48456
rect 49056 48136 49108 48142
rect 49056 48078 49108 48084
rect 49068 47841 49096 48078
rect 49054 47832 49110 47841
rect 49054 47767 49110 47776
rect 49056 47660 49108 47666
rect 49056 47602 49108 47608
rect 49068 47161 49096 47602
rect 49054 47152 49110 47161
rect 49054 47087 49110 47096
rect 49160 46050 49188 51206
rect 49068 46022 49188 46050
rect 49068 45554 49096 46022
rect 49148 45892 49200 45898
rect 49148 45834 49200 45840
rect 49160 45801 49188 45834
rect 49146 45792 49202 45801
rect 49146 45727 49202 45736
rect 49068 45526 49188 45554
rect 48964 36916 49016 36922
rect 48964 36858 49016 36864
rect 48780 36372 48832 36378
rect 48780 36314 48832 36320
rect 49160 35894 49188 45526
rect 48976 35866 49188 35894
rect 48594 35592 48650 35601
rect 48594 35527 48650 35536
rect 48412 35080 48464 35086
rect 48412 35022 48464 35028
rect 47950 34844 48258 34853
rect 47950 34842 47956 34844
rect 48012 34842 48036 34844
rect 48092 34842 48116 34844
rect 48172 34842 48196 34844
rect 48252 34842 48258 34844
rect 48012 34790 48014 34842
rect 48194 34790 48196 34842
rect 47950 34788 47956 34790
rect 48012 34788 48036 34790
rect 48092 34788 48116 34790
rect 48172 34788 48196 34790
rect 48252 34788 48258 34790
rect 47950 34779 48258 34788
rect 48976 34202 49004 35866
rect 49056 35828 49108 35834
rect 49056 35770 49108 35776
rect 49068 34950 49096 35770
rect 49148 35284 49200 35290
rect 49148 35226 49200 35232
rect 49056 34944 49108 34950
rect 49056 34886 49108 34892
rect 49160 34746 49188 35226
rect 49148 34740 49200 34746
rect 49148 34682 49200 34688
rect 48964 34196 49016 34202
rect 48964 34138 49016 34144
rect 49252 33930 49280 51750
rect 49424 50720 49476 50726
rect 49424 50662 49476 50668
rect 49332 38344 49384 38350
rect 49330 38312 49332 38321
rect 49384 38312 49386 38321
rect 49330 38247 49386 38256
rect 49332 37868 49384 37874
rect 49332 37810 49384 37816
rect 49344 37641 49372 37810
rect 49330 37632 49386 37641
rect 49330 37567 49386 37576
rect 49436 37233 49464 50662
rect 49422 37224 49478 37233
rect 49422 37159 49478 37168
rect 49332 36780 49384 36786
rect 49332 36722 49384 36728
rect 49344 36281 49372 36722
rect 49330 36272 49386 36281
rect 49330 36207 49386 36216
rect 49332 35692 49384 35698
rect 49332 35634 49384 35640
rect 49344 35601 49372 35634
rect 49330 35592 49386 35601
rect 49330 35527 49386 35536
rect 49332 35080 49384 35086
rect 49332 35022 49384 35028
rect 49344 34921 49372 35022
rect 49330 34912 49386 34921
rect 49330 34847 49386 34856
rect 49332 34604 49384 34610
rect 49332 34546 49384 34552
rect 49344 34241 49372 34546
rect 49330 34232 49386 34241
rect 49330 34167 49386 34176
rect 49332 33992 49384 33998
rect 49332 33934 49384 33940
rect 49240 33924 49292 33930
rect 49240 33866 49292 33872
rect 47950 33756 48258 33765
rect 47950 33754 47956 33756
rect 48012 33754 48036 33756
rect 48092 33754 48116 33756
rect 48172 33754 48196 33756
rect 48252 33754 48258 33756
rect 48012 33702 48014 33754
rect 48194 33702 48196 33754
rect 47950 33700 47956 33702
rect 48012 33700 48036 33702
rect 48092 33700 48116 33702
rect 48172 33700 48196 33702
rect 48252 33700 48258 33702
rect 47950 33691 48258 33700
rect 49344 33561 49372 33934
rect 49330 33552 49386 33561
rect 49330 33487 49386 33496
rect 48780 33040 48832 33046
rect 48780 32982 48832 32988
rect 47950 32668 48258 32677
rect 47950 32666 47956 32668
rect 48012 32666 48036 32668
rect 48092 32666 48116 32668
rect 48172 32666 48196 32668
rect 48252 32666 48258 32668
rect 48012 32614 48014 32666
rect 48194 32614 48196 32666
rect 47950 32612 47956 32614
rect 48012 32612 48036 32614
rect 48092 32612 48116 32614
rect 48172 32612 48196 32614
rect 48252 32612 48258 32614
rect 47950 32603 48258 32612
rect 48792 32434 48820 32982
rect 49332 32904 49384 32910
rect 49330 32872 49332 32881
rect 49384 32872 49386 32881
rect 49330 32807 49386 32816
rect 49148 32768 49200 32774
rect 49148 32710 49200 32716
rect 49160 32570 49188 32710
rect 49148 32564 49200 32570
rect 49148 32506 49200 32512
rect 48780 32428 48832 32434
rect 48780 32370 48832 32376
rect 48504 32360 48556 32366
rect 48504 32302 48556 32308
rect 48516 32201 48544 32302
rect 48502 32192 48558 32201
rect 48502 32127 48558 32136
rect 48504 31816 48556 31822
rect 48504 31758 48556 31764
rect 47950 31580 48258 31589
rect 47950 31578 47956 31580
rect 48012 31578 48036 31580
rect 48092 31578 48116 31580
rect 48172 31578 48196 31580
rect 48252 31578 48258 31580
rect 48012 31526 48014 31578
rect 48194 31526 48196 31578
rect 47950 31524 47956 31526
rect 48012 31524 48036 31526
rect 48092 31524 48116 31526
rect 48172 31524 48196 31526
rect 48252 31524 48258 31526
rect 47950 31515 48258 31524
rect 48516 31521 48544 31758
rect 48502 31512 48558 31521
rect 47860 31476 47912 31482
rect 48502 31447 48558 31456
rect 47860 31418 47912 31424
rect 48504 31272 48556 31278
rect 48504 31214 48556 31220
rect 47676 30932 47728 30938
rect 47676 30874 47728 30880
rect 48516 30841 48544 31214
rect 48502 30832 48558 30841
rect 48502 30767 48558 30776
rect 48688 30660 48740 30666
rect 48688 30602 48740 30608
rect 47950 30492 48258 30501
rect 47950 30490 47956 30492
rect 48012 30490 48036 30492
rect 48092 30490 48116 30492
rect 48172 30490 48196 30492
rect 48252 30490 48258 30492
rect 48012 30438 48014 30490
rect 48194 30438 48196 30490
rect 47950 30436 47956 30438
rect 48012 30436 48036 30438
rect 48092 30436 48116 30438
rect 48172 30436 48196 30438
rect 48252 30436 48258 30438
rect 47950 30427 48258 30436
rect 48504 29640 48556 29646
rect 48504 29582 48556 29588
rect 48516 29481 48544 29582
rect 48502 29472 48558 29481
rect 47950 29404 48258 29413
rect 48502 29407 48558 29416
rect 47950 29402 47956 29404
rect 48012 29402 48036 29404
rect 48092 29402 48116 29404
rect 48172 29402 48196 29404
rect 48252 29402 48258 29404
rect 48012 29350 48014 29402
rect 48194 29350 48196 29402
rect 47950 29348 47956 29350
rect 48012 29348 48036 29350
rect 48092 29348 48116 29350
rect 48172 29348 48196 29350
rect 48252 29348 48258 29350
rect 47950 29339 48258 29348
rect 47950 28316 48258 28325
rect 47950 28314 47956 28316
rect 48012 28314 48036 28316
rect 48092 28314 48116 28316
rect 48172 28314 48196 28316
rect 48252 28314 48258 28316
rect 48012 28262 48014 28314
rect 48194 28262 48196 28314
rect 47950 28260 47956 28262
rect 48012 28260 48036 28262
rect 48092 28260 48116 28262
rect 48172 28260 48196 28262
rect 48252 28260 48258 28262
rect 47950 28251 48258 28260
rect 47768 27872 47820 27878
rect 47768 27814 47820 27820
rect 47584 27396 47636 27402
rect 47584 27338 47636 27344
rect 47676 27396 47728 27402
rect 47676 27338 47728 27344
rect 47596 22030 47624 27338
rect 47688 26926 47716 27338
rect 47676 26920 47728 26926
rect 47676 26862 47728 26868
rect 47676 26784 47728 26790
rect 47676 26726 47728 26732
rect 47688 23118 47716 26726
rect 47780 24206 47808 27814
rect 48504 27464 48556 27470
rect 48502 27432 48504 27441
rect 48556 27432 48558 27441
rect 48502 27367 48558 27376
rect 47950 27228 48258 27237
rect 47950 27226 47956 27228
rect 48012 27226 48036 27228
rect 48092 27226 48116 27228
rect 48172 27226 48196 27228
rect 48252 27226 48258 27228
rect 48012 27174 48014 27226
rect 48194 27174 48196 27226
rect 47950 27172 47956 27174
rect 48012 27172 48036 27174
rect 48092 27172 48116 27174
rect 48172 27172 48196 27174
rect 48252 27172 48258 27174
rect 47950 27163 48258 27172
rect 48504 26920 48556 26926
rect 48504 26862 48556 26868
rect 48516 26761 48544 26862
rect 48502 26752 48558 26761
rect 48502 26687 48558 26696
rect 48228 26376 48280 26382
rect 48228 26318 48280 26324
rect 48240 26234 48268 26318
rect 48240 26206 48360 26234
rect 47950 26140 48258 26149
rect 47950 26138 47956 26140
rect 48012 26138 48036 26140
rect 48092 26138 48116 26140
rect 48172 26138 48196 26140
rect 48252 26138 48258 26140
rect 48012 26086 48014 26138
rect 48194 26086 48196 26138
rect 47950 26084 47956 26086
rect 48012 26084 48036 26086
rect 48092 26084 48116 26086
rect 48172 26084 48196 26086
rect 48252 26084 48258 26086
rect 47950 26075 48258 26084
rect 48332 26058 48360 26206
rect 48410 26072 48466 26081
rect 48332 26030 48410 26058
rect 48410 26007 48466 26016
rect 47860 25220 47912 25226
rect 47860 25162 47912 25168
rect 47768 24200 47820 24206
rect 47768 24142 47820 24148
rect 47676 23112 47728 23118
rect 47676 23054 47728 23060
rect 47584 22024 47636 22030
rect 47584 21966 47636 21972
rect 47872 20466 47900 25162
rect 47950 25052 48258 25061
rect 47950 25050 47956 25052
rect 48012 25050 48036 25052
rect 48092 25050 48116 25052
rect 48172 25050 48196 25052
rect 48252 25050 48258 25052
rect 48012 24998 48014 25050
rect 48194 24998 48196 25050
rect 47950 24996 47956 24998
rect 48012 24996 48036 24998
rect 48092 24996 48116 24998
rect 48172 24996 48196 24998
rect 48252 24996 48258 24998
rect 47950 24987 48258 24996
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47860 20460 47912 20466
rect 47860 20402 47912 20408
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47860 18692 47912 18698
rect 47860 18634 47912 18640
rect 47872 16114 47900 18634
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 48700 16574 48728 30602
rect 49332 30252 49384 30258
rect 49332 30194 49384 30200
rect 49344 30161 49372 30194
rect 49330 30152 49386 30161
rect 49330 30087 49386 30096
rect 49332 29164 49384 29170
rect 49332 29106 49384 29112
rect 49344 28801 49372 29106
rect 49330 28792 49386 28801
rect 49330 28727 49386 28736
rect 49332 28552 49384 28558
rect 49332 28494 49384 28500
rect 49344 28121 49372 28494
rect 49330 28112 49386 28121
rect 49330 28047 49386 28056
rect 48780 27124 48832 27130
rect 48780 27066 48832 27072
rect 48792 26450 48820 27066
rect 48780 26444 48832 26450
rect 48780 26386 48832 26392
rect 49332 25900 49384 25906
rect 49332 25842 49384 25848
rect 49148 25696 49200 25702
rect 49148 25638 49200 25644
rect 49160 25498 49188 25638
rect 49148 25492 49200 25498
rect 49148 25434 49200 25440
rect 49344 25401 49372 25842
rect 49330 25392 49386 25401
rect 49330 25327 49386 25336
rect 49148 24744 49200 24750
rect 49146 24712 49148 24721
rect 49200 24712 49202 24721
rect 49146 24647 49202 24656
rect 49148 24132 49200 24138
rect 49148 24074 49200 24080
rect 49160 24041 49188 24074
rect 49146 24032 49202 24041
rect 49146 23967 49202 23976
rect 49148 23656 49200 23662
rect 49148 23598 49200 23604
rect 49160 23361 49188 23598
rect 49146 23352 49202 23361
rect 49146 23287 49202 23296
rect 49148 23044 49200 23050
rect 49148 22986 49200 22992
rect 49160 22681 49188 22986
rect 49146 22672 49202 22681
rect 49146 22607 49202 22616
rect 49148 22024 49200 22030
rect 49146 21992 49148 22001
rect 49200 21992 49202 22001
rect 49146 21927 49202 21936
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21321 49188 21422
rect 49146 21312 49202 21321
rect 49146 21247 49202 21256
rect 49148 20868 49200 20874
rect 49148 20810 49200 20816
rect 49160 20641 49188 20810
rect 49146 20632 49202 20641
rect 49146 20567 49202 20576
rect 49148 20392 49200 20398
rect 49148 20334 49200 20340
rect 49160 19961 49188 20334
rect 49146 19952 49202 19961
rect 49146 19887 49202 19896
rect 49148 19372 49200 19378
rect 49148 19314 49200 19320
rect 49160 19281 49188 19314
rect 49146 19272 49202 19281
rect 49146 19207 49202 19216
rect 49148 18692 49200 18698
rect 49148 18634 49200 18640
rect 49160 18601 49188 18634
rect 49146 18592 49202 18601
rect 49146 18527 49202 18536
rect 49148 18216 49200 18222
rect 49148 18158 49200 18164
rect 49160 17921 49188 18158
rect 49146 17912 49202 17921
rect 49146 17847 49202 17856
rect 49148 17604 49200 17610
rect 49148 17546 49200 17552
rect 49160 17241 49188 17546
rect 49146 17232 49202 17241
rect 49146 17167 49202 17176
rect 48700 16546 48820 16574
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47860 16108 47912 16114
rect 47860 16050 47912 16056
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 47780 6914 47808 10610
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 47860 9376 47912 9382
rect 47860 9318 47912 9324
rect 47872 7410 47900 9318
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 47860 7404 47912 7410
rect 47860 7346 47912 7352
rect 47780 6886 47900 6914
rect 47400 6792 47452 6798
rect 47400 6734 47452 6740
rect 46204 5704 46256 5710
rect 46204 5646 46256 5652
rect 46020 4140 46072 4146
rect 46020 4082 46072 4088
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 46032 2650 46060 4082
rect 47412 3058 47440 6734
rect 47492 6656 47544 6662
rect 47492 6598 47544 6604
rect 47504 3058 47532 6598
rect 47872 5030 47900 6886
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 48792 6322 48820 16546
rect 49146 16552 49202 16561
rect 49146 16487 49148 16496
rect 49200 16487 49202 16496
rect 49148 16458 49200 16464
rect 49148 16040 49200 16046
rect 49148 15982 49200 15988
rect 49160 15881 49188 15982
rect 49146 15872 49202 15881
rect 49146 15807 49202 15816
rect 49148 15428 49200 15434
rect 49148 15370 49200 15376
rect 49160 15201 49188 15370
rect 49146 15192 49202 15201
rect 49146 15127 49202 15136
rect 49148 14952 49200 14958
rect 49148 14894 49200 14900
rect 49160 14521 49188 14894
rect 49146 14512 49202 14521
rect 49146 14447 49202 14456
rect 49148 13864 49200 13870
rect 49146 13832 49148 13841
rect 49200 13832 49202 13841
rect 49146 13767 49202 13776
rect 49148 13252 49200 13258
rect 49148 13194 49200 13200
rect 49160 13161 49188 13194
rect 49146 13152 49202 13161
rect 49146 13087 49202 13096
rect 49148 12776 49200 12782
rect 49148 12718 49200 12724
rect 49160 12481 49188 12718
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49148 12164 49200 12170
rect 49148 12106 49200 12112
rect 49160 11801 49188 12106
rect 49146 11792 49202 11801
rect 49146 11727 49202 11736
rect 49148 11144 49200 11150
rect 49146 11112 49148 11121
rect 49200 11112 49202 11121
rect 49146 11047 49202 11056
rect 49148 10600 49200 10606
rect 49148 10542 49200 10548
rect 49160 10441 49188 10542
rect 49146 10432 49202 10441
rect 49146 10367 49202 10376
rect 49148 9988 49200 9994
rect 49148 9930 49200 9936
rect 49160 9761 49188 9930
rect 49146 9752 49202 9761
rect 49146 9687 49202 9696
rect 49148 9512 49200 9518
rect 49148 9454 49200 9460
rect 49160 9081 49188 9454
rect 49146 9072 49202 9081
rect 49146 9007 49202 9016
rect 49148 8424 49200 8430
rect 49146 8392 49148 8401
rect 49200 8392 49202 8401
rect 49146 8327 49202 8336
rect 49148 7812 49200 7818
rect 49148 7754 49200 7760
rect 49160 7721 49188 7754
rect 49146 7712 49202 7721
rect 49146 7647 49202 7656
rect 49148 7336 49200 7342
rect 49148 7278 49200 7284
rect 49160 7041 49188 7278
rect 49146 7032 49202 7041
rect 49146 6967 49202 6976
rect 49148 6724 49200 6730
rect 49148 6666 49200 6672
rect 49160 6361 49188 6666
rect 49146 6352 49202 6361
rect 48780 6316 48832 6322
rect 49146 6287 49202 6296
rect 48780 6258 48832 6264
rect 48320 6112 48372 6118
rect 48320 6054 48372 6060
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 47860 5024 47912 5030
rect 47860 4966 47912 4972
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47400 3052 47452 3058
rect 47400 2994 47452 3000
rect 47492 3052 47544 3058
rect 47492 2994 47544 3000
rect 47124 2984 47176 2990
rect 47124 2926 47176 2932
rect 46388 2848 46440 2854
rect 46388 2790 46440 2796
rect 46020 2644 46072 2650
rect 46020 2586 46072 2592
rect 45652 2372 45704 2378
rect 45652 2314 45704 2320
rect 45664 800 45692 2314
rect 46400 800 46428 2790
rect 47136 800 47164 2926
rect 47780 2446 47808 3878
rect 48332 3534 48360 6054
rect 48792 4146 48820 6258
rect 49148 5704 49200 5710
rect 49146 5672 49148 5681
rect 49200 5672 49202 5681
rect 49146 5607 49202 5616
rect 49332 5024 49384 5030
rect 49330 4992 49332 5001
rect 49384 4992 49386 5001
rect 49330 4927 49386 4936
rect 49148 4548 49200 4554
rect 49148 4490 49200 4496
rect 49160 4321 49188 4490
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 48780 4140 48832 4146
rect 48780 4082 48832 4088
rect 48596 4072 48648 4078
rect 48596 4014 48648 4020
rect 48320 3528 48372 3534
rect 48320 3470 48372 3476
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 47860 2984 47912 2990
rect 47860 2926 47912 2932
rect 47768 2440 47820 2446
rect 47768 2382 47820 2388
rect 47872 800 47900 2926
rect 48320 2848 48372 2854
rect 48320 2790 48372 2796
rect 48332 2514 48360 2790
rect 48320 2508 48372 2514
rect 48320 2450 48372 2456
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 48608 800 48636 4014
rect 49332 3460 49384 3466
rect 49332 3402 49384 3408
rect 49344 800 49372 3402
rect 28092 734 28396 762
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 30930 0 30986 800
rect 31666 0 31722 800
rect 32402 0 32458 800
rect 33138 0 33194 800
rect 33874 0 33930 800
rect 34610 0 34666 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37554 0 37610 800
rect 38290 0 38346 800
rect 39026 0 39082 800
rect 39762 0 39818 800
rect 40498 0 40554 800
rect 41234 0 41290 800
rect 41970 0 42026 800
rect 42706 0 42762 800
rect 43442 0 43498 800
rect 44178 0 44234 800
rect 44914 0 44970 800
rect 45650 0 45706 800
rect 46386 0 46442 800
rect 47122 0 47178 800
rect 47858 0 47914 800
rect 48594 0 48650 800
rect 49330 0 49386 800
<< via2 >>
rect 938 52672 994 52728
rect 2778 54984 2834 55040
rect 938 50360 994 50416
rect 938 48068 994 48104
rect 938 48048 940 48068
rect 940 48048 992 48068
rect 992 48048 994 48068
rect 938 45736 994 45792
rect 1674 41112 1730 41168
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 938 38800 994 38856
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 938 36488 994 36544
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 1766 34176 1822 34232
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 938 31864 994 31920
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 1306 29552 1362 29608
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 1306 27240 1362 27296
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 1306 24928 1362 24984
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 9770 31320 9826 31376
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 8942 24928 8998 24984
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 1306 22616 1362 22672
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 1306 20340 1308 20360
rect 1308 20340 1360 20360
rect 1360 20340 1362 20360
rect 1306 20304 1362 20340
rect 1306 17992 1362 18048
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 1306 15680 1362 15736
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2778 13368 2834 13424
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 3422 11056 3478 11112
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3330 8744 3386 8800
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3422 6432 3478 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3422 4120 3478 4176
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2778 1808 2834 1864
rect 5446 2916 5502 2952
rect 5446 2896 5448 2916
rect 5448 2896 5500 2916
rect 5500 2896 5502 2916
rect 5998 2372 6054 2408
rect 5998 2352 6000 2372
rect 6000 2352 6052 2372
rect 6052 2352 6054 2372
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 9494 25200 9550 25256
rect 9494 24928 9550 24984
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 9586 22616 9642 22672
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12346 2488 12402 2544
rect 11150 1808 11206 1864
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17038 35128 17094 35184
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 27956 54426 28012 54428
rect 28036 54426 28092 54428
rect 28116 54426 28172 54428
rect 28196 54426 28252 54428
rect 27956 54374 28002 54426
rect 28002 54374 28012 54426
rect 28036 54374 28066 54426
rect 28066 54374 28078 54426
rect 28078 54374 28092 54426
rect 28116 54374 28130 54426
rect 28130 54374 28142 54426
rect 28142 54374 28172 54426
rect 28196 54374 28206 54426
rect 28206 54374 28252 54426
rect 27956 54372 28012 54374
rect 28036 54372 28092 54374
rect 28116 54372 28172 54374
rect 28196 54372 28252 54374
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22466 34992 22522 35048
rect 21270 33360 21326 33416
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17958 3032 18014 3088
rect 15290 1944 15346 2000
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 23294 37204 23296 37224
rect 23296 37204 23348 37224
rect 23348 37204 23350 37224
rect 23294 37168 23350 37204
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22742 35128 22798 35184
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22466 31220 22468 31240
rect 22468 31220 22520 31240
rect 22520 31220 22522 31240
rect 22466 31184 22522 31220
rect 22098 30796 22154 30832
rect 22098 30776 22100 30796
rect 22100 30776 22152 30796
rect 22152 30776 22154 30796
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 23294 29164 23350 29200
rect 23294 29144 23296 29164
rect 23296 29144 23348 29164
rect 23348 29144 23350 29164
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 23846 28076 23902 28112
rect 23846 28056 23848 28076
rect 23848 28056 23900 28076
rect 23900 28056 23902 28076
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24858 23432 24914 23488
rect 25042 22924 25044 22944
rect 25044 22924 25096 22944
rect 25096 22924 25098 22944
rect 25042 22888 25098 22924
rect 27956 53338 28012 53340
rect 28036 53338 28092 53340
rect 28116 53338 28172 53340
rect 28196 53338 28252 53340
rect 27956 53286 28002 53338
rect 28002 53286 28012 53338
rect 28036 53286 28066 53338
rect 28066 53286 28078 53338
rect 28078 53286 28092 53338
rect 28116 53286 28130 53338
rect 28130 53286 28142 53338
rect 28142 53286 28172 53338
rect 28196 53286 28206 53338
rect 28206 53286 28252 53338
rect 27956 53284 28012 53286
rect 28036 53284 28092 53286
rect 28116 53284 28172 53286
rect 28196 53284 28252 53286
rect 27956 52250 28012 52252
rect 28036 52250 28092 52252
rect 28116 52250 28172 52252
rect 28196 52250 28252 52252
rect 27956 52198 28002 52250
rect 28002 52198 28012 52250
rect 28036 52198 28066 52250
rect 28066 52198 28078 52250
rect 28078 52198 28092 52250
rect 28116 52198 28130 52250
rect 28130 52198 28142 52250
rect 28142 52198 28172 52250
rect 28196 52198 28206 52250
rect 28206 52198 28252 52250
rect 27956 52196 28012 52198
rect 28036 52196 28092 52198
rect 28116 52196 28172 52198
rect 28196 52196 28252 52198
rect 27956 51162 28012 51164
rect 28036 51162 28092 51164
rect 28116 51162 28172 51164
rect 28196 51162 28252 51164
rect 27956 51110 28002 51162
rect 28002 51110 28012 51162
rect 28036 51110 28066 51162
rect 28066 51110 28078 51162
rect 28078 51110 28092 51162
rect 28116 51110 28130 51162
rect 28130 51110 28142 51162
rect 28142 51110 28172 51162
rect 28196 51110 28206 51162
rect 28206 51110 28252 51162
rect 27956 51108 28012 51110
rect 28036 51108 28092 51110
rect 28116 51108 28172 51110
rect 28196 51108 28252 51110
rect 27956 50074 28012 50076
rect 28036 50074 28092 50076
rect 28116 50074 28172 50076
rect 28196 50074 28252 50076
rect 27956 50022 28002 50074
rect 28002 50022 28012 50074
rect 28036 50022 28066 50074
rect 28066 50022 28078 50074
rect 28078 50022 28092 50074
rect 28116 50022 28130 50074
rect 28130 50022 28142 50074
rect 28142 50022 28172 50074
rect 28196 50022 28206 50074
rect 28206 50022 28252 50074
rect 27956 50020 28012 50022
rect 28036 50020 28092 50022
rect 28116 50020 28172 50022
rect 28196 50020 28252 50022
rect 27956 48986 28012 48988
rect 28036 48986 28092 48988
rect 28116 48986 28172 48988
rect 28196 48986 28252 48988
rect 27956 48934 28002 48986
rect 28002 48934 28012 48986
rect 28036 48934 28066 48986
rect 28066 48934 28078 48986
rect 28078 48934 28092 48986
rect 28116 48934 28130 48986
rect 28130 48934 28142 48986
rect 28142 48934 28172 48986
rect 28196 48934 28206 48986
rect 28206 48934 28252 48986
rect 27956 48932 28012 48934
rect 28036 48932 28092 48934
rect 28116 48932 28172 48934
rect 28196 48932 28252 48934
rect 27956 47898 28012 47900
rect 28036 47898 28092 47900
rect 28116 47898 28172 47900
rect 28196 47898 28252 47900
rect 27956 47846 28002 47898
rect 28002 47846 28012 47898
rect 28036 47846 28066 47898
rect 28066 47846 28078 47898
rect 28078 47846 28092 47898
rect 28116 47846 28130 47898
rect 28130 47846 28142 47898
rect 28142 47846 28172 47898
rect 28196 47846 28206 47898
rect 28206 47846 28252 47898
rect 27956 47844 28012 47846
rect 28036 47844 28092 47846
rect 28116 47844 28172 47846
rect 28196 47844 28252 47846
rect 27956 46810 28012 46812
rect 28036 46810 28092 46812
rect 28116 46810 28172 46812
rect 28196 46810 28252 46812
rect 27956 46758 28002 46810
rect 28002 46758 28012 46810
rect 28036 46758 28066 46810
rect 28066 46758 28078 46810
rect 28078 46758 28092 46810
rect 28116 46758 28130 46810
rect 28130 46758 28142 46810
rect 28142 46758 28172 46810
rect 28196 46758 28206 46810
rect 28206 46758 28252 46810
rect 27956 46756 28012 46758
rect 28036 46756 28092 46758
rect 28116 46756 28172 46758
rect 28196 46756 28252 46758
rect 26790 33360 26846 33416
rect 26790 32816 26846 32872
rect 26238 28092 26240 28112
rect 26240 28092 26292 28112
rect 26292 28092 26294 28112
rect 26238 28056 26294 28092
rect 25962 24692 25964 24712
rect 25964 24692 26016 24712
rect 26016 24692 26018 24712
rect 25962 24656 26018 24692
rect 25502 24268 25558 24304
rect 25502 24248 25504 24268
rect 25504 24248 25556 24268
rect 25556 24248 25558 24268
rect 26330 24792 26386 24848
rect 27526 40468 27528 40488
rect 27528 40468 27580 40488
rect 27580 40468 27582 40488
rect 27526 40432 27582 40468
rect 27956 45722 28012 45724
rect 28036 45722 28092 45724
rect 28116 45722 28172 45724
rect 28196 45722 28252 45724
rect 27956 45670 28002 45722
rect 28002 45670 28012 45722
rect 28036 45670 28066 45722
rect 28066 45670 28078 45722
rect 28078 45670 28092 45722
rect 28116 45670 28130 45722
rect 28130 45670 28142 45722
rect 28142 45670 28172 45722
rect 28196 45670 28206 45722
rect 28206 45670 28252 45722
rect 27956 45668 28012 45670
rect 28036 45668 28092 45670
rect 28116 45668 28172 45670
rect 28196 45668 28252 45670
rect 27956 44634 28012 44636
rect 28036 44634 28092 44636
rect 28116 44634 28172 44636
rect 28196 44634 28252 44636
rect 27956 44582 28002 44634
rect 28002 44582 28012 44634
rect 28036 44582 28066 44634
rect 28066 44582 28078 44634
rect 28078 44582 28092 44634
rect 28116 44582 28130 44634
rect 28130 44582 28142 44634
rect 28142 44582 28172 44634
rect 28196 44582 28206 44634
rect 28206 44582 28252 44634
rect 27956 44580 28012 44582
rect 28036 44580 28092 44582
rect 28116 44580 28172 44582
rect 28196 44580 28252 44582
rect 27956 43546 28012 43548
rect 28036 43546 28092 43548
rect 28116 43546 28172 43548
rect 28196 43546 28252 43548
rect 27956 43494 28002 43546
rect 28002 43494 28012 43546
rect 28036 43494 28066 43546
rect 28066 43494 28078 43546
rect 28078 43494 28092 43546
rect 28116 43494 28130 43546
rect 28130 43494 28142 43546
rect 28142 43494 28172 43546
rect 28196 43494 28206 43546
rect 28206 43494 28252 43546
rect 27956 43492 28012 43494
rect 28036 43492 28092 43494
rect 28116 43492 28172 43494
rect 28196 43492 28252 43494
rect 27956 42458 28012 42460
rect 28036 42458 28092 42460
rect 28116 42458 28172 42460
rect 28196 42458 28252 42460
rect 27956 42406 28002 42458
rect 28002 42406 28012 42458
rect 28036 42406 28066 42458
rect 28066 42406 28078 42458
rect 28078 42406 28092 42458
rect 28116 42406 28130 42458
rect 28130 42406 28142 42458
rect 28142 42406 28172 42458
rect 28196 42406 28206 42458
rect 28206 42406 28252 42458
rect 27956 42404 28012 42406
rect 28036 42404 28092 42406
rect 28116 42404 28172 42406
rect 28196 42404 28252 42406
rect 27956 41370 28012 41372
rect 28036 41370 28092 41372
rect 28116 41370 28172 41372
rect 28196 41370 28252 41372
rect 27956 41318 28002 41370
rect 28002 41318 28012 41370
rect 28036 41318 28066 41370
rect 28066 41318 28078 41370
rect 28078 41318 28092 41370
rect 28116 41318 28130 41370
rect 28130 41318 28142 41370
rect 28142 41318 28172 41370
rect 28196 41318 28206 41370
rect 28206 41318 28252 41370
rect 27956 41316 28012 41318
rect 28036 41316 28092 41318
rect 28116 41316 28172 41318
rect 28196 41316 28252 41318
rect 27956 40282 28012 40284
rect 28036 40282 28092 40284
rect 28116 40282 28172 40284
rect 28196 40282 28252 40284
rect 27956 40230 28002 40282
rect 28002 40230 28012 40282
rect 28036 40230 28066 40282
rect 28066 40230 28078 40282
rect 28078 40230 28092 40282
rect 28116 40230 28130 40282
rect 28130 40230 28142 40282
rect 28142 40230 28172 40282
rect 28196 40230 28206 40282
rect 28206 40230 28252 40282
rect 27956 40228 28012 40230
rect 28036 40228 28092 40230
rect 28116 40228 28172 40230
rect 28196 40228 28252 40230
rect 27956 39194 28012 39196
rect 28036 39194 28092 39196
rect 28116 39194 28172 39196
rect 28196 39194 28252 39196
rect 27956 39142 28002 39194
rect 28002 39142 28012 39194
rect 28036 39142 28066 39194
rect 28066 39142 28078 39194
rect 28078 39142 28092 39194
rect 28116 39142 28130 39194
rect 28130 39142 28142 39194
rect 28142 39142 28172 39194
rect 28196 39142 28206 39194
rect 28206 39142 28252 39194
rect 27956 39140 28012 39142
rect 28036 39140 28092 39142
rect 28116 39140 28172 39142
rect 28196 39140 28252 39142
rect 27956 38106 28012 38108
rect 28036 38106 28092 38108
rect 28116 38106 28172 38108
rect 28196 38106 28252 38108
rect 27956 38054 28002 38106
rect 28002 38054 28012 38106
rect 28036 38054 28066 38106
rect 28066 38054 28078 38106
rect 28078 38054 28092 38106
rect 28116 38054 28130 38106
rect 28130 38054 28142 38106
rect 28142 38054 28172 38106
rect 28196 38054 28206 38106
rect 28206 38054 28252 38106
rect 27956 38052 28012 38054
rect 28036 38052 28092 38054
rect 28116 38052 28172 38054
rect 28196 38052 28252 38054
rect 27956 37018 28012 37020
rect 28036 37018 28092 37020
rect 28116 37018 28172 37020
rect 28196 37018 28252 37020
rect 27956 36966 28002 37018
rect 28002 36966 28012 37018
rect 28036 36966 28066 37018
rect 28066 36966 28078 37018
rect 28078 36966 28092 37018
rect 28116 36966 28130 37018
rect 28130 36966 28142 37018
rect 28142 36966 28172 37018
rect 28196 36966 28206 37018
rect 28206 36966 28252 37018
rect 27956 36964 28012 36966
rect 28036 36964 28092 36966
rect 28116 36964 28172 36966
rect 28196 36964 28252 36966
rect 27956 35930 28012 35932
rect 28036 35930 28092 35932
rect 28116 35930 28172 35932
rect 28196 35930 28252 35932
rect 27956 35878 28002 35930
rect 28002 35878 28012 35930
rect 28036 35878 28066 35930
rect 28066 35878 28078 35930
rect 28078 35878 28092 35930
rect 28116 35878 28130 35930
rect 28130 35878 28142 35930
rect 28142 35878 28172 35930
rect 28196 35878 28206 35930
rect 28206 35878 28252 35930
rect 27956 35876 28012 35878
rect 28036 35876 28092 35878
rect 28116 35876 28172 35878
rect 28196 35876 28252 35878
rect 27710 35672 27766 35728
rect 27956 34842 28012 34844
rect 28036 34842 28092 34844
rect 28116 34842 28172 34844
rect 28196 34842 28252 34844
rect 27956 34790 28002 34842
rect 28002 34790 28012 34842
rect 28036 34790 28066 34842
rect 28066 34790 28078 34842
rect 28078 34790 28092 34842
rect 28116 34790 28130 34842
rect 28130 34790 28142 34842
rect 28142 34790 28172 34842
rect 28196 34790 28206 34842
rect 28206 34790 28252 34842
rect 27956 34788 28012 34790
rect 28036 34788 28092 34790
rect 28116 34788 28172 34790
rect 28196 34788 28252 34790
rect 28262 34584 28318 34640
rect 27956 33754 28012 33756
rect 28036 33754 28092 33756
rect 28116 33754 28172 33756
rect 28196 33754 28252 33756
rect 27956 33702 28002 33754
rect 28002 33702 28012 33754
rect 28036 33702 28066 33754
rect 28066 33702 28078 33754
rect 28078 33702 28092 33754
rect 28116 33702 28130 33754
rect 28130 33702 28142 33754
rect 28142 33702 28172 33754
rect 28196 33702 28206 33754
rect 28206 33702 28252 33754
rect 27956 33700 28012 33702
rect 28036 33700 28092 33702
rect 28116 33700 28172 33702
rect 28196 33700 28252 33702
rect 27956 32666 28012 32668
rect 28036 32666 28092 32668
rect 28116 32666 28172 32668
rect 28196 32666 28252 32668
rect 27956 32614 28002 32666
rect 28002 32614 28012 32666
rect 28036 32614 28066 32666
rect 28066 32614 28078 32666
rect 28078 32614 28092 32666
rect 28116 32614 28130 32666
rect 28130 32614 28142 32666
rect 28142 32614 28172 32666
rect 28196 32614 28206 32666
rect 28206 32614 28252 32666
rect 27956 32612 28012 32614
rect 28036 32612 28092 32614
rect 28116 32612 28172 32614
rect 28196 32612 28252 32614
rect 27250 19216 27306 19272
rect 27956 31578 28012 31580
rect 28036 31578 28092 31580
rect 28116 31578 28172 31580
rect 28196 31578 28252 31580
rect 27956 31526 28002 31578
rect 28002 31526 28012 31578
rect 28036 31526 28066 31578
rect 28066 31526 28078 31578
rect 28078 31526 28092 31578
rect 28116 31526 28130 31578
rect 28130 31526 28142 31578
rect 28142 31526 28172 31578
rect 28196 31526 28206 31578
rect 28206 31526 28252 31578
rect 27956 31524 28012 31526
rect 28036 31524 28092 31526
rect 28116 31524 28172 31526
rect 28196 31524 28252 31526
rect 27956 30490 28012 30492
rect 28036 30490 28092 30492
rect 28116 30490 28172 30492
rect 28196 30490 28252 30492
rect 27956 30438 28002 30490
rect 28002 30438 28012 30490
rect 28036 30438 28066 30490
rect 28066 30438 28078 30490
rect 28078 30438 28092 30490
rect 28116 30438 28130 30490
rect 28130 30438 28142 30490
rect 28142 30438 28172 30490
rect 28196 30438 28206 30490
rect 28206 30438 28252 30490
rect 27956 30436 28012 30438
rect 28036 30436 28092 30438
rect 28116 30436 28172 30438
rect 28196 30436 28252 30438
rect 27956 29402 28012 29404
rect 28036 29402 28092 29404
rect 28116 29402 28172 29404
rect 28196 29402 28252 29404
rect 27956 29350 28002 29402
rect 28002 29350 28012 29402
rect 28036 29350 28066 29402
rect 28066 29350 28078 29402
rect 28078 29350 28092 29402
rect 28116 29350 28130 29402
rect 28130 29350 28142 29402
rect 28142 29350 28172 29402
rect 28196 29350 28206 29402
rect 28206 29350 28252 29402
rect 27956 29348 28012 29350
rect 28036 29348 28092 29350
rect 28116 29348 28172 29350
rect 28196 29348 28252 29350
rect 27956 28314 28012 28316
rect 28036 28314 28092 28316
rect 28116 28314 28172 28316
rect 28196 28314 28252 28316
rect 27956 28262 28002 28314
rect 28002 28262 28012 28314
rect 28036 28262 28066 28314
rect 28066 28262 28078 28314
rect 28078 28262 28092 28314
rect 28116 28262 28130 28314
rect 28130 28262 28142 28314
rect 28142 28262 28172 28314
rect 28196 28262 28206 28314
rect 28206 28262 28252 28314
rect 27956 28260 28012 28262
rect 28036 28260 28092 28262
rect 28116 28260 28172 28262
rect 28196 28260 28252 28262
rect 28722 31628 28724 31648
rect 28724 31628 28776 31648
rect 28776 31628 28778 31648
rect 28722 31592 28778 31628
rect 28722 31456 28778 31512
rect 28722 30776 28778 30832
rect 27956 27226 28012 27228
rect 28036 27226 28092 27228
rect 28116 27226 28172 27228
rect 28196 27226 28252 27228
rect 27956 27174 28002 27226
rect 28002 27174 28012 27226
rect 28036 27174 28066 27226
rect 28066 27174 28078 27226
rect 28078 27174 28092 27226
rect 28116 27174 28130 27226
rect 28130 27174 28142 27226
rect 28142 27174 28172 27226
rect 28196 27174 28206 27226
rect 28206 27174 28252 27226
rect 27956 27172 28012 27174
rect 28036 27172 28092 27174
rect 28116 27172 28172 27174
rect 28196 27172 28252 27174
rect 27956 26138 28012 26140
rect 28036 26138 28092 26140
rect 28116 26138 28172 26140
rect 28196 26138 28252 26140
rect 27956 26086 28002 26138
rect 28002 26086 28012 26138
rect 28036 26086 28066 26138
rect 28066 26086 28078 26138
rect 28078 26086 28092 26138
rect 28116 26086 28130 26138
rect 28130 26086 28142 26138
rect 28142 26086 28172 26138
rect 28196 26086 28206 26138
rect 28206 26086 28252 26138
rect 27956 26084 28012 26086
rect 28036 26084 28092 26086
rect 28116 26084 28172 26086
rect 28196 26084 28252 26086
rect 27956 25050 28012 25052
rect 28036 25050 28092 25052
rect 28116 25050 28172 25052
rect 28196 25050 28252 25052
rect 27956 24998 28002 25050
rect 28002 24998 28012 25050
rect 28036 24998 28066 25050
rect 28066 24998 28078 25050
rect 28078 24998 28092 25050
rect 28116 24998 28130 25050
rect 28130 24998 28142 25050
rect 28142 24998 28172 25050
rect 28196 24998 28206 25050
rect 28206 24998 28252 25050
rect 27956 24996 28012 24998
rect 28036 24996 28092 24998
rect 28116 24996 28172 24998
rect 28196 24996 28252 24998
rect 27894 24828 27896 24848
rect 27896 24828 27948 24848
rect 27948 24828 27950 24848
rect 27894 24792 27950 24828
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27710 18672 27766 18728
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 28538 27512 28594 27568
rect 28538 24792 28594 24848
rect 32956 53882 33012 53884
rect 33036 53882 33092 53884
rect 33116 53882 33172 53884
rect 33196 53882 33252 53884
rect 32956 53830 33002 53882
rect 33002 53830 33012 53882
rect 33036 53830 33066 53882
rect 33066 53830 33078 53882
rect 33078 53830 33092 53882
rect 33116 53830 33130 53882
rect 33130 53830 33142 53882
rect 33142 53830 33172 53882
rect 33196 53830 33206 53882
rect 33206 53830 33252 53882
rect 32956 53828 33012 53830
rect 33036 53828 33092 53830
rect 33116 53828 33172 53830
rect 33196 53828 33252 53830
rect 32956 52794 33012 52796
rect 33036 52794 33092 52796
rect 33116 52794 33172 52796
rect 33196 52794 33252 52796
rect 32956 52742 33002 52794
rect 33002 52742 33012 52794
rect 33036 52742 33066 52794
rect 33066 52742 33078 52794
rect 33078 52742 33092 52794
rect 33116 52742 33130 52794
rect 33130 52742 33142 52794
rect 33142 52742 33172 52794
rect 33196 52742 33206 52794
rect 33206 52742 33252 52794
rect 32956 52740 33012 52742
rect 33036 52740 33092 52742
rect 33116 52740 33172 52742
rect 33196 52740 33252 52742
rect 32956 51706 33012 51708
rect 33036 51706 33092 51708
rect 33116 51706 33172 51708
rect 33196 51706 33252 51708
rect 32956 51654 33002 51706
rect 33002 51654 33012 51706
rect 33036 51654 33066 51706
rect 33066 51654 33078 51706
rect 33078 51654 33092 51706
rect 33116 51654 33130 51706
rect 33130 51654 33142 51706
rect 33142 51654 33172 51706
rect 33196 51654 33206 51706
rect 33206 51654 33252 51706
rect 32956 51652 33012 51654
rect 33036 51652 33092 51654
rect 33116 51652 33172 51654
rect 33196 51652 33252 51654
rect 32956 50618 33012 50620
rect 33036 50618 33092 50620
rect 33116 50618 33172 50620
rect 33196 50618 33252 50620
rect 32956 50566 33002 50618
rect 33002 50566 33012 50618
rect 33036 50566 33066 50618
rect 33066 50566 33078 50618
rect 33078 50566 33092 50618
rect 33116 50566 33130 50618
rect 33130 50566 33142 50618
rect 33142 50566 33172 50618
rect 33196 50566 33206 50618
rect 33206 50566 33252 50618
rect 32956 50564 33012 50566
rect 33036 50564 33092 50566
rect 33116 50564 33172 50566
rect 33196 50564 33252 50566
rect 32956 49530 33012 49532
rect 33036 49530 33092 49532
rect 33116 49530 33172 49532
rect 33196 49530 33252 49532
rect 32956 49478 33002 49530
rect 33002 49478 33012 49530
rect 33036 49478 33066 49530
rect 33066 49478 33078 49530
rect 33078 49478 33092 49530
rect 33116 49478 33130 49530
rect 33130 49478 33142 49530
rect 33142 49478 33172 49530
rect 33196 49478 33206 49530
rect 33206 49478 33252 49530
rect 32956 49476 33012 49478
rect 33036 49476 33092 49478
rect 33116 49476 33172 49478
rect 33196 49476 33252 49478
rect 32956 48442 33012 48444
rect 33036 48442 33092 48444
rect 33116 48442 33172 48444
rect 33196 48442 33252 48444
rect 32956 48390 33002 48442
rect 33002 48390 33012 48442
rect 33036 48390 33066 48442
rect 33066 48390 33078 48442
rect 33078 48390 33092 48442
rect 33116 48390 33130 48442
rect 33130 48390 33142 48442
rect 33142 48390 33172 48442
rect 33196 48390 33206 48442
rect 33206 48390 33252 48442
rect 32956 48388 33012 48390
rect 33036 48388 33092 48390
rect 33116 48388 33172 48390
rect 33196 48388 33252 48390
rect 32956 47354 33012 47356
rect 33036 47354 33092 47356
rect 33116 47354 33172 47356
rect 33196 47354 33252 47356
rect 32956 47302 33002 47354
rect 33002 47302 33012 47354
rect 33036 47302 33066 47354
rect 33066 47302 33078 47354
rect 33078 47302 33092 47354
rect 33116 47302 33130 47354
rect 33130 47302 33142 47354
rect 33142 47302 33172 47354
rect 33196 47302 33206 47354
rect 33206 47302 33252 47354
rect 32956 47300 33012 47302
rect 33036 47300 33092 47302
rect 33116 47300 33172 47302
rect 33196 47300 33252 47302
rect 32956 46266 33012 46268
rect 33036 46266 33092 46268
rect 33116 46266 33172 46268
rect 33196 46266 33252 46268
rect 32956 46214 33002 46266
rect 33002 46214 33012 46266
rect 33036 46214 33066 46266
rect 33066 46214 33078 46266
rect 33078 46214 33092 46266
rect 33116 46214 33130 46266
rect 33130 46214 33142 46266
rect 33142 46214 33172 46266
rect 33196 46214 33206 46266
rect 33206 46214 33252 46266
rect 32956 46212 33012 46214
rect 33036 46212 33092 46214
rect 33116 46212 33172 46214
rect 33196 46212 33252 46214
rect 29826 37168 29882 37224
rect 30102 35536 30158 35592
rect 28814 23432 28870 23488
rect 27710 17076 27712 17096
rect 27712 17076 27764 17096
rect 27764 17076 27766 17096
rect 27710 17040 27766 17076
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27894 18028 27896 18048
rect 27896 18028 27948 18048
rect 27948 18028 27950 18048
rect 27894 17992 27950 18028
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27986 15564 28042 15600
rect 27986 15544 27988 15564
rect 27988 15544 28040 15564
rect 28040 15544 28042 15564
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 28722 18828 28778 18864
rect 28722 18808 28724 18828
rect 28724 18808 28776 18828
rect 28776 18808 28778 18828
rect 28814 15544 28870 15600
rect 28906 12824 28962 12880
rect 30010 29008 30066 29064
rect 30654 40432 30710 40488
rect 30378 34856 30434 34912
rect 30470 29044 30472 29064
rect 30472 29044 30524 29064
rect 30524 29044 30526 29064
rect 30470 29008 30526 29044
rect 30838 37848 30894 37904
rect 30746 35128 30802 35184
rect 31850 36252 31852 36272
rect 31852 36252 31904 36272
rect 31904 36252 31906 36272
rect 31850 36216 31906 36252
rect 31298 35128 31354 35184
rect 31206 34992 31262 35048
rect 31390 35028 31392 35048
rect 31392 35028 31444 35048
rect 31444 35028 31446 35048
rect 31390 34992 31446 35028
rect 31022 31184 31078 31240
rect 31206 29144 31262 29200
rect 31022 27512 31078 27568
rect 30102 23432 30158 23488
rect 30470 22652 30472 22672
rect 30472 22652 30524 22672
rect 30524 22652 30526 22672
rect 30470 22616 30526 22652
rect 30470 20596 30526 20632
rect 30470 20576 30472 20596
rect 30472 20576 30524 20596
rect 30524 20576 30526 20596
rect 31206 27124 31262 27160
rect 31206 27104 31208 27124
rect 31208 27104 31260 27124
rect 31260 27104 31262 27124
rect 31298 26832 31354 26888
rect 31298 19216 31354 19272
rect 32956 45178 33012 45180
rect 33036 45178 33092 45180
rect 33116 45178 33172 45180
rect 33196 45178 33252 45180
rect 32956 45126 33002 45178
rect 33002 45126 33012 45178
rect 33036 45126 33066 45178
rect 33066 45126 33078 45178
rect 33078 45126 33092 45178
rect 33116 45126 33130 45178
rect 33130 45126 33142 45178
rect 33142 45126 33172 45178
rect 33196 45126 33206 45178
rect 33206 45126 33252 45178
rect 32956 45124 33012 45126
rect 33036 45124 33092 45126
rect 33116 45124 33172 45126
rect 33196 45124 33252 45126
rect 32956 44090 33012 44092
rect 33036 44090 33092 44092
rect 33116 44090 33172 44092
rect 33196 44090 33252 44092
rect 32956 44038 33002 44090
rect 33002 44038 33012 44090
rect 33036 44038 33066 44090
rect 33066 44038 33078 44090
rect 33078 44038 33092 44090
rect 33116 44038 33130 44090
rect 33130 44038 33142 44090
rect 33142 44038 33172 44090
rect 33196 44038 33206 44090
rect 33206 44038 33252 44090
rect 32956 44036 33012 44038
rect 33036 44036 33092 44038
rect 33116 44036 33172 44038
rect 33196 44036 33252 44038
rect 32956 43002 33012 43004
rect 33036 43002 33092 43004
rect 33116 43002 33172 43004
rect 33196 43002 33252 43004
rect 32956 42950 33002 43002
rect 33002 42950 33012 43002
rect 33036 42950 33066 43002
rect 33066 42950 33078 43002
rect 33078 42950 33092 43002
rect 33116 42950 33130 43002
rect 33130 42950 33142 43002
rect 33142 42950 33172 43002
rect 33196 42950 33206 43002
rect 33206 42950 33252 43002
rect 32956 42948 33012 42950
rect 33036 42948 33092 42950
rect 33116 42948 33172 42950
rect 33196 42948 33252 42950
rect 32956 41914 33012 41916
rect 33036 41914 33092 41916
rect 33116 41914 33172 41916
rect 33196 41914 33252 41916
rect 32956 41862 33002 41914
rect 33002 41862 33012 41914
rect 33036 41862 33066 41914
rect 33066 41862 33078 41914
rect 33078 41862 33092 41914
rect 33116 41862 33130 41914
rect 33130 41862 33142 41914
rect 33142 41862 33172 41914
rect 33196 41862 33206 41914
rect 33206 41862 33252 41914
rect 32956 41860 33012 41862
rect 33036 41860 33092 41862
rect 33116 41860 33172 41862
rect 33196 41860 33252 41862
rect 32494 36080 32550 36136
rect 32402 30640 32458 30696
rect 32770 35708 32772 35728
rect 32772 35708 32824 35728
rect 32824 35708 32826 35728
rect 32770 35672 32826 35708
rect 32956 40826 33012 40828
rect 33036 40826 33092 40828
rect 33116 40826 33172 40828
rect 33196 40826 33252 40828
rect 32956 40774 33002 40826
rect 33002 40774 33012 40826
rect 33036 40774 33066 40826
rect 33066 40774 33078 40826
rect 33078 40774 33092 40826
rect 33116 40774 33130 40826
rect 33130 40774 33142 40826
rect 33142 40774 33172 40826
rect 33196 40774 33206 40826
rect 33206 40774 33252 40826
rect 32956 40772 33012 40774
rect 33036 40772 33092 40774
rect 33116 40772 33172 40774
rect 33196 40772 33252 40774
rect 32956 39738 33012 39740
rect 33036 39738 33092 39740
rect 33116 39738 33172 39740
rect 33196 39738 33252 39740
rect 32956 39686 33002 39738
rect 33002 39686 33012 39738
rect 33036 39686 33066 39738
rect 33066 39686 33078 39738
rect 33078 39686 33092 39738
rect 33116 39686 33130 39738
rect 33130 39686 33142 39738
rect 33142 39686 33172 39738
rect 33196 39686 33206 39738
rect 33206 39686 33252 39738
rect 32956 39684 33012 39686
rect 33036 39684 33092 39686
rect 33116 39684 33172 39686
rect 33196 39684 33252 39686
rect 32956 38650 33012 38652
rect 33036 38650 33092 38652
rect 33116 38650 33172 38652
rect 33196 38650 33252 38652
rect 32956 38598 33002 38650
rect 33002 38598 33012 38650
rect 33036 38598 33066 38650
rect 33066 38598 33078 38650
rect 33078 38598 33092 38650
rect 33116 38598 33130 38650
rect 33130 38598 33142 38650
rect 33142 38598 33172 38650
rect 33196 38598 33206 38650
rect 33206 38598 33252 38650
rect 32956 38596 33012 38598
rect 33036 38596 33092 38598
rect 33116 38596 33172 38598
rect 33196 38596 33252 38598
rect 32956 37562 33012 37564
rect 33036 37562 33092 37564
rect 33116 37562 33172 37564
rect 33196 37562 33252 37564
rect 32956 37510 33002 37562
rect 33002 37510 33012 37562
rect 33036 37510 33066 37562
rect 33066 37510 33078 37562
rect 33078 37510 33092 37562
rect 33116 37510 33130 37562
rect 33130 37510 33142 37562
rect 33142 37510 33172 37562
rect 33196 37510 33206 37562
rect 33206 37510 33252 37562
rect 32956 37508 33012 37510
rect 33036 37508 33092 37510
rect 33116 37508 33172 37510
rect 33196 37508 33252 37510
rect 33506 37848 33562 37904
rect 33690 37168 33746 37224
rect 32956 36474 33012 36476
rect 33036 36474 33092 36476
rect 33116 36474 33172 36476
rect 33196 36474 33252 36476
rect 32956 36422 33002 36474
rect 33002 36422 33012 36474
rect 33036 36422 33066 36474
rect 33066 36422 33078 36474
rect 33078 36422 33092 36474
rect 33116 36422 33130 36474
rect 33130 36422 33142 36474
rect 33142 36422 33172 36474
rect 33196 36422 33206 36474
rect 33206 36422 33252 36474
rect 32956 36420 33012 36422
rect 33036 36420 33092 36422
rect 33116 36420 33172 36422
rect 33196 36420 33252 36422
rect 32956 35386 33012 35388
rect 33036 35386 33092 35388
rect 33116 35386 33172 35388
rect 33196 35386 33252 35388
rect 32956 35334 33002 35386
rect 33002 35334 33012 35386
rect 33036 35334 33066 35386
rect 33066 35334 33078 35386
rect 33078 35334 33092 35386
rect 33116 35334 33130 35386
rect 33130 35334 33142 35386
rect 33142 35334 33172 35386
rect 33196 35334 33206 35386
rect 33206 35334 33252 35386
rect 32956 35332 33012 35334
rect 33036 35332 33092 35334
rect 33116 35332 33172 35334
rect 33196 35332 33252 35334
rect 32956 34298 33012 34300
rect 33036 34298 33092 34300
rect 33116 34298 33172 34300
rect 33196 34298 33252 34300
rect 32956 34246 33002 34298
rect 33002 34246 33012 34298
rect 33036 34246 33066 34298
rect 33066 34246 33078 34298
rect 33078 34246 33092 34298
rect 33116 34246 33130 34298
rect 33130 34246 33142 34298
rect 33142 34246 33172 34298
rect 33196 34246 33206 34298
rect 33206 34246 33252 34298
rect 32956 34244 33012 34246
rect 33036 34244 33092 34246
rect 33116 34244 33172 34246
rect 33196 34244 33252 34246
rect 32956 33210 33012 33212
rect 33036 33210 33092 33212
rect 33116 33210 33172 33212
rect 33196 33210 33252 33212
rect 32956 33158 33002 33210
rect 33002 33158 33012 33210
rect 33036 33158 33066 33210
rect 33066 33158 33078 33210
rect 33078 33158 33092 33210
rect 33116 33158 33130 33210
rect 33130 33158 33142 33210
rect 33142 33158 33172 33210
rect 33196 33158 33206 33210
rect 33206 33158 33252 33210
rect 32956 33156 33012 33158
rect 33036 33156 33092 33158
rect 33116 33156 33172 33158
rect 33196 33156 33252 33158
rect 32770 32952 32826 33008
rect 32956 32122 33012 32124
rect 33036 32122 33092 32124
rect 33116 32122 33172 32124
rect 33196 32122 33252 32124
rect 32956 32070 33002 32122
rect 33002 32070 33012 32122
rect 33036 32070 33066 32122
rect 33066 32070 33078 32122
rect 33078 32070 33092 32122
rect 33116 32070 33130 32122
rect 33130 32070 33142 32122
rect 33142 32070 33172 32122
rect 33196 32070 33206 32122
rect 33206 32070 33252 32122
rect 32956 32068 33012 32070
rect 33036 32068 33092 32070
rect 33116 32068 33172 32070
rect 33196 32068 33252 32070
rect 32586 27376 32642 27432
rect 31942 21936 31998 21992
rect 32956 31034 33012 31036
rect 33036 31034 33092 31036
rect 33116 31034 33172 31036
rect 33196 31034 33252 31036
rect 32956 30982 33002 31034
rect 33002 30982 33012 31034
rect 33036 30982 33066 31034
rect 33066 30982 33078 31034
rect 33078 30982 33092 31034
rect 33116 30982 33130 31034
rect 33130 30982 33142 31034
rect 33142 30982 33172 31034
rect 33196 30982 33206 31034
rect 33206 30982 33252 31034
rect 32956 30980 33012 30982
rect 33036 30980 33092 30982
rect 33116 30980 33172 30982
rect 33196 30980 33252 30982
rect 32956 29946 33012 29948
rect 33036 29946 33092 29948
rect 33116 29946 33172 29948
rect 33196 29946 33252 29948
rect 32956 29894 33002 29946
rect 33002 29894 33012 29946
rect 33036 29894 33066 29946
rect 33066 29894 33078 29946
rect 33078 29894 33092 29946
rect 33116 29894 33130 29946
rect 33130 29894 33142 29946
rect 33142 29894 33172 29946
rect 33196 29894 33206 29946
rect 33206 29894 33252 29946
rect 32956 29892 33012 29894
rect 33036 29892 33092 29894
rect 33116 29892 33172 29894
rect 33196 29892 33252 29894
rect 32956 28858 33012 28860
rect 33036 28858 33092 28860
rect 33116 28858 33172 28860
rect 33196 28858 33252 28860
rect 32956 28806 33002 28858
rect 33002 28806 33012 28858
rect 33036 28806 33066 28858
rect 33066 28806 33078 28858
rect 33078 28806 33092 28858
rect 33116 28806 33130 28858
rect 33130 28806 33142 28858
rect 33142 28806 33172 28858
rect 33196 28806 33206 28858
rect 33206 28806 33252 28858
rect 32956 28804 33012 28806
rect 33036 28804 33092 28806
rect 33116 28804 33172 28806
rect 33196 28804 33252 28806
rect 33414 34892 33416 34912
rect 33416 34892 33468 34912
rect 33468 34892 33470 34912
rect 33414 34856 33470 34892
rect 35254 44684 35256 44704
rect 35256 44684 35308 44704
rect 35308 44684 35310 44704
rect 35254 44648 35310 44684
rect 32126 21936 32182 21992
rect 32678 25200 32734 25256
rect 32956 27770 33012 27772
rect 33036 27770 33092 27772
rect 33116 27770 33172 27772
rect 33196 27770 33252 27772
rect 32956 27718 33002 27770
rect 33002 27718 33012 27770
rect 33036 27718 33066 27770
rect 33066 27718 33078 27770
rect 33078 27718 33092 27770
rect 33116 27718 33130 27770
rect 33130 27718 33142 27770
rect 33142 27718 33172 27770
rect 33196 27718 33206 27770
rect 33206 27718 33252 27770
rect 32956 27716 33012 27718
rect 33036 27716 33092 27718
rect 33116 27716 33172 27718
rect 33196 27716 33252 27718
rect 33230 26968 33286 27024
rect 32956 26682 33012 26684
rect 33036 26682 33092 26684
rect 33116 26682 33172 26684
rect 33196 26682 33252 26684
rect 32956 26630 33002 26682
rect 33002 26630 33012 26682
rect 33036 26630 33066 26682
rect 33066 26630 33078 26682
rect 33078 26630 33092 26682
rect 33116 26630 33130 26682
rect 33130 26630 33142 26682
rect 33142 26630 33172 26682
rect 33196 26630 33206 26682
rect 33206 26630 33252 26682
rect 32956 26628 33012 26630
rect 33036 26628 33092 26630
rect 33116 26628 33172 26630
rect 33196 26628 33252 26630
rect 32956 25594 33012 25596
rect 33036 25594 33092 25596
rect 33116 25594 33172 25596
rect 33196 25594 33252 25596
rect 32956 25542 33002 25594
rect 33002 25542 33012 25594
rect 33036 25542 33066 25594
rect 33066 25542 33078 25594
rect 33078 25542 33092 25594
rect 33116 25542 33130 25594
rect 33130 25542 33142 25594
rect 33142 25542 33172 25594
rect 33196 25542 33206 25594
rect 33206 25542 33252 25594
rect 32956 25540 33012 25542
rect 33036 25540 33092 25542
rect 33116 25540 33172 25542
rect 33196 25540 33252 25542
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 33874 30368 33930 30424
rect 34058 31320 34114 31376
rect 34150 30252 34206 30288
rect 34150 30232 34152 30252
rect 34152 30232 34204 30252
rect 34204 30232 34206 30252
rect 33690 26968 33746 27024
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 34794 31456 34850 31512
rect 34978 30504 35034 30560
rect 35898 39516 35900 39536
rect 35900 39516 35952 39536
rect 35952 39516 35954 39536
rect 35898 39480 35954 39516
rect 36542 44240 36598 44296
rect 37646 44240 37702 44296
rect 37956 54426 38012 54428
rect 38036 54426 38092 54428
rect 38116 54426 38172 54428
rect 38196 54426 38252 54428
rect 37956 54374 38002 54426
rect 38002 54374 38012 54426
rect 38036 54374 38066 54426
rect 38066 54374 38078 54426
rect 38078 54374 38092 54426
rect 38116 54374 38130 54426
rect 38130 54374 38142 54426
rect 38142 54374 38172 54426
rect 38196 54374 38206 54426
rect 38206 54374 38252 54426
rect 37956 54372 38012 54374
rect 38036 54372 38092 54374
rect 38116 54372 38172 54374
rect 38196 54372 38252 54374
rect 37956 53338 38012 53340
rect 38036 53338 38092 53340
rect 38116 53338 38172 53340
rect 38196 53338 38252 53340
rect 37956 53286 38002 53338
rect 38002 53286 38012 53338
rect 38036 53286 38066 53338
rect 38066 53286 38078 53338
rect 38078 53286 38092 53338
rect 38116 53286 38130 53338
rect 38130 53286 38142 53338
rect 38142 53286 38172 53338
rect 38196 53286 38206 53338
rect 38206 53286 38252 53338
rect 37956 53284 38012 53286
rect 38036 53284 38092 53286
rect 38116 53284 38172 53286
rect 38196 53284 38252 53286
rect 37956 52250 38012 52252
rect 38036 52250 38092 52252
rect 38116 52250 38172 52252
rect 38196 52250 38252 52252
rect 37956 52198 38002 52250
rect 38002 52198 38012 52250
rect 38036 52198 38066 52250
rect 38066 52198 38078 52250
rect 38078 52198 38092 52250
rect 38116 52198 38130 52250
rect 38130 52198 38142 52250
rect 38142 52198 38172 52250
rect 38196 52198 38206 52250
rect 38206 52198 38252 52250
rect 37956 52196 38012 52198
rect 38036 52196 38092 52198
rect 38116 52196 38172 52198
rect 38196 52196 38252 52198
rect 37956 51162 38012 51164
rect 38036 51162 38092 51164
rect 38116 51162 38172 51164
rect 38196 51162 38252 51164
rect 37956 51110 38002 51162
rect 38002 51110 38012 51162
rect 38036 51110 38066 51162
rect 38066 51110 38078 51162
rect 38078 51110 38092 51162
rect 38116 51110 38130 51162
rect 38130 51110 38142 51162
rect 38142 51110 38172 51162
rect 38196 51110 38206 51162
rect 38206 51110 38252 51162
rect 37956 51108 38012 51110
rect 38036 51108 38092 51110
rect 38116 51108 38172 51110
rect 38196 51108 38252 51110
rect 37956 50074 38012 50076
rect 38036 50074 38092 50076
rect 38116 50074 38172 50076
rect 38196 50074 38252 50076
rect 37956 50022 38002 50074
rect 38002 50022 38012 50074
rect 38036 50022 38066 50074
rect 38066 50022 38078 50074
rect 38078 50022 38092 50074
rect 38116 50022 38130 50074
rect 38130 50022 38142 50074
rect 38142 50022 38172 50074
rect 38196 50022 38206 50074
rect 38206 50022 38252 50074
rect 37956 50020 38012 50022
rect 38036 50020 38092 50022
rect 38116 50020 38172 50022
rect 38196 50020 38252 50022
rect 37956 48986 38012 48988
rect 38036 48986 38092 48988
rect 38116 48986 38172 48988
rect 38196 48986 38252 48988
rect 37956 48934 38002 48986
rect 38002 48934 38012 48986
rect 38036 48934 38066 48986
rect 38066 48934 38078 48986
rect 38078 48934 38092 48986
rect 38116 48934 38130 48986
rect 38130 48934 38142 48986
rect 38142 48934 38172 48986
rect 38196 48934 38206 48986
rect 38206 48934 38252 48986
rect 37956 48932 38012 48934
rect 38036 48932 38092 48934
rect 38116 48932 38172 48934
rect 38196 48932 38252 48934
rect 37956 47898 38012 47900
rect 38036 47898 38092 47900
rect 38116 47898 38172 47900
rect 38196 47898 38252 47900
rect 37956 47846 38002 47898
rect 38002 47846 38012 47898
rect 38036 47846 38066 47898
rect 38066 47846 38078 47898
rect 38078 47846 38092 47898
rect 38116 47846 38130 47898
rect 38130 47846 38142 47898
rect 38142 47846 38172 47898
rect 38196 47846 38206 47898
rect 38206 47846 38252 47898
rect 37956 47844 38012 47846
rect 38036 47844 38092 47846
rect 38116 47844 38172 47846
rect 38196 47844 38252 47846
rect 37956 46810 38012 46812
rect 38036 46810 38092 46812
rect 38116 46810 38172 46812
rect 38196 46810 38252 46812
rect 37956 46758 38002 46810
rect 38002 46758 38012 46810
rect 38036 46758 38066 46810
rect 38066 46758 38078 46810
rect 38078 46758 38092 46810
rect 38116 46758 38130 46810
rect 38130 46758 38142 46810
rect 38142 46758 38172 46810
rect 38196 46758 38206 46810
rect 38206 46758 38252 46810
rect 37956 46756 38012 46758
rect 38036 46756 38092 46758
rect 38116 46756 38172 46758
rect 38196 46756 38252 46758
rect 37956 45722 38012 45724
rect 38036 45722 38092 45724
rect 38116 45722 38172 45724
rect 38196 45722 38252 45724
rect 37956 45670 38002 45722
rect 38002 45670 38012 45722
rect 38036 45670 38066 45722
rect 38066 45670 38078 45722
rect 38078 45670 38092 45722
rect 38116 45670 38130 45722
rect 38130 45670 38142 45722
rect 38142 45670 38172 45722
rect 38196 45670 38206 45722
rect 38206 45670 38252 45722
rect 37956 45668 38012 45670
rect 38036 45668 38092 45670
rect 38116 45668 38172 45670
rect 38196 45668 38252 45670
rect 37956 44634 38012 44636
rect 38036 44634 38092 44636
rect 38116 44634 38172 44636
rect 38196 44634 38252 44636
rect 37956 44582 38002 44634
rect 38002 44582 38012 44634
rect 38036 44582 38066 44634
rect 38066 44582 38078 44634
rect 38078 44582 38092 44634
rect 38116 44582 38130 44634
rect 38130 44582 38142 44634
rect 38142 44582 38172 44634
rect 38196 44582 38206 44634
rect 38206 44582 38252 44634
rect 37956 44580 38012 44582
rect 38036 44580 38092 44582
rect 38116 44580 38172 44582
rect 38196 44580 38252 44582
rect 37186 43424 37242 43480
rect 36082 32000 36138 32056
rect 35990 31864 36046 31920
rect 35990 31184 36046 31240
rect 35898 30912 35954 30968
rect 34518 24112 34574 24168
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 34886 24248 34942 24304
rect 35254 27512 35310 27568
rect 37094 39480 37150 39536
rect 37956 43546 38012 43548
rect 38036 43546 38092 43548
rect 38116 43546 38172 43548
rect 38196 43546 38252 43548
rect 37956 43494 38002 43546
rect 38002 43494 38012 43546
rect 38036 43494 38066 43546
rect 38066 43494 38078 43546
rect 38078 43494 38092 43546
rect 38116 43494 38130 43546
rect 38130 43494 38142 43546
rect 38142 43494 38172 43546
rect 38196 43494 38206 43546
rect 38206 43494 38252 43546
rect 37956 43492 38012 43494
rect 38036 43492 38092 43494
rect 38116 43492 38172 43494
rect 38196 43492 38252 43494
rect 37956 42458 38012 42460
rect 38036 42458 38092 42460
rect 38116 42458 38172 42460
rect 38196 42458 38252 42460
rect 37956 42406 38002 42458
rect 38002 42406 38012 42458
rect 38036 42406 38066 42458
rect 38066 42406 38078 42458
rect 38078 42406 38092 42458
rect 38116 42406 38130 42458
rect 38130 42406 38142 42458
rect 38142 42406 38172 42458
rect 38196 42406 38206 42458
rect 38206 42406 38252 42458
rect 37956 42404 38012 42406
rect 38036 42404 38092 42406
rect 38116 42404 38172 42406
rect 38196 42404 38252 42406
rect 37956 41370 38012 41372
rect 38036 41370 38092 41372
rect 38116 41370 38172 41372
rect 38196 41370 38252 41372
rect 37956 41318 38002 41370
rect 38002 41318 38012 41370
rect 38036 41318 38066 41370
rect 38066 41318 38078 41370
rect 38078 41318 38092 41370
rect 38116 41318 38130 41370
rect 38130 41318 38142 41370
rect 38142 41318 38172 41370
rect 38196 41318 38206 41370
rect 38206 41318 38252 41370
rect 37956 41316 38012 41318
rect 38036 41316 38092 41318
rect 38116 41316 38172 41318
rect 38196 41316 38252 41318
rect 37002 33380 37058 33416
rect 37002 33360 37004 33380
rect 37004 33360 37056 33380
rect 37056 33360 37058 33380
rect 36910 33224 36966 33280
rect 36634 32000 36690 32056
rect 36726 30368 36782 30424
rect 36818 28464 36874 28520
rect 37956 40282 38012 40284
rect 38036 40282 38092 40284
rect 38116 40282 38172 40284
rect 38196 40282 38252 40284
rect 37956 40230 38002 40282
rect 38002 40230 38012 40282
rect 38036 40230 38066 40282
rect 38066 40230 38078 40282
rect 38078 40230 38092 40282
rect 38116 40230 38130 40282
rect 38130 40230 38142 40282
rect 38142 40230 38172 40282
rect 38196 40230 38206 40282
rect 38206 40230 38252 40282
rect 37956 40228 38012 40230
rect 38036 40228 38092 40230
rect 38116 40228 38172 40230
rect 38196 40228 38252 40230
rect 37956 39194 38012 39196
rect 38036 39194 38092 39196
rect 38116 39194 38172 39196
rect 38196 39194 38252 39196
rect 37956 39142 38002 39194
rect 38002 39142 38012 39194
rect 38036 39142 38066 39194
rect 38066 39142 38078 39194
rect 38078 39142 38092 39194
rect 38116 39142 38130 39194
rect 38130 39142 38142 39194
rect 38142 39142 38172 39194
rect 38196 39142 38206 39194
rect 38206 39142 38252 39194
rect 37956 39140 38012 39142
rect 38036 39140 38092 39142
rect 38116 39140 38172 39142
rect 38196 39140 38252 39142
rect 37956 38106 38012 38108
rect 38036 38106 38092 38108
rect 38116 38106 38172 38108
rect 38196 38106 38252 38108
rect 37956 38054 38002 38106
rect 38002 38054 38012 38106
rect 38036 38054 38066 38106
rect 38066 38054 38078 38106
rect 38078 38054 38092 38106
rect 38116 38054 38130 38106
rect 38130 38054 38142 38106
rect 38142 38054 38172 38106
rect 38196 38054 38206 38106
rect 38206 38054 38252 38106
rect 37956 38052 38012 38054
rect 38036 38052 38092 38054
rect 38116 38052 38172 38054
rect 38196 38052 38252 38054
rect 38106 37168 38162 37224
rect 37956 37018 38012 37020
rect 38036 37018 38092 37020
rect 38116 37018 38172 37020
rect 38196 37018 38252 37020
rect 37956 36966 38002 37018
rect 38002 36966 38012 37018
rect 38036 36966 38066 37018
rect 38066 36966 38078 37018
rect 38078 36966 38092 37018
rect 38116 36966 38130 37018
rect 38130 36966 38142 37018
rect 38142 36966 38172 37018
rect 38196 36966 38206 37018
rect 38206 36966 38252 37018
rect 37956 36964 38012 36966
rect 38036 36964 38092 36966
rect 38116 36964 38172 36966
rect 38196 36964 38252 36966
rect 37956 35930 38012 35932
rect 38036 35930 38092 35932
rect 38116 35930 38172 35932
rect 38196 35930 38252 35932
rect 37956 35878 38002 35930
rect 38002 35878 38012 35930
rect 38036 35878 38066 35930
rect 38066 35878 38078 35930
rect 38078 35878 38092 35930
rect 38116 35878 38130 35930
rect 38130 35878 38142 35930
rect 38142 35878 38172 35930
rect 38196 35878 38206 35930
rect 38206 35878 38252 35930
rect 37956 35876 38012 35878
rect 38036 35876 38092 35878
rect 38116 35876 38172 35878
rect 38196 35876 38252 35878
rect 38382 36216 38438 36272
rect 38382 35672 38438 35728
rect 37956 34842 38012 34844
rect 38036 34842 38092 34844
rect 38116 34842 38172 34844
rect 38196 34842 38252 34844
rect 37956 34790 38002 34842
rect 38002 34790 38012 34842
rect 38036 34790 38066 34842
rect 38066 34790 38078 34842
rect 38078 34790 38092 34842
rect 38116 34790 38130 34842
rect 38130 34790 38142 34842
rect 38142 34790 38172 34842
rect 38196 34790 38206 34842
rect 38206 34790 38252 34842
rect 37956 34788 38012 34790
rect 38036 34788 38092 34790
rect 38116 34788 38172 34790
rect 38196 34788 38252 34790
rect 37462 33224 37518 33280
rect 37278 30504 37334 30560
rect 37956 33754 38012 33756
rect 38036 33754 38092 33756
rect 38116 33754 38172 33756
rect 38196 33754 38252 33756
rect 37956 33702 38002 33754
rect 38002 33702 38012 33754
rect 38036 33702 38066 33754
rect 38066 33702 38078 33754
rect 38078 33702 38092 33754
rect 38116 33702 38130 33754
rect 38130 33702 38142 33754
rect 38142 33702 38172 33754
rect 38196 33702 38206 33754
rect 38206 33702 38252 33754
rect 37956 33700 38012 33702
rect 38036 33700 38092 33702
rect 38116 33700 38172 33702
rect 38196 33700 38252 33702
rect 37830 33516 37886 33552
rect 37830 33496 37832 33516
rect 37832 33496 37884 33516
rect 37884 33496 37886 33516
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 37956 32666 38012 32668
rect 38036 32666 38092 32668
rect 38116 32666 38172 32668
rect 38196 32666 38252 32668
rect 37956 32614 38002 32666
rect 38002 32614 38012 32666
rect 38036 32614 38066 32666
rect 38066 32614 38078 32666
rect 38078 32614 38092 32666
rect 38116 32614 38130 32666
rect 38130 32614 38142 32666
rect 38142 32614 38172 32666
rect 38196 32614 38206 32666
rect 38206 32614 38252 32666
rect 37956 32612 38012 32614
rect 38036 32612 38092 32614
rect 38116 32612 38172 32614
rect 38196 32612 38252 32614
rect 37738 31456 37794 31512
rect 37554 31320 37610 31376
rect 37370 27104 37426 27160
rect 37462 26968 37518 27024
rect 38290 32408 38346 32464
rect 37956 31578 38012 31580
rect 38036 31578 38092 31580
rect 38116 31578 38172 31580
rect 38196 31578 38252 31580
rect 37956 31526 38002 31578
rect 38002 31526 38012 31578
rect 38036 31526 38066 31578
rect 38066 31526 38078 31578
rect 38078 31526 38092 31578
rect 38116 31526 38130 31578
rect 38130 31526 38142 31578
rect 38142 31526 38172 31578
rect 38196 31526 38206 31578
rect 38206 31526 38252 31578
rect 37956 31524 38012 31526
rect 38036 31524 38092 31526
rect 38116 31524 38172 31526
rect 38196 31524 38252 31526
rect 38198 31356 38200 31376
rect 38200 31356 38252 31376
rect 38252 31356 38254 31376
rect 38198 31320 38254 31356
rect 37956 30490 38012 30492
rect 38036 30490 38092 30492
rect 38116 30490 38172 30492
rect 38196 30490 38252 30492
rect 37956 30438 38002 30490
rect 38002 30438 38012 30490
rect 38036 30438 38066 30490
rect 38066 30438 38078 30490
rect 38078 30438 38092 30490
rect 38116 30438 38130 30490
rect 38130 30438 38142 30490
rect 38142 30438 38172 30490
rect 38196 30438 38206 30490
rect 38206 30438 38252 30490
rect 37956 30436 38012 30438
rect 38036 30436 38092 30438
rect 38116 30436 38172 30438
rect 38196 30436 38252 30438
rect 37956 29402 38012 29404
rect 38036 29402 38092 29404
rect 38116 29402 38172 29404
rect 38196 29402 38252 29404
rect 37956 29350 38002 29402
rect 38002 29350 38012 29402
rect 38036 29350 38066 29402
rect 38066 29350 38078 29402
rect 38078 29350 38092 29402
rect 38116 29350 38130 29402
rect 38130 29350 38142 29402
rect 38142 29350 38172 29402
rect 38196 29350 38206 29402
rect 38206 29350 38252 29402
rect 37956 29348 38012 29350
rect 38036 29348 38092 29350
rect 38116 29348 38172 29350
rect 38196 29348 38252 29350
rect 37956 28314 38012 28316
rect 38036 28314 38092 28316
rect 38116 28314 38172 28316
rect 38196 28314 38252 28316
rect 37956 28262 38002 28314
rect 38002 28262 38012 28314
rect 38036 28262 38066 28314
rect 38066 28262 38078 28314
rect 38078 28262 38092 28314
rect 38116 28262 38130 28314
rect 38130 28262 38142 28314
rect 38142 28262 38172 28314
rect 38196 28262 38206 28314
rect 38206 28262 38252 28314
rect 37956 28260 38012 28262
rect 38036 28260 38092 28262
rect 38116 28260 38172 28262
rect 38196 28260 38252 28262
rect 39118 37204 39120 37224
rect 39120 37204 39172 37224
rect 39172 37204 39174 37224
rect 39118 37168 39174 37204
rect 38658 31748 38714 31784
rect 38658 31728 38660 31748
rect 38660 31728 38712 31748
rect 38712 31728 38714 31748
rect 37956 27226 38012 27228
rect 38036 27226 38092 27228
rect 38116 27226 38172 27228
rect 38196 27226 38252 27228
rect 37956 27174 38002 27226
rect 38002 27174 38012 27226
rect 38036 27174 38066 27226
rect 38066 27174 38078 27226
rect 38078 27174 38092 27226
rect 38116 27174 38130 27226
rect 38130 27174 38142 27226
rect 38142 27174 38172 27226
rect 38196 27174 38206 27226
rect 38206 27174 38252 27226
rect 37956 27172 38012 27174
rect 38036 27172 38092 27174
rect 38116 27172 38172 27174
rect 38196 27172 38252 27174
rect 37956 26138 38012 26140
rect 38036 26138 38092 26140
rect 38116 26138 38172 26140
rect 38196 26138 38252 26140
rect 37956 26086 38002 26138
rect 38002 26086 38012 26138
rect 38036 26086 38066 26138
rect 38066 26086 38078 26138
rect 38078 26086 38092 26138
rect 38116 26086 38130 26138
rect 38130 26086 38142 26138
rect 38142 26086 38172 26138
rect 38196 26086 38206 26138
rect 38206 26086 38252 26138
rect 37956 26084 38012 26086
rect 38036 26084 38092 26086
rect 38116 26084 38172 26086
rect 38196 26084 38252 26086
rect 37956 25050 38012 25052
rect 38036 25050 38092 25052
rect 38116 25050 38172 25052
rect 38196 25050 38252 25052
rect 37956 24998 38002 25050
rect 38002 24998 38012 25050
rect 38036 24998 38066 25050
rect 38066 24998 38078 25050
rect 38078 24998 38092 25050
rect 38116 24998 38130 25050
rect 38130 24998 38142 25050
rect 38142 24998 38172 25050
rect 38196 24998 38206 25050
rect 38206 24998 38252 25050
rect 37956 24996 38012 24998
rect 38036 24996 38092 24998
rect 38116 24996 38172 24998
rect 38196 24996 38252 24998
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 39026 31340 39082 31376
rect 39026 31320 39028 31340
rect 39028 31320 39080 31340
rect 39080 31320 39082 31340
rect 39394 36080 39450 36136
rect 39302 35536 39358 35592
rect 40406 41656 40462 41712
rect 42956 53882 43012 53884
rect 43036 53882 43092 53884
rect 43116 53882 43172 53884
rect 43196 53882 43252 53884
rect 42956 53830 43002 53882
rect 43002 53830 43012 53882
rect 43036 53830 43066 53882
rect 43066 53830 43078 53882
rect 43078 53830 43092 53882
rect 43116 53830 43130 53882
rect 43130 53830 43142 53882
rect 43142 53830 43172 53882
rect 43196 53830 43206 53882
rect 43206 53830 43252 53882
rect 42956 53828 43012 53830
rect 43036 53828 43092 53830
rect 43116 53828 43172 53830
rect 43196 53828 43252 53830
rect 42956 52794 43012 52796
rect 43036 52794 43092 52796
rect 43116 52794 43172 52796
rect 43196 52794 43252 52796
rect 42956 52742 43002 52794
rect 43002 52742 43012 52794
rect 43036 52742 43066 52794
rect 43066 52742 43078 52794
rect 43078 52742 43092 52794
rect 43116 52742 43130 52794
rect 43130 52742 43142 52794
rect 43142 52742 43172 52794
rect 43196 52742 43206 52794
rect 43206 52742 43252 52794
rect 42956 52740 43012 52742
rect 43036 52740 43092 52742
rect 43116 52740 43172 52742
rect 43196 52740 43252 52742
rect 42956 51706 43012 51708
rect 43036 51706 43092 51708
rect 43116 51706 43172 51708
rect 43196 51706 43252 51708
rect 42956 51654 43002 51706
rect 43002 51654 43012 51706
rect 43036 51654 43066 51706
rect 43066 51654 43078 51706
rect 43078 51654 43092 51706
rect 43116 51654 43130 51706
rect 43130 51654 43142 51706
rect 43142 51654 43172 51706
rect 43196 51654 43206 51706
rect 43206 51654 43252 51706
rect 42956 51652 43012 51654
rect 43036 51652 43092 51654
rect 43116 51652 43172 51654
rect 43196 51652 43252 51654
rect 42956 50618 43012 50620
rect 43036 50618 43092 50620
rect 43116 50618 43172 50620
rect 43196 50618 43252 50620
rect 42956 50566 43002 50618
rect 43002 50566 43012 50618
rect 43036 50566 43066 50618
rect 43066 50566 43078 50618
rect 43078 50566 43092 50618
rect 43116 50566 43130 50618
rect 43130 50566 43142 50618
rect 43142 50566 43172 50618
rect 43196 50566 43206 50618
rect 43206 50566 43252 50618
rect 42956 50564 43012 50566
rect 43036 50564 43092 50566
rect 43116 50564 43172 50566
rect 43196 50564 43252 50566
rect 42956 49530 43012 49532
rect 43036 49530 43092 49532
rect 43116 49530 43172 49532
rect 43196 49530 43252 49532
rect 42956 49478 43002 49530
rect 43002 49478 43012 49530
rect 43036 49478 43066 49530
rect 43066 49478 43078 49530
rect 43078 49478 43092 49530
rect 43116 49478 43130 49530
rect 43130 49478 43142 49530
rect 43142 49478 43172 49530
rect 43196 49478 43206 49530
rect 43206 49478 43252 49530
rect 42956 49476 43012 49478
rect 43036 49476 43092 49478
rect 43116 49476 43172 49478
rect 43196 49476 43252 49478
rect 42956 48442 43012 48444
rect 43036 48442 43092 48444
rect 43116 48442 43172 48444
rect 43196 48442 43252 48444
rect 42956 48390 43002 48442
rect 43002 48390 43012 48442
rect 43036 48390 43066 48442
rect 43066 48390 43078 48442
rect 43078 48390 43092 48442
rect 43116 48390 43130 48442
rect 43130 48390 43142 48442
rect 43142 48390 43172 48442
rect 43196 48390 43206 48442
rect 43206 48390 43252 48442
rect 42956 48388 43012 48390
rect 43036 48388 43092 48390
rect 43116 48388 43172 48390
rect 43196 48388 43252 48390
rect 42956 47354 43012 47356
rect 43036 47354 43092 47356
rect 43116 47354 43172 47356
rect 43196 47354 43252 47356
rect 42956 47302 43002 47354
rect 43002 47302 43012 47354
rect 43036 47302 43066 47354
rect 43066 47302 43078 47354
rect 43078 47302 43092 47354
rect 43116 47302 43130 47354
rect 43130 47302 43142 47354
rect 43142 47302 43172 47354
rect 43196 47302 43206 47354
rect 43206 47302 43252 47354
rect 42956 47300 43012 47302
rect 43036 47300 43092 47302
rect 43116 47300 43172 47302
rect 43196 47300 43252 47302
rect 42956 46266 43012 46268
rect 43036 46266 43092 46268
rect 43116 46266 43172 46268
rect 43196 46266 43252 46268
rect 42956 46214 43002 46266
rect 43002 46214 43012 46266
rect 43036 46214 43066 46266
rect 43066 46214 43078 46266
rect 43078 46214 43092 46266
rect 43116 46214 43130 46266
rect 43130 46214 43142 46266
rect 43142 46214 43172 46266
rect 43196 46214 43206 46266
rect 43206 46214 43252 46266
rect 42956 46212 43012 46214
rect 43036 46212 43092 46214
rect 43116 46212 43172 46214
rect 43196 46212 43252 46214
rect 42956 45178 43012 45180
rect 43036 45178 43092 45180
rect 43116 45178 43172 45180
rect 43196 45178 43252 45180
rect 42956 45126 43002 45178
rect 43002 45126 43012 45178
rect 43036 45126 43066 45178
rect 43066 45126 43078 45178
rect 43078 45126 43092 45178
rect 43116 45126 43130 45178
rect 43130 45126 43142 45178
rect 43142 45126 43172 45178
rect 43196 45126 43206 45178
rect 43206 45126 43252 45178
rect 42956 45124 43012 45126
rect 43036 45124 43092 45126
rect 43116 45124 43172 45126
rect 43196 45124 43252 45126
rect 42956 44090 43012 44092
rect 43036 44090 43092 44092
rect 43116 44090 43172 44092
rect 43196 44090 43252 44092
rect 42956 44038 43002 44090
rect 43002 44038 43012 44090
rect 43036 44038 43066 44090
rect 43066 44038 43078 44090
rect 43078 44038 43092 44090
rect 43116 44038 43130 44090
rect 43130 44038 43142 44090
rect 43142 44038 43172 44090
rect 43196 44038 43206 44090
rect 43206 44038 43252 44090
rect 42956 44036 43012 44038
rect 43036 44036 43092 44038
rect 43116 44036 43172 44038
rect 43196 44036 43252 44038
rect 39302 30640 39358 30696
rect 40866 34992 40922 35048
rect 41326 42064 41382 42120
rect 42956 43002 43012 43004
rect 43036 43002 43092 43004
rect 43116 43002 43172 43004
rect 43196 43002 43252 43004
rect 42956 42950 43002 43002
rect 43002 42950 43012 43002
rect 43036 42950 43066 43002
rect 43066 42950 43078 43002
rect 43078 42950 43092 43002
rect 43116 42950 43130 43002
rect 43130 42950 43142 43002
rect 43142 42950 43172 43002
rect 43196 42950 43206 43002
rect 43206 42950 43252 43002
rect 42956 42948 43012 42950
rect 43036 42948 43092 42950
rect 43116 42948 43172 42950
rect 43196 42948 43252 42950
rect 40590 31900 40592 31920
rect 40592 31900 40644 31920
rect 40644 31900 40646 31920
rect 40590 31864 40646 31900
rect 40590 27124 40646 27160
rect 40590 27104 40592 27124
rect 40592 27104 40644 27124
rect 40644 27104 40646 27124
rect 42956 41914 43012 41916
rect 43036 41914 43092 41916
rect 43116 41914 43172 41916
rect 43196 41914 43252 41916
rect 42956 41862 43002 41914
rect 43002 41862 43012 41914
rect 43036 41862 43066 41914
rect 43066 41862 43078 41914
rect 43078 41862 43092 41914
rect 43116 41862 43130 41914
rect 43130 41862 43142 41914
rect 43142 41862 43172 41914
rect 43196 41862 43206 41914
rect 43206 41862 43252 41914
rect 42956 41860 43012 41862
rect 43036 41860 43092 41862
rect 43116 41860 43172 41862
rect 43196 41860 43252 41862
rect 42956 40826 43012 40828
rect 43036 40826 43092 40828
rect 43116 40826 43172 40828
rect 43196 40826 43252 40828
rect 42956 40774 43002 40826
rect 43002 40774 43012 40826
rect 43036 40774 43066 40826
rect 43066 40774 43078 40826
rect 43078 40774 43092 40826
rect 43116 40774 43130 40826
rect 43130 40774 43142 40826
rect 43142 40774 43172 40826
rect 43196 40774 43206 40826
rect 43206 40774 43252 40826
rect 42956 40772 43012 40774
rect 43036 40772 43092 40774
rect 43116 40772 43172 40774
rect 43196 40772 43252 40774
rect 42956 39738 43012 39740
rect 43036 39738 43092 39740
rect 43116 39738 43172 39740
rect 43196 39738 43252 39740
rect 42956 39686 43002 39738
rect 43002 39686 43012 39738
rect 43036 39686 43066 39738
rect 43066 39686 43078 39738
rect 43078 39686 43092 39738
rect 43116 39686 43130 39738
rect 43130 39686 43142 39738
rect 43142 39686 43172 39738
rect 43196 39686 43206 39738
rect 43206 39686 43252 39738
rect 42956 39684 43012 39686
rect 43036 39684 43092 39686
rect 43116 39684 43172 39686
rect 43196 39684 43252 39686
rect 42956 38650 43012 38652
rect 43036 38650 43092 38652
rect 43116 38650 43172 38652
rect 43196 38650 43252 38652
rect 42956 38598 43002 38650
rect 43002 38598 43012 38650
rect 43036 38598 43066 38650
rect 43066 38598 43078 38650
rect 43078 38598 43092 38650
rect 43116 38598 43130 38650
rect 43130 38598 43142 38650
rect 43142 38598 43172 38650
rect 43196 38598 43206 38650
rect 43206 38598 43252 38650
rect 42956 38596 43012 38598
rect 43036 38596 43092 38598
rect 43116 38596 43172 38598
rect 43196 38596 43252 38598
rect 42956 37562 43012 37564
rect 43036 37562 43092 37564
rect 43116 37562 43172 37564
rect 43196 37562 43252 37564
rect 42956 37510 43002 37562
rect 43002 37510 43012 37562
rect 43036 37510 43066 37562
rect 43066 37510 43078 37562
rect 43078 37510 43092 37562
rect 43116 37510 43130 37562
rect 43130 37510 43142 37562
rect 43142 37510 43172 37562
rect 43196 37510 43206 37562
rect 43206 37510 43252 37562
rect 42956 37508 43012 37510
rect 43036 37508 43092 37510
rect 43116 37508 43172 37510
rect 43196 37508 43252 37510
rect 42956 36474 43012 36476
rect 43036 36474 43092 36476
rect 43116 36474 43172 36476
rect 43196 36474 43252 36476
rect 42956 36422 43002 36474
rect 43002 36422 43012 36474
rect 43036 36422 43066 36474
rect 43066 36422 43078 36474
rect 43078 36422 43092 36474
rect 43116 36422 43130 36474
rect 43130 36422 43142 36474
rect 43142 36422 43172 36474
rect 43196 36422 43206 36474
rect 43206 36422 43252 36474
rect 42956 36420 43012 36422
rect 43036 36420 43092 36422
rect 43116 36420 43172 36422
rect 43196 36420 43252 36422
rect 42956 35386 43012 35388
rect 43036 35386 43092 35388
rect 43116 35386 43172 35388
rect 43196 35386 43252 35388
rect 42956 35334 43002 35386
rect 43002 35334 43012 35386
rect 43036 35334 43066 35386
rect 43066 35334 43078 35386
rect 43078 35334 43092 35386
rect 43116 35334 43130 35386
rect 43130 35334 43142 35386
rect 43142 35334 43172 35386
rect 43196 35334 43206 35386
rect 43206 35334 43252 35386
rect 42956 35332 43012 35334
rect 43036 35332 43092 35334
rect 43116 35332 43172 35334
rect 43196 35332 43252 35334
rect 42956 34298 43012 34300
rect 43036 34298 43092 34300
rect 43116 34298 43172 34300
rect 43196 34298 43252 34300
rect 42956 34246 43002 34298
rect 43002 34246 43012 34298
rect 43036 34246 43066 34298
rect 43066 34246 43078 34298
rect 43078 34246 43092 34298
rect 43116 34246 43130 34298
rect 43130 34246 43142 34298
rect 43142 34246 43172 34298
rect 43196 34246 43206 34298
rect 43206 34246 43252 34298
rect 42956 34244 43012 34246
rect 43036 34244 43092 34246
rect 43116 34244 43172 34246
rect 43196 34244 43252 34246
rect 42956 33210 43012 33212
rect 43036 33210 43092 33212
rect 43116 33210 43172 33212
rect 43196 33210 43252 33212
rect 42956 33158 43002 33210
rect 43002 33158 43012 33210
rect 43036 33158 43066 33210
rect 43066 33158 43078 33210
rect 43078 33158 43092 33210
rect 43116 33158 43130 33210
rect 43130 33158 43142 33210
rect 43142 33158 43172 33210
rect 43196 33158 43206 33210
rect 43206 33158 43252 33210
rect 42956 33156 43012 33158
rect 43036 33156 43092 33158
rect 43116 33156 43172 33158
rect 43196 33156 43252 33158
rect 42956 32122 43012 32124
rect 43036 32122 43092 32124
rect 43116 32122 43172 32124
rect 43196 32122 43252 32124
rect 42956 32070 43002 32122
rect 43002 32070 43012 32122
rect 43036 32070 43066 32122
rect 43066 32070 43078 32122
rect 43078 32070 43092 32122
rect 43116 32070 43130 32122
rect 43130 32070 43142 32122
rect 43142 32070 43172 32122
rect 43196 32070 43206 32122
rect 43206 32070 43252 32122
rect 42956 32068 43012 32070
rect 43036 32068 43092 32070
rect 43116 32068 43172 32070
rect 43196 32068 43252 32070
rect 47956 54426 48012 54428
rect 48036 54426 48092 54428
rect 48116 54426 48172 54428
rect 48196 54426 48252 54428
rect 47956 54374 48002 54426
rect 48002 54374 48012 54426
rect 48036 54374 48066 54426
rect 48066 54374 48078 54426
rect 48078 54374 48092 54426
rect 48116 54374 48130 54426
rect 48130 54374 48142 54426
rect 48142 54374 48172 54426
rect 48196 54374 48206 54426
rect 48206 54374 48252 54426
rect 47956 54372 48012 54374
rect 48036 54372 48092 54374
rect 48116 54372 48172 54374
rect 48196 54372 48252 54374
rect 43994 31728 44050 31784
rect 42956 31034 43012 31036
rect 43036 31034 43092 31036
rect 43116 31034 43172 31036
rect 43196 31034 43252 31036
rect 42956 30982 43002 31034
rect 43002 30982 43012 31034
rect 43036 30982 43066 31034
rect 43066 30982 43078 31034
rect 43078 30982 43092 31034
rect 43116 30982 43130 31034
rect 43130 30982 43142 31034
rect 43142 30982 43172 31034
rect 43196 30982 43206 31034
rect 43206 30982 43252 31034
rect 42956 30980 43012 30982
rect 43036 30980 43092 30982
rect 43116 30980 43172 30982
rect 43196 30980 43252 30982
rect 42956 29946 43012 29948
rect 43036 29946 43092 29948
rect 43116 29946 43172 29948
rect 43196 29946 43252 29948
rect 42956 29894 43002 29946
rect 43002 29894 43012 29946
rect 43036 29894 43066 29946
rect 43066 29894 43078 29946
rect 43078 29894 43092 29946
rect 43116 29894 43130 29946
rect 43130 29894 43142 29946
rect 43142 29894 43172 29946
rect 43196 29894 43206 29946
rect 43206 29894 43252 29946
rect 42956 29892 43012 29894
rect 43036 29892 43092 29894
rect 43116 29892 43172 29894
rect 43196 29892 43252 29894
rect 42956 28858 43012 28860
rect 43036 28858 43092 28860
rect 43116 28858 43172 28860
rect 43196 28858 43252 28860
rect 42956 28806 43002 28858
rect 43002 28806 43012 28858
rect 43036 28806 43066 28858
rect 43066 28806 43078 28858
rect 43078 28806 43092 28858
rect 43116 28806 43130 28858
rect 43130 28806 43142 28858
rect 43142 28806 43172 28858
rect 43196 28806 43206 28858
rect 43206 28806 43252 28858
rect 42956 28804 43012 28806
rect 43036 28804 43092 28806
rect 43116 28804 43172 28806
rect 43196 28804 43252 28806
rect 42956 27770 43012 27772
rect 43036 27770 43092 27772
rect 43116 27770 43172 27772
rect 43196 27770 43252 27772
rect 42956 27718 43002 27770
rect 43002 27718 43012 27770
rect 43036 27718 43066 27770
rect 43066 27718 43078 27770
rect 43078 27718 43092 27770
rect 43116 27718 43130 27770
rect 43130 27718 43142 27770
rect 43142 27718 43172 27770
rect 43196 27718 43206 27770
rect 43206 27718 43252 27770
rect 42956 27716 43012 27718
rect 43036 27716 43092 27718
rect 43116 27716 43172 27718
rect 43196 27716 43252 27718
rect 42154 27124 42210 27160
rect 42154 27104 42156 27124
rect 42156 27104 42208 27124
rect 42208 27104 42210 27124
rect 42956 26682 43012 26684
rect 43036 26682 43092 26684
rect 43116 26682 43172 26684
rect 43196 26682 43252 26684
rect 42956 26630 43002 26682
rect 43002 26630 43012 26682
rect 43036 26630 43066 26682
rect 43066 26630 43078 26682
rect 43078 26630 43092 26682
rect 43116 26630 43130 26682
rect 43130 26630 43142 26682
rect 43142 26630 43172 26682
rect 43196 26630 43206 26682
rect 43206 26630 43252 26682
rect 42956 26628 43012 26630
rect 43036 26628 43092 26630
rect 43116 26628 43172 26630
rect 43196 26628 43252 26630
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 42956 25594 43012 25596
rect 43036 25594 43092 25596
rect 43116 25594 43172 25596
rect 43196 25594 43252 25596
rect 42956 25542 43002 25594
rect 43002 25542 43012 25594
rect 43036 25542 43066 25594
rect 43066 25542 43078 25594
rect 43078 25542 43092 25594
rect 43116 25542 43130 25594
rect 43130 25542 43142 25594
rect 43142 25542 43172 25594
rect 43196 25542 43206 25594
rect 43206 25542 43252 25594
rect 42956 25540 43012 25542
rect 43036 25540 43092 25542
rect 43116 25540 43172 25542
rect 43196 25540 43252 25542
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 53338 48012 53340
rect 48036 53338 48092 53340
rect 48116 53338 48172 53340
rect 48196 53338 48252 53340
rect 47956 53286 48002 53338
rect 48002 53286 48012 53338
rect 48036 53286 48066 53338
rect 48066 53286 48078 53338
rect 48078 53286 48092 53338
rect 48116 53286 48130 53338
rect 48130 53286 48142 53338
rect 48142 53286 48172 53338
rect 48196 53286 48206 53338
rect 48206 53286 48252 53338
rect 47956 53284 48012 53286
rect 48036 53284 48092 53286
rect 48116 53284 48172 53286
rect 48196 53284 48252 53286
rect 47956 52250 48012 52252
rect 48036 52250 48092 52252
rect 48116 52250 48172 52252
rect 48196 52250 48252 52252
rect 47956 52198 48002 52250
rect 48002 52198 48012 52250
rect 48036 52198 48066 52250
rect 48066 52198 48078 52250
rect 48078 52198 48092 52250
rect 48116 52198 48130 52250
rect 48130 52198 48142 52250
rect 48142 52198 48172 52250
rect 48196 52198 48206 52250
rect 48206 52198 48252 52250
rect 47956 52196 48012 52198
rect 48036 52196 48092 52198
rect 48116 52196 48172 52198
rect 48196 52196 48252 52198
rect 49054 51856 49110 51912
rect 49054 51176 49110 51232
rect 47956 51162 48012 51164
rect 48036 51162 48092 51164
rect 48116 51162 48172 51164
rect 48196 51162 48252 51164
rect 47956 51110 48002 51162
rect 48002 51110 48012 51162
rect 48036 51110 48066 51162
rect 48066 51110 48078 51162
rect 48078 51110 48092 51162
rect 48116 51110 48130 51162
rect 48130 51110 48142 51162
rect 48142 51110 48172 51162
rect 48196 51110 48206 51162
rect 48206 51110 48252 51162
rect 47956 51108 48012 51110
rect 48036 51108 48092 51110
rect 48116 51108 48172 51110
rect 48196 51108 48252 51110
rect 48962 50496 49018 50552
rect 47956 50074 48012 50076
rect 48036 50074 48092 50076
rect 48116 50074 48172 50076
rect 48196 50074 48252 50076
rect 47956 50022 48002 50074
rect 48002 50022 48012 50074
rect 48036 50022 48066 50074
rect 48066 50022 48078 50074
rect 48078 50022 48092 50074
rect 48116 50022 48130 50074
rect 48130 50022 48142 50074
rect 48142 50022 48172 50074
rect 48196 50022 48206 50074
rect 48206 50022 48252 50074
rect 47956 50020 48012 50022
rect 48036 50020 48092 50022
rect 48116 50020 48172 50022
rect 48196 50020 48252 50022
rect 47956 48986 48012 48988
rect 48036 48986 48092 48988
rect 48116 48986 48172 48988
rect 48196 48986 48252 48988
rect 47956 48934 48002 48986
rect 48002 48934 48012 48986
rect 48036 48934 48066 48986
rect 48066 48934 48078 48986
rect 48078 48934 48092 48986
rect 48116 48934 48130 48986
rect 48130 48934 48142 48986
rect 48142 48934 48172 48986
rect 48196 48934 48206 48986
rect 48206 48934 48252 48986
rect 47956 48932 48012 48934
rect 48036 48932 48092 48934
rect 48116 48932 48172 48934
rect 48196 48932 48252 48934
rect 47956 47898 48012 47900
rect 48036 47898 48092 47900
rect 48116 47898 48172 47900
rect 48196 47898 48252 47900
rect 47956 47846 48002 47898
rect 48002 47846 48012 47898
rect 48036 47846 48066 47898
rect 48066 47846 48078 47898
rect 48078 47846 48092 47898
rect 48116 47846 48130 47898
rect 48130 47846 48142 47898
rect 48142 47846 48172 47898
rect 48196 47846 48206 47898
rect 48206 47846 48252 47898
rect 47956 47844 48012 47846
rect 48036 47844 48092 47846
rect 48116 47844 48172 47846
rect 48196 47844 48252 47846
rect 47956 46810 48012 46812
rect 48036 46810 48092 46812
rect 48116 46810 48172 46812
rect 48196 46810 48252 46812
rect 47956 46758 48002 46810
rect 48002 46758 48012 46810
rect 48036 46758 48066 46810
rect 48066 46758 48078 46810
rect 48078 46758 48092 46810
rect 48116 46758 48130 46810
rect 48130 46758 48142 46810
rect 48142 46758 48172 46810
rect 48196 46758 48206 46810
rect 48206 46758 48252 46810
rect 47956 46756 48012 46758
rect 48036 46756 48092 46758
rect 48116 46756 48172 46758
rect 48196 46756 48252 46758
rect 47956 45722 48012 45724
rect 48036 45722 48092 45724
rect 48116 45722 48172 45724
rect 48196 45722 48252 45724
rect 47956 45670 48002 45722
rect 48002 45670 48012 45722
rect 48036 45670 48066 45722
rect 48066 45670 48078 45722
rect 48078 45670 48092 45722
rect 48116 45670 48130 45722
rect 48130 45670 48142 45722
rect 48142 45670 48172 45722
rect 48196 45670 48206 45722
rect 48206 45670 48252 45722
rect 47956 45668 48012 45670
rect 48036 45668 48092 45670
rect 48116 45668 48172 45670
rect 48196 45668 48252 45670
rect 48318 45056 48374 45112
rect 47956 44634 48012 44636
rect 48036 44634 48092 44636
rect 48116 44634 48172 44636
rect 48196 44634 48252 44636
rect 47956 44582 48002 44634
rect 48002 44582 48012 44634
rect 48036 44582 48066 44634
rect 48066 44582 48078 44634
rect 48078 44582 48092 44634
rect 48116 44582 48130 44634
rect 48130 44582 48142 44634
rect 48142 44582 48172 44634
rect 48196 44582 48206 44634
rect 48206 44582 48252 44634
rect 47956 44580 48012 44582
rect 48036 44580 48092 44582
rect 48116 44580 48172 44582
rect 48196 44580 48252 44582
rect 47956 43546 48012 43548
rect 48036 43546 48092 43548
rect 48116 43546 48172 43548
rect 48196 43546 48252 43548
rect 47956 43494 48002 43546
rect 48002 43494 48012 43546
rect 48036 43494 48066 43546
rect 48066 43494 48078 43546
rect 48078 43494 48092 43546
rect 48116 43494 48130 43546
rect 48130 43494 48142 43546
rect 48142 43494 48172 43546
rect 48196 43494 48206 43546
rect 48206 43494 48252 43546
rect 47956 43492 48012 43494
rect 48036 43492 48092 43494
rect 48116 43492 48172 43494
rect 48196 43492 48252 43494
rect 47956 42458 48012 42460
rect 48036 42458 48092 42460
rect 48116 42458 48172 42460
rect 48196 42458 48252 42460
rect 47956 42406 48002 42458
rect 48002 42406 48012 42458
rect 48036 42406 48066 42458
rect 48066 42406 48078 42458
rect 48078 42406 48092 42458
rect 48116 42406 48130 42458
rect 48130 42406 48142 42458
rect 48142 42406 48172 42458
rect 48196 42406 48206 42458
rect 48206 42406 48252 42458
rect 47956 42404 48012 42406
rect 48036 42404 48092 42406
rect 48116 42404 48172 42406
rect 48196 42404 48252 42406
rect 47956 41370 48012 41372
rect 48036 41370 48092 41372
rect 48116 41370 48172 41372
rect 48196 41370 48252 41372
rect 47956 41318 48002 41370
rect 48002 41318 48012 41370
rect 48036 41318 48066 41370
rect 48066 41318 48078 41370
rect 48078 41318 48092 41370
rect 48116 41318 48130 41370
rect 48130 41318 48142 41370
rect 48142 41318 48172 41370
rect 48196 41318 48206 41370
rect 48206 41318 48252 41370
rect 47956 41316 48012 41318
rect 48036 41316 48092 41318
rect 48116 41316 48172 41318
rect 48196 41316 48252 41318
rect 49054 49816 49110 49872
rect 49054 49172 49056 49192
rect 49056 49172 49108 49192
rect 49108 49172 49110 49192
rect 49054 49136 49110 49172
rect 48502 44376 48558 44432
rect 48502 43732 48504 43752
rect 48504 43732 48556 43752
rect 48556 43732 48558 43752
rect 48502 43696 48558 43732
rect 48502 43016 48558 43072
rect 48502 42336 48558 42392
rect 48502 41656 48558 41712
rect 48502 41012 48504 41032
rect 48504 41012 48556 41032
rect 48556 41012 48558 41032
rect 48502 40976 48558 41012
rect 47956 40282 48012 40284
rect 48036 40282 48092 40284
rect 48116 40282 48172 40284
rect 48196 40282 48252 40284
rect 47956 40230 48002 40282
rect 48002 40230 48012 40282
rect 48036 40230 48066 40282
rect 48066 40230 48078 40282
rect 48078 40230 48092 40282
rect 48116 40230 48130 40282
rect 48130 40230 48142 40282
rect 48142 40230 48172 40282
rect 48196 40230 48206 40282
rect 48206 40230 48252 40282
rect 47956 40228 48012 40230
rect 48036 40228 48092 40230
rect 48116 40228 48172 40230
rect 48196 40228 48252 40230
rect 47956 39194 48012 39196
rect 48036 39194 48092 39196
rect 48116 39194 48172 39196
rect 48196 39194 48252 39196
rect 47956 39142 48002 39194
rect 48002 39142 48012 39194
rect 48036 39142 48066 39194
rect 48066 39142 48078 39194
rect 48078 39142 48092 39194
rect 48116 39142 48130 39194
rect 48130 39142 48142 39194
rect 48142 39142 48172 39194
rect 48196 39142 48206 39194
rect 48206 39142 48252 39194
rect 47956 39140 48012 39142
rect 48036 39140 48092 39142
rect 48116 39140 48172 39142
rect 48196 39140 48252 39142
rect 47956 38106 48012 38108
rect 48036 38106 48092 38108
rect 48116 38106 48172 38108
rect 48196 38106 48252 38108
rect 47956 38054 48002 38106
rect 48002 38054 48012 38106
rect 48036 38054 48066 38106
rect 48066 38054 48078 38106
rect 48078 38054 48092 38106
rect 48116 38054 48130 38106
rect 48130 38054 48142 38106
rect 48142 38054 48172 38106
rect 48196 38054 48206 38106
rect 48206 38054 48252 38106
rect 47956 38052 48012 38054
rect 48036 38052 48092 38054
rect 48116 38052 48172 38054
rect 48196 38052 48252 38054
rect 47956 37018 48012 37020
rect 48036 37018 48092 37020
rect 48116 37018 48172 37020
rect 48196 37018 48252 37020
rect 47956 36966 48002 37018
rect 48002 36966 48012 37018
rect 48036 36966 48066 37018
rect 48066 36966 48078 37018
rect 48078 36966 48092 37018
rect 48116 36966 48130 37018
rect 48130 36966 48142 37018
rect 48142 36966 48172 37018
rect 48196 36966 48206 37018
rect 48206 36966 48252 37018
rect 47956 36964 48012 36966
rect 48036 36964 48092 36966
rect 48116 36964 48172 36966
rect 48196 36964 48252 36966
rect 47956 35930 48012 35932
rect 48036 35930 48092 35932
rect 48116 35930 48172 35932
rect 48196 35930 48252 35932
rect 47956 35878 48002 35930
rect 48002 35878 48012 35930
rect 48036 35878 48066 35930
rect 48066 35878 48078 35930
rect 48078 35878 48092 35930
rect 48116 35878 48130 35930
rect 48130 35878 48142 35930
rect 48142 35878 48172 35930
rect 48196 35878 48206 35930
rect 48206 35878 48252 35930
rect 47956 35876 48012 35878
rect 48036 35876 48092 35878
rect 48116 35876 48172 35878
rect 48196 35876 48252 35878
rect 48502 40296 48558 40352
rect 48502 39616 48558 39672
rect 48502 38936 48558 38992
rect 48502 36896 48558 36952
rect 48778 39500 48834 39536
rect 48778 39480 48780 39500
rect 48780 39480 48832 39500
rect 48832 39480 48834 39500
rect 49054 48456 49110 48512
rect 49054 47776 49110 47832
rect 49054 47096 49110 47152
rect 49146 45736 49202 45792
rect 48594 35536 48650 35592
rect 47956 34842 48012 34844
rect 48036 34842 48092 34844
rect 48116 34842 48172 34844
rect 48196 34842 48252 34844
rect 47956 34790 48002 34842
rect 48002 34790 48012 34842
rect 48036 34790 48066 34842
rect 48066 34790 48078 34842
rect 48078 34790 48092 34842
rect 48116 34790 48130 34842
rect 48130 34790 48142 34842
rect 48142 34790 48172 34842
rect 48196 34790 48206 34842
rect 48206 34790 48252 34842
rect 47956 34788 48012 34790
rect 48036 34788 48092 34790
rect 48116 34788 48172 34790
rect 48196 34788 48252 34790
rect 49330 38292 49332 38312
rect 49332 38292 49384 38312
rect 49384 38292 49386 38312
rect 49330 38256 49386 38292
rect 49330 37576 49386 37632
rect 49422 37168 49478 37224
rect 49330 36216 49386 36272
rect 49330 35536 49386 35592
rect 49330 34856 49386 34912
rect 49330 34176 49386 34232
rect 47956 33754 48012 33756
rect 48036 33754 48092 33756
rect 48116 33754 48172 33756
rect 48196 33754 48252 33756
rect 47956 33702 48002 33754
rect 48002 33702 48012 33754
rect 48036 33702 48066 33754
rect 48066 33702 48078 33754
rect 48078 33702 48092 33754
rect 48116 33702 48130 33754
rect 48130 33702 48142 33754
rect 48142 33702 48172 33754
rect 48196 33702 48206 33754
rect 48206 33702 48252 33754
rect 47956 33700 48012 33702
rect 48036 33700 48092 33702
rect 48116 33700 48172 33702
rect 48196 33700 48252 33702
rect 49330 33496 49386 33552
rect 47956 32666 48012 32668
rect 48036 32666 48092 32668
rect 48116 32666 48172 32668
rect 48196 32666 48252 32668
rect 47956 32614 48002 32666
rect 48002 32614 48012 32666
rect 48036 32614 48066 32666
rect 48066 32614 48078 32666
rect 48078 32614 48092 32666
rect 48116 32614 48130 32666
rect 48130 32614 48142 32666
rect 48142 32614 48172 32666
rect 48196 32614 48206 32666
rect 48206 32614 48252 32666
rect 47956 32612 48012 32614
rect 48036 32612 48092 32614
rect 48116 32612 48172 32614
rect 48196 32612 48252 32614
rect 49330 32852 49332 32872
rect 49332 32852 49384 32872
rect 49384 32852 49386 32872
rect 49330 32816 49386 32852
rect 48502 32136 48558 32192
rect 47956 31578 48012 31580
rect 48036 31578 48092 31580
rect 48116 31578 48172 31580
rect 48196 31578 48252 31580
rect 47956 31526 48002 31578
rect 48002 31526 48012 31578
rect 48036 31526 48066 31578
rect 48066 31526 48078 31578
rect 48078 31526 48092 31578
rect 48116 31526 48130 31578
rect 48130 31526 48142 31578
rect 48142 31526 48172 31578
rect 48196 31526 48206 31578
rect 48206 31526 48252 31578
rect 47956 31524 48012 31526
rect 48036 31524 48092 31526
rect 48116 31524 48172 31526
rect 48196 31524 48252 31526
rect 48502 31456 48558 31512
rect 48502 30776 48558 30832
rect 47956 30490 48012 30492
rect 48036 30490 48092 30492
rect 48116 30490 48172 30492
rect 48196 30490 48252 30492
rect 47956 30438 48002 30490
rect 48002 30438 48012 30490
rect 48036 30438 48066 30490
rect 48066 30438 48078 30490
rect 48078 30438 48092 30490
rect 48116 30438 48130 30490
rect 48130 30438 48142 30490
rect 48142 30438 48172 30490
rect 48196 30438 48206 30490
rect 48206 30438 48252 30490
rect 47956 30436 48012 30438
rect 48036 30436 48092 30438
rect 48116 30436 48172 30438
rect 48196 30436 48252 30438
rect 48502 29416 48558 29472
rect 47956 29402 48012 29404
rect 48036 29402 48092 29404
rect 48116 29402 48172 29404
rect 48196 29402 48252 29404
rect 47956 29350 48002 29402
rect 48002 29350 48012 29402
rect 48036 29350 48066 29402
rect 48066 29350 48078 29402
rect 48078 29350 48092 29402
rect 48116 29350 48130 29402
rect 48130 29350 48142 29402
rect 48142 29350 48172 29402
rect 48196 29350 48206 29402
rect 48206 29350 48252 29402
rect 47956 29348 48012 29350
rect 48036 29348 48092 29350
rect 48116 29348 48172 29350
rect 48196 29348 48252 29350
rect 47956 28314 48012 28316
rect 48036 28314 48092 28316
rect 48116 28314 48172 28316
rect 48196 28314 48252 28316
rect 47956 28262 48002 28314
rect 48002 28262 48012 28314
rect 48036 28262 48066 28314
rect 48066 28262 48078 28314
rect 48078 28262 48092 28314
rect 48116 28262 48130 28314
rect 48130 28262 48142 28314
rect 48142 28262 48172 28314
rect 48196 28262 48206 28314
rect 48206 28262 48252 28314
rect 47956 28260 48012 28262
rect 48036 28260 48092 28262
rect 48116 28260 48172 28262
rect 48196 28260 48252 28262
rect 48502 27412 48504 27432
rect 48504 27412 48556 27432
rect 48556 27412 48558 27432
rect 48502 27376 48558 27412
rect 47956 27226 48012 27228
rect 48036 27226 48092 27228
rect 48116 27226 48172 27228
rect 48196 27226 48252 27228
rect 47956 27174 48002 27226
rect 48002 27174 48012 27226
rect 48036 27174 48066 27226
rect 48066 27174 48078 27226
rect 48078 27174 48092 27226
rect 48116 27174 48130 27226
rect 48130 27174 48142 27226
rect 48142 27174 48172 27226
rect 48196 27174 48206 27226
rect 48206 27174 48252 27226
rect 47956 27172 48012 27174
rect 48036 27172 48092 27174
rect 48116 27172 48172 27174
rect 48196 27172 48252 27174
rect 48502 26696 48558 26752
rect 47956 26138 48012 26140
rect 48036 26138 48092 26140
rect 48116 26138 48172 26140
rect 48196 26138 48252 26140
rect 47956 26086 48002 26138
rect 48002 26086 48012 26138
rect 48036 26086 48066 26138
rect 48066 26086 48078 26138
rect 48078 26086 48092 26138
rect 48116 26086 48130 26138
rect 48130 26086 48142 26138
rect 48142 26086 48172 26138
rect 48196 26086 48206 26138
rect 48206 26086 48252 26138
rect 47956 26084 48012 26086
rect 48036 26084 48092 26086
rect 48116 26084 48172 26086
rect 48196 26084 48252 26086
rect 48410 26016 48466 26072
rect 47956 25050 48012 25052
rect 48036 25050 48092 25052
rect 48116 25050 48172 25052
rect 48196 25050 48252 25052
rect 47956 24998 48002 25050
rect 48002 24998 48012 25050
rect 48036 24998 48066 25050
rect 48066 24998 48078 25050
rect 48078 24998 48092 25050
rect 48116 24998 48130 25050
rect 48130 24998 48142 25050
rect 48142 24998 48172 25050
rect 48196 24998 48206 25050
rect 48206 24998 48252 25050
rect 47956 24996 48012 24998
rect 48036 24996 48092 24998
rect 48116 24996 48172 24998
rect 48196 24996 48252 24998
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 49330 30096 49386 30152
rect 49330 28736 49386 28792
rect 49330 28056 49386 28112
rect 49330 25336 49386 25392
rect 49146 24692 49148 24712
rect 49148 24692 49200 24712
rect 49200 24692 49202 24712
rect 49146 24656 49202 24692
rect 49146 23976 49202 24032
rect 49146 23296 49202 23352
rect 49146 22616 49202 22672
rect 49146 21972 49148 21992
rect 49148 21972 49200 21992
rect 49200 21972 49202 21992
rect 49146 21936 49202 21972
rect 49146 21256 49202 21312
rect 49146 20576 49202 20632
rect 49146 19896 49202 19952
rect 49146 19216 49202 19272
rect 49146 18536 49202 18592
rect 49146 17856 49202 17912
rect 49146 17176 49202 17232
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 49146 16516 49202 16552
rect 49146 16496 49148 16516
rect 49148 16496 49200 16516
rect 49200 16496 49202 16516
rect 49146 15816 49202 15872
rect 49146 15136 49202 15192
rect 49146 14456 49202 14512
rect 49146 13812 49148 13832
rect 49148 13812 49200 13832
rect 49200 13812 49202 13832
rect 49146 13776 49202 13812
rect 49146 13096 49202 13152
rect 49146 12416 49202 12472
rect 49146 11736 49202 11792
rect 49146 11092 49148 11112
rect 49148 11092 49200 11112
rect 49200 11092 49202 11112
rect 49146 11056 49202 11092
rect 49146 10376 49202 10432
rect 49146 9696 49202 9752
rect 49146 9016 49202 9072
rect 49146 8372 49148 8392
rect 49148 8372 49200 8392
rect 49200 8372 49202 8392
rect 49146 8336 49202 8372
rect 49146 7656 49202 7712
rect 49146 6976 49202 7032
rect 49146 6296 49202 6352
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 5652 49148 5672
rect 49148 5652 49200 5672
rect 49200 5652 49202 5672
rect 49146 5616 49202 5652
rect 49330 4972 49332 4992
rect 49332 4972 49384 4992
rect 49384 4972 49386 4992
rect 49330 4936 49386 4972
rect 49146 4256 49202 4312
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 55042 800 55072
rect 2773 55042 2839 55045
rect 0 55040 2839 55042
rect 0 54984 2778 55040
rect 2834 54984 2839 55040
rect 0 54982 2839 54984
rect 0 54952 800 54982
rect 2773 54979 2839 54982
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 27946 54432 28262 54433
rect 27946 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28262 54432
rect 27946 54367 28262 54368
rect 37946 54432 38262 54433
rect 37946 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38262 54432
rect 37946 54367 38262 54368
rect 47946 54432 48262 54433
rect 47946 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48262 54432
rect 47946 54367 48262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 32946 53888 33262 53889
rect 32946 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33262 53888
rect 32946 53823 33262 53824
rect 42946 53888 43262 53889
rect 42946 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43262 53888
rect 42946 53823 43262 53824
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 27946 53344 28262 53345
rect 27946 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28262 53344
rect 27946 53279 28262 53280
rect 37946 53344 38262 53345
rect 37946 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38262 53344
rect 37946 53279 38262 53280
rect 47946 53344 48262 53345
rect 47946 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48262 53344
rect 47946 53279 48262 53280
rect 2946 52800 3262 52801
rect 0 52730 800 52760
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 32946 52800 33262 52801
rect 32946 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33262 52800
rect 32946 52735 33262 52736
rect 42946 52800 43262 52801
rect 42946 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43262 52800
rect 42946 52735 43262 52736
rect 933 52730 999 52733
rect 0 52728 999 52730
rect 0 52672 938 52728
rect 994 52672 999 52728
rect 0 52670 999 52672
rect 0 52640 800 52670
rect 933 52667 999 52670
rect 50200 52504 51000 52624
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 27946 52256 28262 52257
rect 27946 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28262 52256
rect 27946 52191 28262 52192
rect 37946 52256 38262 52257
rect 37946 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38262 52256
rect 37946 52191 38262 52192
rect 47946 52256 48262 52257
rect 47946 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48262 52256
rect 47946 52191 48262 52192
rect 49049 51914 49115 51917
rect 50200 51914 51000 51944
rect 49049 51912 51000 51914
rect 49049 51856 49054 51912
rect 49110 51856 51000 51912
rect 49049 51854 51000 51856
rect 49049 51851 49115 51854
rect 50200 51824 51000 51854
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 32946 51712 33262 51713
rect 32946 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33262 51712
rect 32946 51647 33262 51648
rect 42946 51712 43262 51713
rect 42946 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43262 51712
rect 42946 51647 43262 51648
rect 49049 51234 49115 51237
rect 50200 51234 51000 51264
rect 49049 51232 51000 51234
rect 49049 51176 49054 51232
rect 49110 51176 51000 51232
rect 49049 51174 51000 51176
rect 49049 51171 49115 51174
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 27946 51168 28262 51169
rect 27946 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28262 51168
rect 27946 51103 28262 51104
rect 37946 51168 38262 51169
rect 37946 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38262 51168
rect 37946 51103 38262 51104
rect 47946 51168 48262 51169
rect 47946 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48262 51168
rect 50200 51144 51000 51174
rect 47946 51103 48262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 32946 50624 33262 50625
rect 32946 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33262 50624
rect 32946 50559 33262 50560
rect 42946 50624 43262 50625
rect 42946 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43262 50624
rect 42946 50559 43262 50560
rect 48957 50554 49023 50557
rect 50200 50554 51000 50584
rect 48957 50552 51000 50554
rect 48957 50496 48962 50552
rect 49018 50496 51000 50552
rect 48957 50494 51000 50496
rect 48957 50491 49023 50494
rect 50200 50464 51000 50494
rect 0 50418 800 50448
rect 933 50418 999 50421
rect 0 50416 999 50418
rect 0 50360 938 50416
rect 994 50360 999 50416
rect 0 50358 999 50360
rect 0 50328 800 50358
rect 933 50355 999 50358
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 27946 50080 28262 50081
rect 27946 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28262 50080
rect 27946 50015 28262 50016
rect 37946 50080 38262 50081
rect 37946 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38262 50080
rect 37946 50015 38262 50016
rect 47946 50080 48262 50081
rect 47946 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48262 50080
rect 47946 50015 48262 50016
rect 49049 49874 49115 49877
rect 50200 49874 51000 49904
rect 49049 49872 51000 49874
rect 49049 49816 49054 49872
rect 49110 49816 51000 49872
rect 49049 49814 51000 49816
rect 49049 49811 49115 49814
rect 50200 49784 51000 49814
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 32946 49536 33262 49537
rect 32946 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33262 49536
rect 32946 49471 33262 49472
rect 42946 49536 43262 49537
rect 42946 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43262 49536
rect 42946 49471 43262 49472
rect 49049 49194 49115 49197
rect 50200 49194 51000 49224
rect 49049 49192 51000 49194
rect 49049 49136 49054 49192
rect 49110 49136 51000 49192
rect 49049 49134 51000 49136
rect 49049 49131 49115 49134
rect 50200 49104 51000 49134
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 27946 48992 28262 48993
rect 27946 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28262 48992
rect 27946 48927 28262 48928
rect 37946 48992 38262 48993
rect 37946 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38262 48992
rect 37946 48927 38262 48928
rect 47946 48992 48262 48993
rect 47946 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48262 48992
rect 47946 48927 48262 48928
rect 49049 48514 49115 48517
rect 50200 48514 51000 48544
rect 49049 48512 51000 48514
rect 49049 48456 49054 48512
rect 49110 48456 51000 48512
rect 49049 48454 51000 48456
rect 49049 48451 49115 48454
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 32946 48448 33262 48449
rect 32946 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33262 48448
rect 32946 48383 33262 48384
rect 42946 48448 43262 48449
rect 42946 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43262 48448
rect 50200 48424 51000 48454
rect 42946 48383 43262 48384
rect 0 48106 800 48136
rect 933 48106 999 48109
rect 0 48104 999 48106
rect 0 48048 938 48104
rect 994 48048 999 48104
rect 0 48046 999 48048
rect 0 48016 800 48046
rect 933 48043 999 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 27946 47904 28262 47905
rect 27946 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28262 47904
rect 27946 47839 28262 47840
rect 37946 47904 38262 47905
rect 37946 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38262 47904
rect 37946 47839 38262 47840
rect 47946 47904 48262 47905
rect 47946 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48262 47904
rect 47946 47839 48262 47840
rect 49049 47834 49115 47837
rect 50200 47834 51000 47864
rect 49049 47832 51000 47834
rect 49049 47776 49054 47832
rect 49110 47776 51000 47832
rect 49049 47774 51000 47776
rect 49049 47771 49115 47774
rect 50200 47744 51000 47774
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 32946 47360 33262 47361
rect 32946 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33262 47360
rect 32946 47295 33262 47296
rect 42946 47360 43262 47361
rect 42946 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43262 47360
rect 42946 47295 43262 47296
rect 49049 47154 49115 47157
rect 50200 47154 51000 47184
rect 49049 47152 51000 47154
rect 49049 47096 49054 47152
rect 49110 47096 51000 47152
rect 49049 47094 51000 47096
rect 49049 47091 49115 47094
rect 50200 47064 51000 47094
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 27946 46816 28262 46817
rect 27946 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28262 46816
rect 27946 46751 28262 46752
rect 37946 46816 38262 46817
rect 37946 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38262 46816
rect 37946 46751 38262 46752
rect 47946 46816 48262 46817
rect 47946 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48262 46816
rect 47946 46751 48262 46752
rect 50200 46384 51000 46504
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 32946 46272 33262 46273
rect 32946 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33262 46272
rect 32946 46207 33262 46208
rect 42946 46272 43262 46273
rect 42946 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43262 46272
rect 42946 46207 43262 46208
rect 0 45794 800 45824
rect 933 45794 999 45797
rect 0 45792 999 45794
rect 0 45736 938 45792
rect 994 45736 999 45792
rect 0 45734 999 45736
rect 0 45704 800 45734
rect 933 45731 999 45734
rect 49141 45794 49207 45797
rect 50200 45794 51000 45824
rect 49141 45792 51000 45794
rect 49141 45736 49146 45792
rect 49202 45736 51000 45792
rect 49141 45734 51000 45736
rect 49141 45731 49207 45734
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 27946 45728 28262 45729
rect 27946 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28262 45728
rect 27946 45663 28262 45664
rect 37946 45728 38262 45729
rect 37946 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38262 45728
rect 37946 45663 38262 45664
rect 47946 45728 48262 45729
rect 47946 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48262 45728
rect 50200 45704 51000 45734
rect 47946 45663 48262 45664
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 32946 45184 33262 45185
rect 32946 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33262 45184
rect 32946 45119 33262 45120
rect 42946 45184 43262 45185
rect 42946 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43262 45184
rect 42946 45119 43262 45120
rect 48313 45114 48379 45117
rect 50200 45114 51000 45144
rect 48313 45112 51000 45114
rect 48313 45056 48318 45112
rect 48374 45056 51000 45112
rect 48313 45054 51000 45056
rect 48313 45051 48379 45054
rect 50200 45024 51000 45054
rect 35249 44706 35315 44709
rect 35382 44706 35388 44708
rect 35249 44704 35388 44706
rect 35249 44648 35254 44704
rect 35310 44648 35388 44704
rect 35249 44646 35388 44648
rect 35249 44643 35315 44646
rect 35382 44644 35388 44646
rect 35452 44644 35458 44708
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 27946 44640 28262 44641
rect 27946 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28262 44640
rect 27946 44575 28262 44576
rect 37946 44640 38262 44641
rect 37946 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38262 44640
rect 37946 44575 38262 44576
rect 47946 44640 48262 44641
rect 47946 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48262 44640
rect 47946 44575 48262 44576
rect 48497 44434 48563 44437
rect 50200 44434 51000 44464
rect 48497 44432 51000 44434
rect 48497 44376 48502 44432
rect 48558 44376 51000 44432
rect 48497 44374 51000 44376
rect 48497 44371 48563 44374
rect 50200 44344 51000 44374
rect 36537 44298 36603 44301
rect 36670 44298 36676 44300
rect 36537 44296 36676 44298
rect 36537 44240 36542 44296
rect 36598 44240 36676 44296
rect 36537 44238 36676 44240
rect 36537 44235 36603 44238
rect 36670 44236 36676 44238
rect 36740 44236 36746 44300
rect 37222 44236 37228 44300
rect 37292 44298 37298 44300
rect 37641 44298 37707 44301
rect 37292 44296 37707 44298
rect 37292 44240 37646 44296
rect 37702 44240 37707 44296
rect 37292 44238 37707 44240
rect 37292 44236 37298 44238
rect 37641 44235 37707 44238
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 32946 44096 33262 44097
rect 32946 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33262 44096
rect 32946 44031 33262 44032
rect 42946 44096 43262 44097
rect 42946 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43262 44096
rect 42946 44031 43262 44032
rect 48497 43754 48563 43757
rect 50200 43754 51000 43784
rect 48497 43752 51000 43754
rect 48497 43696 48502 43752
rect 48558 43696 51000 43752
rect 48497 43694 51000 43696
rect 48497 43691 48563 43694
rect 50200 43664 51000 43694
rect 7946 43552 8262 43553
rect 0 43392 800 43512
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 27946 43552 28262 43553
rect 27946 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28262 43552
rect 27946 43487 28262 43488
rect 37946 43552 38262 43553
rect 37946 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38262 43552
rect 37946 43487 38262 43488
rect 47946 43552 48262 43553
rect 47946 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48262 43552
rect 47946 43487 48262 43488
rect 35934 43420 35940 43484
rect 36004 43482 36010 43484
rect 37181 43482 37247 43485
rect 36004 43480 37247 43482
rect 36004 43424 37186 43480
rect 37242 43424 37247 43480
rect 36004 43422 37247 43424
rect 36004 43420 36010 43422
rect 37181 43419 37247 43422
rect 48497 43074 48563 43077
rect 50200 43074 51000 43104
rect 48497 43072 51000 43074
rect 48497 43016 48502 43072
rect 48558 43016 51000 43072
rect 48497 43014 51000 43016
rect 48497 43011 48563 43014
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 32946 43008 33262 43009
rect 32946 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33262 43008
rect 32946 42943 33262 42944
rect 42946 43008 43262 43009
rect 42946 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43262 43008
rect 50200 42984 51000 43014
rect 42946 42943 43262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 27946 42464 28262 42465
rect 27946 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28262 42464
rect 27946 42399 28262 42400
rect 37946 42464 38262 42465
rect 37946 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38262 42464
rect 37946 42399 38262 42400
rect 47946 42464 48262 42465
rect 47946 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48262 42464
rect 47946 42399 48262 42400
rect 48497 42394 48563 42397
rect 50200 42394 51000 42424
rect 48497 42392 51000 42394
rect 48497 42336 48502 42392
rect 48558 42336 51000 42392
rect 48497 42334 51000 42336
rect 48497 42331 48563 42334
rect 50200 42304 51000 42334
rect 39982 42060 39988 42124
rect 40052 42122 40058 42124
rect 41321 42122 41387 42125
rect 40052 42120 41387 42122
rect 40052 42064 41326 42120
rect 41382 42064 41387 42120
rect 40052 42062 41387 42064
rect 40052 42060 40058 42062
rect 41321 42059 41387 42062
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 32946 41920 33262 41921
rect 32946 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33262 41920
rect 32946 41855 33262 41856
rect 42946 41920 43262 41921
rect 42946 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43262 41920
rect 42946 41855 43262 41856
rect 40401 41714 40467 41717
rect 40534 41714 40540 41716
rect 40401 41712 40540 41714
rect 40401 41656 40406 41712
rect 40462 41656 40540 41712
rect 40401 41654 40540 41656
rect 40401 41651 40467 41654
rect 40534 41652 40540 41654
rect 40604 41652 40610 41716
rect 48497 41714 48563 41717
rect 50200 41714 51000 41744
rect 48497 41712 51000 41714
rect 48497 41656 48502 41712
rect 48558 41656 51000 41712
rect 48497 41654 51000 41656
rect 48497 41651 48563 41654
rect 50200 41624 51000 41654
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 27946 41376 28262 41377
rect 27946 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28262 41376
rect 27946 41311 28262 41312
rect 37946 41376 38262 41377
rect 37946 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38262 41376
rect 37946 41311 38262 41312
rect 47946 41376 48262 41377
rect 47946 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48262 41376
rect 47946 41311 48262 41312
rect 0 41170 800 41200
rect 1669 41170 1735 41173
rect 0 41168 1735 41170
rect 0 41112 1674 41168
rect 1730 41112 1735 41168
rect 0 41110 1735 41112
rect 0 41080 800 41110
rect 1669 41107 1735 41110
rect 48497 41034 48563 41037
rect 50200 41034 51000 41064
rect 48497 41032 51000 41034
rect 48497 40976 48502 41032
rect 48558 40976 51000 41032
rect 48497 40974 51000 40976
rect 48497 40971 48563 40974
rect 50200 40944 51000 40974
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 32946 40832 33262 40833
rect 32946 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33262 40832
rect 32946 40767 33262 40768
rect 42946 40832 43262 40833
rect 42946 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43262 40832
rect 42946 40767 43262 40768
rect 27521 40490 27587 40493
rect 30649 40490 30715 40493
rect 27521 40488 30715 40490
rect 27521 40432 27526 40488
rect 27582 40432 30654 40488
rect 30710 40432 30715 40488
rect 27521 40430 30715 40432
rect 27521 40427 27587 40430
rect 30649 40427 30715 40430
rect 48497 40354 48563 40357
rect 50200 40354 51000 40384
rect 48497 40352 51000 40354
rect 48497 40296 48502 40352
rect 48558 40296 51000 40352
rect 48497 40294 51000 40296
rect 48497 40291 48563 40294
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 27946 40288 28262 40289
rect 27946 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28262 40288
rect 27946 40223 28262 40224
rect 37946 40288 38262 40289
rect 37946 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38262 40288
rect 37946 40223 38262 40224
rect 47946 40288 48262 40289
rect 47946 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48262 40288
rect 50200 40264 51000 40294
rect 47946 40223 48262 40224
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 32946 39744 33262 39745
rect 32946 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33262 39744
rect 32946 39679 33262 39680
rect 42946 39744 43262 39745
rect 42946 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43262 39744
rect 42946 39679 43262 39680
rect 48497 39674 48563 39677
rect 50200 39674 51000 39704
rect 48497 39672 51000 39674
rect 48497 39616 48502 39672
rect 48558 39616 51000 39672
rect 48497 39614 51000 39616
rect 48497 39611 48563 39614
rect 50200 39584 51000 39614
rect 35893 39538 35959 39541
rect 37089 39538 37155 39541
rect 48773 39538 48839 39541
rect 35893 39536 48839 39538
rect 35893 39480 35898 39536
rect 35954 39480 37094 39536
rect 37150 39480 48778 39536
rect 48834 39480 48839 39536
rect 35893 39478 48839 39480
rect 35893 39475 35959 39478
rect 37089 39475 37155 39478
rect 48773 39475 48839 39478
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 27946 39200 28262 39201
rect 27946 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28262 39200
rect 27946 39135 28262 39136
rect 37946 39200 38262 39201
rect 37946 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38262 39200
rect 37946 39135 38262 39136
rect 47946 39200 48262 39201
rect 47946 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48262 39200
rect 47946 39135 48262 39136
rect 48497 38994 48563 38997
rect 50200 38994 51000 39024
rect 48497 38992 51000 38994
rect 48497 38936 48502 38992
rect 48558 38936 51000 38992
rect 48497 38934 51000 38936
rect 48497 38931 48563 38934
rect 50200 38904 51000 38934
rect 0 38858 800 38888
rect 933 38858 999 38861
rect 0 38856 999 38858
rect 0 38800 938 38856
rect 994 38800 999 38856
rect 0 38798 999 38800
rect 0 38768 800 38798
rect 933 38795 999 38798
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 32946 38656 33262 38657
rect 32946 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33262 38656
rect 32946 38591 33262 38592
rect 42946 38656 43262 38657
rect 42946 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43262 38656
rect 42946 38591 43262 38592
rect 49325 38314 49391 38317
rect 50200 38314 51000 38344
rect 49325 38312 51000 38314
rect 49325 38256 49330 38312
rect 49386 38256 51000 38312
rect 49325 38254 51000 38256
rect 49325 38251 49391 38254
rect 50200 38224 51000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 27946 38112 28262 38113
rect 27946 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28262 38112
rect 27946 38047 28262 38048
rect 37946 38112 38262 38113
rect 37946 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38262 38112
rect 37946 38047 38262 38048
rect 47946 38112 48262 38113
rect 47946 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48262 38112
rect 47946 38047 48262 38048
rect 30833 37906 30899 37909
rect 33501 37906 33567 37909
rect 30833 37904 33567 37906
rect 30833 37848 30838 37904
rect 30894 37848 33506 37904
rect 33562 37848 33567 37904
rect 30833 37846 33567 37848
rect 30833 37843 30899 37846
rect 33501 37843 33567 37846
rect 49325 37634 49391 37637
rect 50200 37634 51000 37664
rect 49325 37632 51000 37634
rect 49325 37576 49330 37632
rect 49386 37576 51000 37632
rect 49325 37574 51000 37576
rect 49325 37571 49391 37574
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 32946 37568 33262 37569
rect 32946 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33262 37568
rect 32946 37503 33262 37504
rect 42946 37568 43262 37569
rect 42946 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43262 37568
rect 50200 37544 51000 37574
rect 42946 37503 43262 37504
rect 23289 37226 23355 37229
rect 25630 37226 25636 37228
rect 23289 37224 25636 37226
rect 23289 37168 23294 37224
rect 23350 37168 25636 37224
rect 23289 37166 25636 37168
rect 23289 37163 23355 37166
rect 25630 37164 25636 37166
rect 25700 37226 25706 37228
rect 29821 37226 29887 37229
rect 25700 37224 29887 37226
rect 25700 37168 29826 37224
rect 29882 37168 29887 37224
rect 25700 37166 29887 37168
rect 25700 37164 25706 37166
rect 29821 37163 29887 37166
rect 33685 37226 33751 37229
rect 38101 37226 38167 37229
rect 33685 37224 38167 37226
rect 33685 37168 33690 37224
rect 33746 37168 38106 37224
rect 38162 37168 38167 37224
rect 33685 37166 38167 37168
rect 33685 37163 33751 37166
rect 38101 37163 38167 37166
rect 39113 37226 39179 37229
rect 49417 37226 49483 37229
rect 39113 37224 49483 37226
rect 39113 37168 39118 37224
rect 39174 37168 49422 37224
rect 49478 37168 49483 37224
rect 39113 37166 49483 37168
rect 39113 37163 39179 37166
rect 49417 37163 49483 37166
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 27946 37024 28262 37025
rect 27946 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28262 37024
rect 27946 36959 28262 36960
rect 37946 37024 38262 37025
rect 37946 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38262 37024
rect 37946 36959 38262 36960
rect 47946 37024 48262 37025
rect 47946 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48262 37024
rect 47946 36959 48262 36960
rect 48497 36954 48563 36957
rect 50200 36954 51000 36984
rect 48497 36952 51000 36954
rect 48497 36896 48502 36952
rect 48558 36896 51000 36952
rect 48497 36894 51000 36896
rect 48497 36891 48563 36894
rect 50200 36864 51000 36894
rect 0 36546 800 36576
rect 933 36546 999 36549
rect 0 36544 999 36546
rect 0 36488 938 36544
rect 994 36488 999 36544
rect 0 36486 999 36488
rect 0 36456 800 36486
rect 933 36483 999 36486
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 32946 36480 33262 36481
rect 32946 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33262 36480
rect 32946 36415 33262 36416
rect 42946 36480 43262 36481
rect 42946 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43262 36480
rect 42946 36415 43262 36416
rect 31845 36274 31911 36277
rect 38377 36274 38443 36277
rect 31845 36272 38443 36274
rect 31845 36216 31850 36272
rect 31906 36216 38382 36272
rect 38438 36216 38443 36272
rect 31845 36214 38443 36216
rect 31845 36211 31911 36214
rect 38377 36211 38443 36214
rect 49325 36274 49391 36277
rect 50200 36274 51000 36304
rect 49325 36272 51000 36274
rect 49325 36216 49330 36272
rect 49386 36216 51000 36272
rect 49325 36214 51000 36216
rect 49325 36211 49391 36214
rect 50200 36184 51000 36214
rect 32489 36138 32555 36141
rect 39389 36138 39455 36141
rect 32489 36136 39455 36138
rect 32489 36080 32494 36136
rect 32550 36080 39394 36136
rect 39450 36080 39455 36136
rect 32489 36078 39455 36080
rect 32489 36075 32555 36078
rect 39389 36075 39455 36078
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 27946 35936 28262 35937
rect 27946 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28262 35936
rect 27946 35871 28262 35872
rect 37946 35936 38262 35937
rect 37946 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38262 35936
rect 37946 35871 38262 35872
rect 47946 35936 48262 35937
rect 47946 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48262 35936
rect 47946 35871 48262 35872
rect 27705 35730 27771 35733
rect 28390 35730 28396 35732
rect 27705 35728 28396 35730
rect 27705 35672 27710 35728
rect 27766 35672 28396 35728
rect 27705 35670 28396 35672
rect 27705 35667 27771 35670
rect 28390 35668 28396 35670
rect 28460 35730 28466 35732
rect 32765 35730 32831 35733
rect 38377 35732 38443 35733
rect 28460 35728 32831 35730
rect 28460 35672 32770 35728
rect 32826 35672 32831 35728
rect 28460 35670 32831 35672
rect 28460 35668 28466 35670
rect 32765 35667 32831 35670
rect 38326 35668 38332 35732
rect 38396 35730 38443 35732
rect 38396 35728 38488 35730
rect 38438 35672 38488 35728
rect 38396 35670 38488 35672
rect 38396 35668 38443 35670
rect 38377 35667 38443 35668
rect 30097 35594 30163 35597
rect 39297 35594 39363 35597
rect 48589 35594 48655 35597
rect 30097 35592 48655 35594
rect 30097 35536 30102 35592
rect 30158 35536 39302 35592
rect 39358 35536 48594 35592
rect 48650 35536 48655 35592
rect 30097 35534 48655 35536
rect 30097 35531 30163 35534
rect 39297 35531 39363 35534
rect 48589 35531 48655 35534
rect 49325 35594 49391 35597
rect 50200 35594 51000 35624
rect 49325 35592 51000 35594
rect 49325 35536 49330 35592
rect 49386 35536 51000 35592
rect 49325 35534 51000 35536
rect 49325 35531 49391 35534
rect 50200 35504 51000 35534
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 32946 35392 33262 35393
rect 32946 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33262 35392
rect 32946 35327 33262 35328
rect 42946 35392 43262 35393
rect 42946 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43262 35392
rect 42946 35327 43262 35328
rect 17033 35186 17099 35189
rect 22737 35186 22803 35189
rect 30741 35186 30807 35189
rect 31293 35186 31359 35189
rect 17033 35184 19350 35186
rect 17033 35128 17038 35184
rect 17094 35128 19350 35184
rect 17033 35126 19350 35128
rect 17033 35123 17099 35126
rect 19290 35050 19350 35126
rect 22737 35184 31359 35186
rect 22737 35128 22742 35184
rect 22798 35128 30746 35184
rect 30802 35128 31298 35184
rect 31354 35128 31359 35184
rect 22737 35126 31359 35128
rect 22737 35123 22803 35126
rect 30741 35123 30807 35126
rect 31293 35123 31359 35126
rect 22461 35050 22527 35053
rect 31201 35050 31267 35053
rect 19290 35048 31267 35050
rect 19290 34992 22466 35048
rect 22522 34992 31206 35048
rect 31262 34992 31267 35048
rect 19290 34990 31267 34992
rect 22461 34987 22527 34990
rect 31201 34987 31267 34990
rect 31385 35050 31451 35053
rect 40861 35050 40927 35053
rect 31385 35048 40927 35050
rect 31385 34992 31390 35048
rect 31446 34992 40866 35048
rect 40922 34992 40927 35048
rect 31385 34990 40927 34992
rect 31385 34987 31451 34990
rect 40861 34987 40927 34990
rect 30373 34914 30439 34917
rect 33409 34914 33475 34917
rect 30373 34912 33475 34914
rect 30373 34856 30378 34912
rect 30434 34856 33414 34912
rect 33470 34856 33475 34912
rect 30373 34854 33475 34856
rect 30373 34851 30439 34854
rect 33409 34851 33475 34854
rect 49325 34914 49391 34917
rect 50200 34914 51000 34944
rect 49325 34912 51000 34914
rect 49325 34856 49330 34912
rect 49386 34856 51000 34912
rect 49325 34854 51000 34856
rect 49325 34851 49391 34854
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 27946 34848 28262 34849
rect 27946 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28262 34848
rect 27946 34783 28262 34784
rect 37946 34848 38262 34849
rect 37946 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38262 34848
rect 37946 34783 38262 34784
rect 47946 34848 48262 34849
rect 47946 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48262 34848
rect 50200 34824 51000 34854
rect 47946 34783 48262 34784
rect 28257 34642 28323 34645
rect 28574 34642 28580 34644
rect 28257 34640 28580 34642
rect 28257 34584 28262 34640
rect 28318 34584 28580 34640
rect 28257 34582 28580 34584
rect 28257 34579 28323 34582
rect 28574 34580 28580 34582
rect 28644 34580 28650 34644
rect 2946 34304 3262 34305
rect 0 34234 800 34264
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 32946 34304 33262 34305
rect 32946 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33262 34304
rect 32946 34239 33262 34240
rect 42946 34304 43262 34305
rect 42946 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43262 34304
rect 42946 34239 43262 34240
rect 1761 34234 1827 34237
rect 0 34232 1827 34234
rect 0 34176 1766 34232
rect 1822 34176 1827 34232
rect 0 34174 1827 34176
rect 0 34144 800 34174
rect 1761 34171 1827 34174
rect 49325 34234 49391 34237
rect 50200 34234 51000 34264
rect 49325 34232 51000 34234
rect 49325 34176 49330 34232
rect 49386 34176 51000 34232
rect 49325 34174 51000 34176
rect 49325 34171 49391 34174
rect 50200 34144 51000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 27946 33760 28262 33761
rect 27946 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28262 33760
rect 27946 33695 28262 33696
rect 37946 33760 38262 33761
rect 37946 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38262 33760
rect 37946 33695 38262 33696
rect 47946 33760 48262 33761
rect 47946 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48262 33760
rect 47946 33695 48262 33696
rect 37825 33554 37891 33557
rect 31710 33552 37891 33554
rect 31710 33496 37830 33552
rect 37886 33496 37891 33552
rect 31710 33494 37891 33496
rect 21265 33418 21331 33421
rect 26785 33418 26851 33421
rect 31710 33418 31770 33494
rect 37825 33491 37891 33494
rect 49325 33554 49391 33557
rect 50200 33554 51000 33584
rect 49325 33552 51000 33554
rect 49325 33496 49330 33552
rect 49386 33496 51000 33552
rect 49325 33494 51000 33496
rect 49325 33491 49391 33494
rect 50200 33464 51000 33494
rect 21265 33416 31770 33418
rect 21265 33360 21270 33416
rect 21326 33360 26790 33416
rect 26846 33360 31770 33416
rect 21265 33358 31770 33360
rect 36997 33418 37063 33421
rect 38193 33418 38259 33421
rect 36997 33416 38259 33418
rect 36997 33360 37002 33416
rect 37058 33360 38198 33416
rect 38254 33360 38259 33416
rect 36997 33358 38259 33360
rect 21265 33355 21331 33358
rect 26785 33355 26851 33358
rect 36997 33355 37063 33358
rect 38193 33355 38259 33358
rect 36905 33282 36971 33285
rect 37457 33282 37523 33285
rect 36905 33280 37523 33282
rect 36905 33224 36910 33280
rect 36966 33224 37462 33280
rect 37518 33224 37523 33280
rect 36905 33222 37523 33224
rect 36905 33219 36971 33222
rect 37457 33219 37523 33222
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 32946 33216 33262 33217
rect 32946 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33262 33216
rect 32946 33151 33262 33152
rect 42946 33216 43262 33217
rect 42946 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43262 33216
rect 42946 33151 43262 33152
rect 32765 33010 32831 33013
rect 35382 33010 35388 33012
rect 32765 33008 35388 33010
rect 32765 32952 32770 33008
rect 32826 32952 35388 33008
rect 32765 32950 35388 32952
rect 32765 32947 32831 32950
rect 35382 32948 35388 32950
rect 35452 32948 35458 33012
rect 26785 32874 26851 32877
rect 27102 32874 27108 32876
rect 26785 32872 27108 32874
rect 26785 32816 26790 32872
rect 26846 32816 27108 32872
rect 26785 32814 27108 32816
rect 26785 32811 26851 32814
rect 27102 32812 27108 32814
rect 27172 32812 27178 32876
rect 49325 32874 49391 32877
rect 50200 32874 51000 32904
rect 49325 32872 51000 32874
rect 49325 32816 49330 32872
rect 49386 32816 51000 32872
rect 49325 32814 51000 32816
rect 49325 32811 49391 32814
rect 50200 32784 51000 32814
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 27946 32672 28262 32673
rect 27946 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28262 32672
rect 27946 32607 28262 32608
rect 37946 32672 38262 32673
rect 37946 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38262 32672
rect 37946 32607 38262 32608
rect 47946 32672 48262 32673
rect 47946 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48262 32672
rect 47946 32607 48262 32608
rect 38285 32468 38351 32469
rect 38285 32464 38332 32468
rect 38396 32466 38402 32468
rect 38285 32408 38290 32464
rect 38285 32404 38332 32408
rect 38396 32406 38442 32466
rect 38396 32404 38402 32406
rect 38285 32403 38351 32404
rect 48497 32194 48563 32197
rect 50200 32194 51000 32224
rect 48497 32192 51000 32194
rect 48497 32136 48502 32192
rect 48558 32136 51000 32192
rect 48497 32134 51000 32136
rect 48497 32131 48563 32134
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 32946 32128 33262 32129
rect 32946 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33262 32128
rect 32946 32063 33262 32064
rect 42946 32128 43262 32129
rect 42946 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43262 32128
rect 50200 32104 51000 32134
rect 42946 32063 43262 32064
rect 36077 32058 36143 32061
rect 36629 32058 36695 32061
rect 36077 32056 36695 32058
rect 36077 32000 36082 32056
rect 36138 32000 36634 32056
rect 36690 32000 36695 32056
rect 36077 31998 36695 32000
rect 36077 31995 36143 31998
rect 36629 31995 36695 31998
rect 0 31922 800 31952
rect 933 31922 999 31925
rect 0 31920 999 31922
rect 0 31864 938 31920
rect 994 31864 999 31920
rect 0 31862 999 31864
rect 0 31832 800 31862
rect 933 31859 999 31862
rect 35985 31922 36051 31925
rect 40585 31922 40651 31925
rect 35985 31920 40651 31922
rect 35985 31864 35990 31920
rect 36046 31864 40590 31920
rect 40646 31864 40651 31920
rect 35985 31862 40651 31864
rect 35985 31859 36051 31862
rect 40585 31859 40651 31862
rect 38510 31724 38516 31788
rect 38580 31786 38586 31788
rect 38653 31786 38719 31789
rect 43989 31786 44055 31789
rect 38580 31784 44055 31786
rect 38580 31728 38658 31784
rect 38714 31728 43994 31784
rect 44050 31728 44055 31784
rect 38580 31726 44055 31728
rect 38580 31724 38586 31726
rect 38653 31723 38719 31726
rect 43989 31723 44055 31726
rect 28390 31588 28396 31652
rect 28460 31650 28466 31652
rect 28717 31650 28783 31653
rect 28460 31648 28783 31650
rect 28460 31592 28722 31648
rect 28778 31592 28783 31648
rect 28460 31590 28783 31592
rect 28460 31588 28466 31590
rect 28717 31587 28783 31590
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 27946 31584 28262 31585
rect 27946 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28262 31584
rect 27946 31519 28262 31520
rect 37946 31584 38262 31585
rect 37946 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38262 31584
rect 37946 31519 38262 31520
rect 47946 31584 48262 31585
rect 47946 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48262 31584
rect 47946 31519 48262 31520
rect 28574 31452 28580 31516
rect 28644 31514 28650 31516
rect 28717 31514 28783 31517
rect 28644 31512 28783 31514
rect 28644 31456 28722 31512
rect 28778 31456 28783 31512
rect 28644 31454 28783 31456
rect 28644 31452 28650 31454
rect 28717 31451 28783 31454
rect 34789 31514 34855 31517
rect 37733 31514 37799 31517
rect 34789 31512 37799 31514
rect 34789 31456 34794 31512
rect 34850 31456 37738 31512
rect 37794 31456 37799 31512
rect 34789 31454 37799 31456
rect 34789 31451 34855 31454
rect 37733 31451 37799 31454
rect 48497 31514 48563 31517
rect 50200 31514 51000 31544
rect 48497 31512 51000 31514
rect 48497 31456 48502 31512
rect 48558 31456 51000 31512
rect 48497 31454 51000 31456
rect 48497 31451 48563 31454
rect 50200 31424 51000 31454
rect 9765 31378 9831 31381
rect 34053 31378 34119 31381
rect 37549 31378 37615 31381
rect 9765 31376 12450 31378
rect 9765 31320 9770 31376
rect 9826 31320 12450 31376
rect 9765 31318 12450 31320
rect 9765 31315 9831 31318
rect 12390 31242 12450 31318
rect 34053 31376 37615 31378
rect 34053 31320 34058 31376
rect 34114 31320 37554 31376
rect 37610 31320 37615 31376
rect 34053 31318 37615 31320
rect 34053 31315 34119 31318
rect 37549 31315 37615 31318
rect 38193 31378 38259 31381
rect 39021 31378 39087 31381
rect 38193 31376 39087 31378
rect 38193 31320 38198 31376
rect 38254 31320 39026 31376
rect 39082 31320 39087 31376
rect 38193 31318 39087 31320
rect 38193 31315 38259 31318
rect 39021 31315 39087 31318
rect 22461 31242 22527 31245
rect 22686 31242 22692 31244
rect 12390 31240 22692 31242
rect 12390 31184 22466 31240
rect 22522 31184 22692 31240
rect 12390 31182 22692 31184
rect 22461 31179 22527 31182
rect 22686 31180 22692 31182
rect 22756 31180 22762 31244
rect 31017 31242 31083 31245
rect 35985 31242 36051 31245
rect 31017 31240 36051 31242
rect 31017 31184 31022 31240
rect 31078 31184 35990 31240
rect 36046 31184 36051 31240
rect 31017 31182 36051 31184
rect 31017 31179 31083 31182
rect 35985 31179 36051 31182
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 32946 31040 33262 31041
rect 32946 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33262 31040
rect 32946 30975 33262 30976
rect 42946 31040 43262 31041
rect 42946 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43262 31040
rect 42946 30975 43262 30976
rect 35893 30970 35959 30973
rect 36670 30970 36676 30972
rect 35893 30968 36676 30970
rect 35893 30912 35898 30968
rect 35954 30912 36676 30968
rect 35893 30910 36676 30912
rect 35893 30907 35959 30910
rect 36670 30908 36676 30910
rect 36740 30908 36746 30972
rect 22093 30834 22159 30837
rect 28717 30834 28783 30837
rect 22093 30832 28783 30834
rect 22093 30776 22098 30832
rect 22154 30776 28722 30832
rect 28778 30776 28783 30832
rect 22093 30774 28783 30776
rect 22093 30771 22159 30774
rect 28717 30771 28783 30774
rect 48497 30834 48563 30837
rect 50200 30834 51000 30864
rect 48497 30832 51000 30834
rect 48497 30776 48502 30832
rect 48558 30776 51000 30832
rect 48497 30774 51000 30776
rect 48497 30771 48563 30774
rect 50200 30744 51000 30774
rect 32397 30698 32463 30701
rect 39297 30698 39363 30701
rect 32397 30696 39363 30698
rect 32397 30640 32402 30696
rect 32458 30640 39302 30696
rect 39358 30640 39363 30696
rect 32397 30638 39363 30640
rect 32397 30635 32463 30638
rect 39297 30635 39363 30638
rect 34973 30562 35039 30565
rect 37273 30562 37339 30565
rect 34973 30560 37339 30562
rect 34973 30504 34978 30560
rect 35034 30504 37278 30560
rect 37334 30504 37339 30560
rect 34973 30502 37339 30504
rect 34973 30499 35039 30502
rect 37273 30499 37339 30502
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 27946 30496 28262 30497
rect 27946 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28262 30496
rect 27946 30431 28262 30432
rect 37946 30496 38262 30497
rect 37946 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38262 30496
rect 37946 30431 38262 30432
rect 47946 30496 48262 30497
rect 47946 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48262 30496
rect 47946 30431 48262 30432
rect 33869 30426 33935 30429
rect 36721 30426 36787 30429
rect 37222 30426 37228 30428
rect 33869 30424 37228 30426
rect 33869 30368 33874 30424
rect 33930 30368 36726 30424
rect 36782 30368 37228 30424
rect 33869 30366 37228 30368
rect 33869 30363 33935 30366
rect 36721 30363 36787 30366
rect 37222 30364 37228 30366
rect 37292 30364 37298 30428
rect 34145 30290 34211 30293
rect 35934 30290 35940 30292
rect 34145 30288 35940 30290
rect 34145 30232 34150 30288
rect 34206 30232 35940 30288
rect 34145 30230 35940 30232
rect 34145 30227 34211 30230
rect 35934 30228 35940 30230
rect 36004 30228 36010 30292
rect 49325 30154 49391 30157
rect 50200 30154 51000 30184
rect 49325 30152 51000 30154
rect 49325 30096 49330 30152
rect 49386 30096 51000 30152
rect 49325 30094 51000 30096
rect 49325 30091 49391 30094
rect 50200 30064 51000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 32946 29952 33262 29953
rect 32946 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33262 29952
rect 32946 29887 33262 29888
rect 42946 29952 43262 29953
rect 42946 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43262 29952
rect 42946 29887 43262 29888
rect 0 29610 800 29640
rect 1301 29610 1367 29613
rect 0 29608 1367 29610
rect 0 29552 1306 29608
rect 1362 29552 1367 29608
rect 0 29550 1367 29552
rect 0 29520 800 29550
rect 1301 29547 1367 29550
rect 48497 29474 48563 29477
rect 50200 29474 51000 29504
rect 48497 29472 51000 29474
rect 48497 29416 48502 29472
rect 48558 29416 51000 29472
rect 48497 29414 51000 29416
rect 48497 29411 48563 29414
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 27946 29408 28262 29409
rect 27946 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28262 29408
rect 27946 29343 28262 29344
rect 37946 29408 38262 29409
rect 37946 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38262 29408
rect 37946 29343 38262 29344
rect 47946 29408 48262 29409
rect 47946 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48262 29408
rect 50200 29384 51000 29414
rect 47946 29343 48262 29344
rect 23289 29202 23355 29205
rect 31201 29202 31267 29205
rect 23289 29200 31267 29202
rect 23289 29144 23294 29200
rect 23350 29144 31206 29200
rect 31262 29144 31267 29200
rect 23289 29142 31267 29144
rect 23289 29139 23355 29142
rect 31201 29139 31267 29142
rect 30005 29066 30071 29069
rect 30465 29066 30531 29069
rect 30005 29064 30531 29066
rect 30005 29008 30010 29064
rect 30066 29008 30470 29064
rect 30526 29008 30531 29064
rect 30005 29006 30531 29008
rect 30005 29003 30071 29006
rect 30465 29003 30531 29006
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 32946 28864 33262 28865
rect 32946 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33262 28864
rect 32946 28799 33262 28800
rect 42946 28864 43262 28865
rect 42946 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43262 28864
rect 42946 28799 43262 28800
rect 49325 28794 49391 28797
rect 50200 28794 51000 28824
rect 49325 28792 51000 28794
rect 49325 28736 49330 28792
rect 49386 28736 51000 28792
rect 49325 28734 51000 28736
rect 49325 28731 49391 28734
rect 50200 28704 51000 28734
rect 36813 28522 36879 28525
rect 40534 28522 40540 28524
rect 36813 28520 40540 28522
rect 36813 28464 36818 28520
rect 36874 28464 40540 28520
rect 36813 28462 40540 28464
rect 36813 28459 36879 28462
rect 40534 28460 40540 28462
rect 40604 28460 40610 28524
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 27946 28320 28262 28321
rect 27946 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28262 28320
rect 27946 28255 28262 28256
rect 37946 28320 38262 28321
rect 37946 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38262 28320
rect 37946 28255 38262 28256
rect 47946 28320 48262 28321
rect 47946 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48262 28320
rect 47946 28255 48262 28256
rect 23841 28114 23907 28117
rect 26233 28114 26299 28117
rect 23841 28112 26299 28114
rect 23841 28056 23846 28112
rect 23902 28056 26238 28112
rect 26294 28056 26299 28112
rect 23841 28054 26299 28056
rect 23841 28051 23907 28054
rect 26233 28051 26299 28054
rect 49325 28114 49391 28117
rect 50200 28114 51000 28144
rect 49325 28112 51000 28114
rect 49325 28056 49330 28112
rect 49386 28056 51000 28112
rect 49325 28054 51000 28056
rect 49325 28051 49391 28054
rect 50200 28024 51000 28054
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 32946 27776 33262 27777
rect 32946 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33262 27776
rect 32946 27711 33262 27712
rect 42946 27776 43262 27777
rect 42946 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43262 27776
rect 42946 27711 43262 27712
rect 28533 27570 28599 27573
rect 31017 27570 31083 27573
rect 35249 27570 35315 27573
rect 28533 27568 35315 27570
rect 28533 27512 28538 27568
rect 28594 27512 31022 27568
rect 31078 27512 35254 27568
rect 35310 27512 35315 27568
rect 28533 27510 35315 27512
rect 28533 27507 28599 27510
rect 31017 27507 31083 27510
rect 35249 27507 35315 27510
rect 32581 27434 32647 27437
rect 38510 27434 38516 27436
rect 32581 27432 38516 27434
rect 32581 27376 32586 27432
rect 32642 27376 38516 27432
rect 32581 27374 38516 27376
rect 32581 27371 32647 27374
rect 38510 27372 38516 27374
rect 38580 27372 38586 27436
rect 48497 27434 48563 27437
rect 50200 27434 51000 27464
rect 48497 27432 51000 27434
rect 48497 27376 48502 27432
rect 48558 27376 51000 27432
rect 48497 27374 51000 27376
rect 48497 27371 48563 27374
rect 50200 27344 51000 27374
rect 0 27298 800 27328
rect 1301 27298 1367 27301
rect 0 27296 1367 27298
rect 0 27240 1306 27296
rect 1362 27240 1367 27296
rect 0 27238 1367 27240
rect 0 27208 800 27238
rect 1301 27235 1367 27238
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 27946 27232 28262 27233
rect 27946 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28262 27232
rect 27946 27167 28262 27168
rect 37946 27232 38262 27233
rect 37946 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38262 27232
rect 37946 27167 38262 27168
rect 47946 27232 48262 27233
rect 47946 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48262 27232
rect 47946 27167 48262 27168
rect 31201 27162 31267 27165
rect 37365 27162 37431 27165
rect 31201 27160 37431 27162
rect 31201 27104 31206 27160
rect 31262 27104 37370 27160
rect 37426 27104 37431 27160
rect 31201 27102 37431 27104
rect 31201 27099 31267 27102
rect 37365 27099 37431 27102
rect 40585 27162 40651 27165
rect 42149 27162 42215 27165
rect 40585 27160 42215 27162
rect 40585 27104 40590 27160
rect 40646 27104 42154 27160
rect 42210 27104 42215 27160
rect 40585 27102 42215 27104
rect 40585 27099 40651 27102
rect 42149 27099 42215 27102
rect 33225 27026 33291 27029
rect 33685 27026 33751 27029
rect 37457 27026 37523 27029
rect 39982 27026 39988 27028
rect 33225 27024 39988 27026
rect 33225 26968 33230 27024
rect 33286 26968 33690 27024
rect 33746 26968 37462 27024
rect 37518 26968 39988 27024
rect 33225 26966 39988 26968
rect 33225 26963 33291 26966
rect 33685 26963 33751 26966
rect 37457 26963 37523 26966
rect 39982 26964 39988 26966
rect 40052 26964 40058 27028
rect 30598 26828 30604 26892
rect 30668 26890 30674 26892
rect 31293 26890 31359 26893
rect 30668 26888 31359 26890
rect 30668 26832 31298 26888
rect 31354 26832 31359 26888
rect 30668 26830 31359 26832
rect 30668 26828 30674 26830
rect 31293 26827 31359 26830
rect 48497 26754 48563 26757
rect 50200 26754 51000 26784
rect 48497 26752 51000 26754
rect 48497 26696 48502 26752
rect 48558 26696 51000 26752
rect 48497 26694 51000 26696
rect 48497 26691 48563 26694
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 32946 26688 33262 26689
rect 32946 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33262 26688
rect 32946 26623 33262 26624
rect 42946 26688 43262 26689
rect 42946 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43262 26688
rect 50200 26664 51000 26694
rect 42946 26623 43262 26624
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 27946 26144 28262 26145
rect 27946 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28262 26144
rect 27946 26079 28262 26080
rect 37946 26144 38262 26145
rect 37946 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38262 26144
rect 37946 26079 38262 26080
rect 47946 26144 48262 26145
rect 47946 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48262 26144
rect 47946 26079 48262 26080
rect 48405 26074 48471 26077
rect 50200 26074 51000 26104
rect 48405 26072 51000 26074
rect 48405 26016 48410 26072
rect 48466 26016 51000 26072
rect 48405 26014 51000 26016
rect 48405 26011 48471 26014
rect 50200 25984 51000 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 32946 25600 33262 25601
rect 32946 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33262 25600
rect 32946 25535 33262 25536
rect 42946 25600 43262 25601
rect 42946 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43262 25600
rect 42946 25535 43262 25536
rect 49325 25394 49391 25397
rect 50200 25394 51000 25424
rect 49325 25392 51000 25394
rect 49325 25336 49330 25392
rect 49386 25336 51000 25392
rect 49325 25334 51000 25336
rect 49325 25331 49391 25334
rect 50200 25304 51000 25334
rect 9489 25258 9555 25261
rect 30414 25258 30420 25260
rect 9489 25256 30420 25258
rect 9489 25200 9494 25256
rect 9550 25200 30420 25256
rect 9489 25198 30420 25200
rect 9489 25195 9555 25198
rect 30414 25196 30420 25198
rect 30484 25258 30490 25260
rect 32673 25258 32739 25261
rect 30484 25256 32739 25258
rect 30484 25200 32678 25256
rect 32734 25200 32739 25256
rect 30484 25198 32739 25200
rect 30484 25196 30490 25198
rect 32673 25195 32739 25198
rect 7946 25056 8262 25057
rect 0 24986 800 25016
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 27946 25056 28262 25057
rect 27946 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28262 25056
rect 27946 24991 28262 24992
rect 37946 25056 38262 25057
rect 37946 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38262 25056
rect 37946 24991 38262 24992
rect 47946 25056 48262 25057
rect 47946 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48262 25056
rect 47946 24991 48262 24992
rect 1301 24986 1367 24989
rect 0 24984 1367 24986
rect 0 24928 1306 24984
rect 1362 24928 1367 24984
rect 0 24926 1367 24928
rect 0 24896 800 24926
rect 1301 24923 1367 24926
rect 8937 24986 9003 24989
rect 9489 24986 9555 24989
rect 8937 24984 9555 24986
rect 8937 24928 8942 24984
rect 8998 24928 9494 24984
rect 9550 24928 9555 24984
rect 8937 24926 9555 24928
rect 8937 24923 9003 24926
rect 9489 24923 9555 24926
rect 26325 24850 26391 24853
rect 27889 24850 27955 24853
rect 28533 24850 28599 24853
rect 26325 24848 28599 24850
rect 26325 24792 26330 24848
rect 26386 24792 27894 24848
rect 27950 24792 28538 24848
rect 28594 24792 28599 24848
rect 26325 24790 28599 24792
rect 26325 24787 26391 24790
rect 27889 24787 27955 24790
rect 28533 24787 28599 24790
rect 25957 24716 26023 24717
rect 25957 24714 26004 24716
rect 25912 24712 26004 24714
rect 25912 24656 25962 24712
rect 25912 24654 26004 24656
rect 25957 24652 26004 24654
rect 26068 24652 26074 24716
rect 49141 24714 49207 24717
rect 50200 24714 51000 24744
rect 49141 24712 51000 24714
rect 49141 24656 49146 24712
rect 49202 24656 51000 24712
rect 49141 24654 51000 24656
rect 25957 24651 26023 24652
rect 49141 24651 49207 24654
rect 50200 24624 51000 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 25497 24306 25563 24309
rect 25630 24306 25636 24308
rect 25497 24304 25636 24306
rect 25497 24248 25502 24304
rect 25558 24248 25636 24304
rect 25497 24246 25636 24248
rect 25497 24243 25563 24246
rect 25630 24244 25636 24246
rect 25700 24244 25706 24308
rect 34881 24306 34947 24309
rect 34654 24304 34947 24306
rect 34654 24248 34886 24304
rect 34942 24248 34947 24304
rect 34654 24246 34947 24248
rect 34513 24170 34579 24173
rect 34654 24170 34714 24246
rect 34881 24243 34947 24246
rect 34513 24168 34714 24170
rect 34513 24112 34518 24168
rect 34574 24112 34714 24168
rect 34513 24110 34714 24112
rect 34513 24107 34579 24110
rect 49141 24034 49207 24037
rect 50200 24034 51000 24064
rect 49141 24032 51000 24034
rect 49141 23976 49146 24032
rect 49202 23976 51000 24032
rect 49141 23974 51000 23976
rect 49141 23971 49207 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 50200 23944 51000 23974
rect 47946 23903 48262 23904
rect 24853 23490 24919 23493
rect 28809 23490 28875 23493
rect 30097 23490 30163 23493
rect 24853 23488 30163 23490
rect 24853 23432 24858 23488
rect 24914 23432 28814 23488
rect 28870 23432 30102 23488
rect 30158 23432 30163 23488
rect 24853 23430 30163 23432
rect 24853 23427 24919 23430
rect 28809 23427 28875 23430
rect 30097 23427 30163 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 49141 23354 49207 23357
rect 50200 23354 51000 23384
rect 49141 23352 51000 23354
rect 49141 23296 49146 23352
rect 49202 23296 51000 23352
rect 49141 23294 51000 23296
rect 49141 23291 49207 23294
rect 50200 23264 51000 23294
rect 22686 22884 22692 22948
rect 22756 22946 22762 22948
rect 25037 22946 25103 22949
rect 22756 22944 25103 22946
rect 22756 22888 25042 22944
rect 25098 22888 25103 22944
rect 22756 22886 25103 22888
rect 22756 22884 22762 22886
rect 25037 22883 25103 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 0 22674 800 22704
rect 1301 22674 1367 22677
rect 0 22672 1367 22674
rect 0 22616 1306 22672
rect 1362 22616 1367 22672
rect 0 22614 1367 22616
rect 0 22584 800 22614
rect 1301 22611 1367 22614
rect 9581 22674 9647 22677
rect 30465 22674 30531 22677
rect 9581 22672 30531 22674
rect 9581 22616 9586 22672
rect 9642 22616 30470 22672
rect 30526 22616 30531 22672
rect 9581 22614 30531 22616
rect 9581 22611 9647 22614
rect 30465 22611 30531 22614
rect 49141 22674 49207 22677
rect 50200 22674 51000 22704
rect 49141 22672 51000 22674
rect 49141 22616 49146 22672
rect 49202 22616 51000 22672
rect 49141 22614 51000 22616
rect 49141 22611 49207 22614
rect 50200 22584 51000 22614
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 31937 21994 32003 21997
rect 32121 21994 32187 21997
rect 31937 21992 32187 21994
rect 31937 21936 31942 21992
rect 31998 21936 32126 21992
rect 32182 21936 32187 21992
rect 31937 21934 32187 21936
rect 31937 21931 32003 21934
rect 32121 21931 32187 21934
rect 49141 21994 49207 21997
rect 50200 21994 51000 22024
rect 49141 21992 51000 21994
rect 49141 21936 49146 21992
rect 49202 21936 51000 21992
rect 49141 21934 51000 21936
rect 49141 21931 49207 21934
rect 50200 21904 51000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 49141 21314 49207 21317
rect 50200 21314 51000 21344
rect 49141 21312 51000 21314
rect 49141 21256 49146 21312
rect 49202 21256 51000 21312
rect 49141 21254 51000 21256
rect 49141 21251 49207 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 50200 21224 51000 21254
rect 42946 21183 43262 21184
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 30465 20636 30531 20637
rect 30414 20572 30420 20636
rect 30484 20634 30531 20636
rect 49141 20634 49207 20637
rect 50200 20634 51000 20664
rect 30484 20632 30576 20634
rect 30526 20576 30576 20632
rect 30484 20574 30576 20576
rect 49141 20632 51000 20634
rect 49141 20576 49146 20632
rect 49202 20576 51000 20632
rect 49141 20574 51000 20576
rect 30484 20572 30531 20574
rect 30465 20571 30531 20572
rect 49141 20571 49207 20574
rect 50200 20544 51000 20574
rect 0 20362 800 20392
rect 1301 20362 1367 20365
rect 0 20360 1367 20362
rect 0 20304 1306 20360
rect 1362 20304 1367 20360
rect 0 20302 1367 20304
rect 0 20272 800 20302
rect 1301 20299 1367 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 49141 19954 49207 19957
rect 50200 19954 51000 19984
rect 49141 19952 51000 19954
rect 49141 19896 49146 19952
rect 49202 19896 51000 19952
rect 49141 19894 51000 19896
rect 49141 19891 49207 19894
rect 50200 19864 51000 19894
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 26734 19212 26740 19276
rect 26804 19274 26810 19276
rect 27245 19274 27311 19277
rect 31293 19274 31359 19277
rect 26804 19272 31359 19274
rect 26804 19216 27250 19272
rect 27306 19216 31298 19272
rect 31354 19216 31359 19272
rect 26804 19214 31359 19216
rect 26804 19212 26810 19214
rect 27245 19211 27311 19214
rect 31293 19211 31359 19214
rect 49141 19274 49207 19277
rect 50200 19274 51000 19304
rect 49141 19272 51000 19274
rect 49141 19216 49146 19272
rect 49202 19216 51000 19272
rect 49141 19214 51000 19216
rect 49141 19211 49207 19214
rect 50200 19184 51000 19214
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 27102 18804 27108 18868
rect 27172 18866 27178 18868
rect 28717 18866 28783 18869
rect 27172 18864 28783 18866
rect 27172 18808 28722 18864
rect 28778 18808 28783 18864
rect 27172 18806 28783 18808
rect 27172 18804 27178 18806
rect 28717 18803 28783 18806
rect 27705 18732 27771 18733
rect 27654 18668 27660 18732
rect 27724 18730 27771 18732
rect 27724 18728 27816 18730
rect 27766 18672 27816 18728
rect 27724 18670 27816 18672
rect 27724 18668 27771 18670
rect 27705 18667 27771 18668
rect 49141 18594 49207 18597
rect 50200 18594 51000 18624
rect 49141 18592 51000 18594
rect 49141 18536 49146 18592
rect 49202 18536 51000 18592
rect 49141 18534 51000 18536
rect 49141 18531 49207 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 50200 18504 51000 18534
rect 47946 18463 48262 18464
rect 0 18050 800 18080
rect 1301 18050 1367 18053
rect 0 18048 1367 18050
rect 0 17992 1306 18048
rect 1362 17992 1367 18048
rect 0 17990 1367 17992
rect 0 17960 800 17990
rect 1301 17987 1367 17990
rect 27889 18050 27955 18053
rect 30598 18050 30604 18052
rect 27889 18048 30604 18050
rect 27889 17992 27894 18048
rect 27950 17992 30604 18048
rect 27889 17990 30604 17992
rect 27889 17987 27955 17990
rect 30598 17988 30604 17990
rect 30668 17988 30674 18052
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 49141 17914 49207 17917
rect 50200 17914 51000 17944
rect 49141 17912 51000 17914
rect 49141 17856 49146 17912
rect 49202 17856 51000 17912
rect 49141 17854 51000 17856
rect 49141 17851 49207 17854
rect 50200 17824 51000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 49141 17234 49207 17237
rect 50200 17234 51000 17264
rect 49141 17232 51000 17234
rect 49141 17176 49146 17232
rect 49202 17176 51000 17232
rect 49141 17174 51000 17176
rect 49141 17171 49207 17174
rect 50200 17144 51000 17174
rect 27705 17100 27771 17101
rect 27654 17036 27660 17100
rect 27724 17098 27771 17100
rect 27724 17096 27816 17098
rect 27766 17040 27816 17096
rect 27724 17038 27816 17040
rect 27724 17036 27771 17038
rect 27705 17035 27771 17036
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 49141 16554 49207 16557
rect 50200 16554 51000 16584
rect 49141 16552 51000 16554
rect 49141 16496 49146 16552
rect 49202 16496 51000 16552
rect 49141 16494 51000 16496
rect 49141 16491 49207 16494
rect 50200 16464 51000 16494
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 49141 15874 49207 15877
rect 50200 15874 51000 15904
rect 49141 15872 51000 15874
rect 49141 15816 49146 15872
rect 49202 15816 51000 15872
rect 49141 15814 51000 15816
rect 49141 15811 49207 15814
rect 2946 15808 3262 15809
rect 0 15738 800 15768
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 50200 15784 51000 15814
rect 42946 15743 43262 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 27981 15602 28047 15605
rect 28809 15602 28875 15605
rect 27981 15600 28875 15602
rect 27981 15544 27986 15600
rect 28042 15544 28814 15600
rect 28870 15544 28875 15600
rect 27981 15542 28875 15544
rect 27981 15539 28047 15542
rect 28809 15539 28875 15542
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 49141 15194 49207 15197
rect 50200 15194 51000 15224
rect 49141 15192 51000 15194
rect 49141 15136 49146 15192
rect 49202 15136 51000 15192
rect 49141 15134 51000 15136
rect 49141 15131 49207 15134
rect 50200 15104 51000 15134
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 49141 14514 49207 14517
rect 50200 14514 51000 14544
rect 49141 14512 51000 14514
rect 49141 14456 49146 14512
rect 49202 14456 51000 14512
rect 49141 14454 51000 14456
rect 49141 14451 49207 14454
rect 50200 14424 51000 14454
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 49141 13834 49207 13837
rect 50200 13834 51000 13864
rect 49141 13832 51000 13834
rect 49141 13776 49146 13832
rect 49202 13776 51000 13832
rect 49141 13774 51000 13776
rect 49141 13771 49207 13774
rect 50200 13744 51000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 0 13426 800 13456
rect 2773 13426 2839 13429
rect 0 13424 2839 13426
rect 0 13368 2778 13424
rect 2834 13368 2839 13424
rect 0 13366 2839 13368
rect 0 13336 800 13366
rect 2773 13363 2839 13366
rect 49141 13154 49207 13157
rect 50200 13154 51000 13184
rect 49141 13152 51000 13154
rect 49141 13096 49146 13152
rect 49202 13096 51000 13152
rect 49141 13094 51000 13096
rect 49141 13091 49207 13094
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 50200 13064 51000 13094
rect 47946 13023 48262 13024
rect 28901 12882 28967 12885
rect 30598 12882 30604 12884
rect 28901 12880 30604 12882
rect 28901 12824 28906 12880
rect 28962 12824 30604 12880
rect 28901 12822 30604 12824
rect 28901 12819 28967 12822
rect 30598 12820 30604 12822
rect 30668 12820 30674 12884
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 49141 12411 49207 12414
rect 50200 12384 51000 12414
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 49141 11794 49207 11797
rect 50200 11794 51000 11824
rect 49141 11792 51000 11794
rect 49141 11736 49146 11792
rect 49202 11736 51000 11792
rect 49141 11734 51000 11736
rect 49141 11731 49207 11734
rect 50200 11704 51000 11734
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 0 11114 800 11144
rect 3417 11114 3483 11117
rect 0 11112 3483 11114
rect 0 11056 3422 11112
rect 3478 11056 3483 11112
rect 0 11054 3483 11056
rect 0 11024 800 11054
rect 3417 11051 3483 11054
rect 49141 11114 49207 11117
rect 50200 11114 51000 11144
rect 49141 11112 51000 11114
rect 49141 11056 49146 11112
rect 49202 11056 51000 11112
rect 49141 11054 51000 11056
rect 49141 11051 49207 11054
rect 50200 11024 51000 11054
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 49141 10434 49207 10437
rect 50200 10434 51000 10464
rect 49141 10432 51000 10434
rect 49141 10376 49146 10432
rect 49202 10376 51000 10432
rect 49141 10374 51000 10376
rect 49141 10371 49207 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 49141 9754 49207 9757
rect 50200 9754 51000 9784
rect 49141 9752 51000 9754
rect 49141 9696 49146 9752
rect 49202 9696 51000 9752
rect 49141 9694 51000 9696
rect 49141 9691 49207 9694
rect 50200 9664 51000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 49141 9074 49207 9077
rect 50200 9074 51000 9104
rect 49141 9072 51000 9074
rect 49141 9016 49146 9072
rect 49202 9016 51000 9072
rect 49141 9014 51000 9016
rect 49141 9011 49207 9014
rect 50200 8984 51000 9014
rect 0 8802 800 8832
rect 3325 8802 3391 8805
rect 0 8800 3391 8802
rect 0 8744 3330 8800
rect 3386 8744 3391 8800
rect 0 8742 3391 8744
rect 0 8712 800 8742
rect 3325 8739 3391 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 49141 8394 49207 8397
rect 50200 8394 51000 8424
rect 49141 8392 51000 8394
rect 49141 8336 49146 8392
rect 49202 8336 51000 8392
rect 49141 8334 51000 8336
rect 49141 8331 49207 8334
rect 50200 8304 51000 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 49141 7714 49207 7717
rect 50200 7714 51000 7744
rect 49141 7712 51000 7714
rect 49141 7656 49146 7712
rect 49202 7656 51000 7712
rect 49141 7654 51000 7656
rect 49141 7651 49207 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 50200 7624 51000 7654
rect 47946 7583 48262 7584
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 49141 7034 49207 7037
rect 50200 7034 51000 7064
rect 49141 7032 51000 7034
rect 49141 6976 49146 7032
rect 49202 6976 51000 7032
rect 49141 6974 51000 6976
rect 49141 6971 49207 6974
rect 50200 6944 51000 6974
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 3417 6490 3483 6493
rect 0 6488 3483 6490
rect 0 6432 3422 6488
rect 3478 6432 3483 6488
rect 0 6430 3483 6432
rect 0 6400 800 6430
rect 3417 6427 3483 6430
rect 49141 6354 49207 6357
rect 50200 6354 51000 6384
rect 49141 6352 51000 6354
rect 49141 6296 49146 6352
rect 49202 6296 51000 6352
rect 49141 6294 51000 6296
rect 49141 6291 49207 6294
rect 50200 6264 51000 6294
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5674 49207 5677
rect 50200 5674 51000 5704
rect 49141 5672 51000 5674
rect 49141 5616 49146 5672
rect 49202 5616 51000 5672
rect 49141 5614 51000 5616
rect 49141 5611 49207 5614
rect 50200 5584 51000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 49325 4994 49391 4997
rect 50200 4994 51000 5024
rect 49325 4992 51000 4994
rect 49325 4936 49330 4992
rect 49386 4936 51000 4992
rect 49325 4934 51000 4936
rect 49325 4931 49391 4934
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 50200 4904 51000 4934
rect 42946 4863 43262 4864
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4178 800 4208
rect 3417 4178 3483 4181
rect 0 4176 3483 4178
rect 0 4120 3422 4176
rect 3478 4120 3483 4176
rect 0 4118 3483 4120
rect 0 4088 800 4118
rect 3417 4115 3483 4118
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 17953 3090 18019 3093
rect 27102 3090 27108 3092
rect 17953 3088 27108 3090
rect 17953 3032 17958 3088
rect 18014 3032 27108 3088
rect 17953 3030 27108 3032
rect 17953 3027 18019 3030
rect 27102 3028 27108 3030
rect 27172 3028 27178 3092
rect 5441 2954 5507 2957
rect 22686 2954 22692 2956
rect 5441 2952 22692 2954
rect 5441 2896 5446 2952
rect 5502 2896 22692 2952
rect 5441 2894 22692 2896
rect 5441 2891 5507 2894
rect 22686 2892 22692 2894
rect 22756 2892 22762 2956
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 12341 2546 12407 2549
rect 27654 2546 27660 2548
rect 12341 2544 27660 2546
rect 12341 2488 12346 2544
rect 12402 2488 27660 2544
rect 12341 2486 27660 2488
rect 12341 2483 12407 2486
rect 27654 2484 27660 2486
rect 27724 2484 27730 2548
rect 5993 2410 6059 2413
rect 25998 2410 26004 2412
rect 5993 2408 26004 2410
rect 5993 2352 5998 2408
rect 6054 2352 26004 2408
rect 5993 2350 26004 2352
rect 5993 2347 6059 2350
rect 25998 2348 26004 2350
rect 26068 2348 26074 2412
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 15285 2002 15351 2005
rect 26734 2002 26740 2004
rect 15285 2000 26740 2002
rect 15285 1944 15290 2000
rect 15346 1944 26740 2000
rect 15285 1942 26740 1944
rect 15285 1939 15351 1942
rect 26734 1940 26740 1942
rect 26804 1940 26810 2004
rect 0 1866 800 1896
rect 2773 1866 2839 1869
rect 0 1864 2839 1866
rect 0 1808 2778 1864
rect 2834 1808 2839 1864
rect 0 1806 2839 1808
rect 0 1776 800 1806
rect 2773 1803 2839 1806
rect 11145 1866 11211 1869
rect 25630 1866 25636 1868
rect 11145 1864 25636 1866
rect 11145 1808 11150 1864
rect 11206 1808 25636 1864
rect 11145 1806 25636 1808
rect 11145 1803 11211 1806
rect 25630 1804 25636 1806
rect 25700 1804 25706 1868
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 27952 54428 28016 54432
rect 27952 54372 27956 54428
rect 27956 54372 28012 54428
rect 28012 54372 28016 54428
rect 27952 54368 28016 54372
rect 28032 54428 28096 54432
rect 28032 54372 28036 54428
rect 28036 54372 28092 54428
rect 28092 54372 28096 54428
rect 28032 54368 28096 54372
rect 28112 54428 28176 54432
rect 28112 54372 28116 54428
rect 28116 54372 28172 54428
rect 28172 54372 28176 54428
rect 28112 54368 28176 54372
rect 28192 54428 28256 54432
rect 28192 54372 28196 54428
rect 28196 54372 28252 54428
rect 28252 54372 28256 54428
rect 28192 54368 28256 54372
rect 37952 54428 38016 54432
rect 37952 54372 37956 54428
rect 37956 54372 38012 54428
rect 38012 54372 38016 54428
rect 37952 54368 38016 54372
rect 38032 54428 38096 54432
rect 38032 54372 38036 54428
rect 38036 54372 38092 54428
rect 38092 54372 38096 54428
rect 38032 54368 38096 54372
rect 38112 54428 38176 54432
rect 38112 54372 38116 54428
rect 38116 54372 38172 54428
rect 38172 54372 38176 54428
rect 38112 54368 38176 54372
rect 38192 54428 38256 54432
rect 38192 54372 38196 54428
rect 38196 54372 38252 54428
rect 38252 54372 38256 54428
rect 38192 54368 38256 54372
rect 47952 54428 48016 54432
rect 47952 54372 47956 54428
rect 47956 54372 48012 54428
rect 48012 54372 48016 54428
rect 47952 54368 48016 54372
rect 48032 54428 48096 54432
rect 48032 54372 48036 54428
rect 48036 54372 48092 54428
rect 48092 54372 48096 54428
rect 48032 54368 48096 54372
rect 48112 54428 48176 54432
rect 48112 54372 48116 54428
rect 48116 54372 48172 54428
rect 48172 54372 48176 54428
rect 48112 54368 48176 54372
rect 48192 54428 48256 54432
rect 48192 54372 48196 54428
rect 48196 54372 48252 54428
rect 48252 54372 48256 54428
rect 48192 54368 48256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 32952 53884 33016 53888
rect 32952 53828 32956 53884
rect 32956 53828 33012 53884
rect 33012 53828 33016 53884
rect 32952 53824 33016 53828
rect 33032 53884 33096 53888
rect 33032 53828 33036 53884
rect 33036 53828 33092 53884
rect 33092 53828 33096 53884
rect 33032 53824 33096 53828
rect 33112 53884 33176 53888
rect 33112 53828 33116 53884
rect 33116 53828 33172 53884
rect 33172 53828 33176 53884
rect 33112 53824 33176 53828
rect 33192 53884 33256 53888
rect 33192 53828 33196 53884
rect 33196 53828 33252 53884
rect 33252 53828 33256 53884
rect 33192 53824 33256 53828
rect 42952 53884 43016 53888
rect 42952 53828 42956 53884
rect 42956 53828 43012 53884
rect 43012 53828 43016 53884
rect 42952 53824 43016 53828
rect 43032 53884 43096 53888
rect 43032 53828 43036 53884
rect 43036 53828 43092 53884
rect 43092 53828 43096 53884
rect 43032 53824 43096 53828
rect 43112 53884 43176 53888
rect 43112 53828 43116 53884
rect 43116 53828 43172 53884
rect 43172 53828 43176 53884
rect 43112 53824 43176 53828
rect 43192 53884 43256 53888
rect 43192 53828 43196 53884
rect 43196 53828 43252 53884
rect 43252 53828 43256 53884
rect 43192 53824 43256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 27952 53340 28016 53344
rect 27952 53284 27956 53340
rect 27956 53284 28012 53340
rect 28012 53284 28016 53340
rect 27952 53280 28016 53284
rect 28032 53340 28096 53344
rect 28032 53284 28036 53340
rect 28036 53284 28092 53340
rect 28092 53284 28096 53340
rect 28032 53280 28096 53284
rect 28112 53340 28176 53344
rect 28112 53284 28116 53340
rect 28116 53284 28172 53340
rect 28172 53284 28176 53340
rect 28112 53280 28176 53284
rect 28192 53340 28256 53344
rect 28192 53284 28196 53340
rect 28196 53284 28252 53340
rect 28252 53284 28256 53340
rect 28192 53280 28256 53284
rect 37952 53340 38016 53344
rect 37952 53284 37956 53340
rect 37956 53284 38012 53340
rect 38012 53284 38016 53340
rect 37952 53280 38016 53284
rect 38032 53340 38096 53344
rect 38032 53284 38036 53340
rect 38036 53284 38092 53340
rect 38092 53284 38096 53340
rect 38032 53280 38096 53284
rect 38112 53340 38176 53344
rect 38112 53284 38116 53340
rect 38116 53284 38172 53340
rect 38172 53284 38176 53340
rect 38112 53280 38176 53284
rect 38192 53340 38256 53344
rect 38192 53284 38196 53340
rect 38196 53284 38252 53340
rect 38252 53284 38256 53340
rect 38192 53280 38256 53284
rect 47952 53340 48016 53344
rect 47952 53284 47956 53340
rect 47956 53284 48012 53340
rect 48012 53284 48016 53340
rect 47952 53280 48016 53284
rect 48032 53340 48096 53344
rect 48032 53284 48036 53340
rect 48036 53284 48092 53340
rect 48092 53284 48096 53340
rect 48032 53280 48096 53284
rect 48112 53340 48176 53344
rect 48112 53284 48116 53340
rect 48116 53284 48172 53340
rect 48172 53284 48176 53340
rect 48112 53280 48176 53284
rect 48192 53340 48256 53344
rect 48192 53284 48196 53340
rect 48196 53284 48252 53340
rect 48252 53284 48256 53340
rect 48192 53280 48256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 32952 52796 33016 52800
rect 32952 52740 32956 52796
rect 32956 52740 33012 52796
rect 33012 52740 33016 52796
rect 32952 52736 33016 52740
rect 33032 52796 33096 52800
rect 33032 52740 33036 52796
rect 33036 52740 33092 52796
rect 33092 52740 33096 52796
rect 33032 52736 33096 52740
rect 33112 52796 33176 52800
rect 33112 52740 33116 52796
rect 33116 52740 33172 52796
rect 33172 52740 33176 52796
rect 33112 52736 33176 52740
rect 33192 52796 33256 52800
rect 33192 52740 33196 52796
rect 33196 52740 33252 52796
rect 33252 52740 33256 52796
rect 33192 52736 33256 52740
rect 42952 52796 43016 52800
rect 42952 52740 42956 52796
rect 42956 52740 43012 52796
rect 43012 52740 43016 52796
rect 42952 52736 43016 52740
rect 43032 52796 43096 52800
rect 43032 52740 43036 52796
rect 43036 52740 43092 52796
rect 43092 52740 43096 52796
rect 43032 52736 43096 52740
rect 43112 52796 43176 52800
rect 43112 52740 43116 52796
rect 43116 52740 43172 52796
rect 43172 52740 43176 52796
rect 43112 52736 43176 52740
rect 43192 52796 43256 52800
rect 43192 52740 43196 52796
rect 43196 52740 43252 52796
rect 43252 52740 43256 52796
rect 43192 52736 43256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 27952 52252 28016 52256
rect 27952 52196 27956 52252
rect 27956 52196 28012 52252
rect 28012 52196 28016 52252
rect 27952 52192 28016 52196
rect 28032 52252 28096 52256
rect 28032 52196 28036 52252
rect 28036 52196 28092 52252
rect 28092 52196 28096 52252
rect 28032 52192 28096 52196
rect 28112 52252 28176 52256
rect 28112 52196 28116 52252
rect 28116 52196 28172 52252
rect 28172 52196 28176 52252
rect 28112 52192 28176 52196
rect 28192 52252 28256 52256
rect 28192 52196 28196 52252
rect 28196 52196 28252 52252
rect 28252 52196 28256 52252
rect 28192 52192 28256 52196
rect 37952 52252 38016 52256
rect 37952 52196 37956 52252
rect 37956 52196 38012 52252
rect 38012 52196 38016 52252
rect 37952 52192 38016 52196
rect 38032 52252 38096 52256
rect 38032 52196 38036 52252
rect 38036 52196 38092 52252
rect 38092 52196 38096 52252
rect 38032 52192 38096 52196
rect 38112 52252 38176 52256
rect 38112 52196 38116 52252
rect 38116 52196 38172 52252
rect 38172 52196 38176 52252
rect 38112 52192 38176 52196
rect 38192 52252 38256 52256
rect 38192 52196 38196 52252
rect 38196 52196 38252 52252
rect 38252 52196 38256 52252
rect 38192 52192 38256 52196
rect 47952 52252 48016 52256
rect 47952 52196 47956 52252
rect 47956 52196 48012 52252
rect 48012 52196 48016 52252
rect 47952 52192 48016 52196
rect 48032 52252 48096 52256
rect 48032 52196 48036 52252
rect 48036 52196 48092 52252
rect 48092 52196 48096 52252
rect 48032 52192 48096 52196
rect 48112 52252 48176 52256
rect 48112 52196 48116 52252
rect 48116 52196 48172 52252
rect 48172 52196 48176 52252
rect 48112 52192 48176 52196
rect 48192 52252 48256 52256
rect 48192 52196 48196 52252
rect 48196 52196 48252 52252
rect 48252 52196 48256 52252
rect 48192 52192 48256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 32952 51708 33016 51712
rect 32952 51652 32956 51708
rect 32956 51652 33012 51708
rect 33012 51652 33016 51708
rect 32952 51648 33016 51652
rect 33032 51708 33096 51712
rect 33032 51652 33036 51708
rect 33036 51652 33092 51708
rect 33092 51652 33096 51708
rect 33032 51648 33096 51652
rect 33112 51708 33176 51712
rect 33112 51652 33116 51708
rect 33116 51652 33172 51708
rect 33172 51652 33176 51708
rect 33112 51648 33176 51652
rect 33192 51708 33256 51712
rect 33192 51652 33196 51708
rect 33196 51652 33252 51708
rect 33252 51652 33256 51708
rect 33192 51648 33256 51652
rect 42952 51708 43016 51712
rect 42952 51652 42956 51708
rect 42956 51652 43012 51708
rect 43012 51652 43016 51708
rect 42952 51648 43016 51652
rect 43032 51708 43096 51712
rect 43032 51652 43036 51708
rect 43036 51652 43092 51708
rect 43092 51652 43096 51708
rect 43032 51648 43096 51652
rect 43112 51708 43176 51712
rect 43112 51652 43116 51708
rect 43116 51652 43172 51708
rect 43172 51652 43176 51708
rect 43112 51648 43176 51652
rect 43192 51708 43256 51712
rect 43192 51652 43196 51708
rect 43196 51652 43252 51708
rect 43252 51652 43256 51708
rect 43192 51648 43256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 27952 51164 28016 51168
rect 27952 51108 27956 51164
rect 27956 51108 28012 51164
rect 28012 51108 28016 51164
rect 27952 51104 28016 51108
rect 28032 51164 28096 51168
rect 28032 51108 28036 51164
rect 28036 51108 28092 51164
rect 28092 51108 28096 51164
rect 28032 51104 28096 51108
rect 28112 51164 28176 51168
rect 28112 51108 28116 51164
rect 28116 51108 28172 51164
rect 28172 51108 28176 51164
rect 28112 51104 28176 51108
rect 28192 51164 28256 51168
rect 28192 51108 28196 51164
rect 28196 51108 28252 51164
rect 28252 51108 28256 51164
rect 28192 51104 28256 51108
rect 37952 51164 38016 51168
rect 37952 51108 37956 51164
rect 37956 51108 38012 51164
rect 38012 51108 38016 51164
rect 37952 51104 38016 51108
rect 38032 51164 38096 51168
rect 38032 51108 38036 51164
rect 38036 51108 38092 51164
rect 38092 51108 38096 51164
rect 38032 51104 38096 51108
rect 38112 51164 38176 51168
rect 38112 51108 38116 51164
rect 38116 51108 38172 51164
rect 38172 51108 38176 51164
rect 38112 51104 38176 51108
rect 38192 51164 38256 51168
rect 38192 51108 38196 51164
rect 38196 51108 38252 51164
rect 38252 51108 38256 51164
rect 38192 51104 38256 51108
rect 47952 51164 48016 51168
rect 47952 51108 47956 51164
rect 47956 51108 48012 51164
rect 48012 51108 48016 51164
rect 47952 51104 48016 51108
rect 48032 51164 48096 51168
rect 48032 51108 48036 51164
rect 48036 51108 48092 51164
rect 48092 51108 48096 51164
rect 48032 51104 48096 51108
rect 48112 51164 48176 51168
rect 48112 51108 48116 51164
rect 48116 51108 48172 51164
rect 48172 51108 48176 51164
rect 48112 51104 48176 51108
rect 48192 51164 48256 51168
rect 48192 51108 48196 51164
rect 48196 51108 48252 51164
rect 48252 51108 48256 51164
rect 48192 51104 48256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 32952 50620 33016 50624
rect 32952 50564 32956 50620
rect 32956 50564 33012 50620
rect 33012 50564 33016 50620
rect 32952 50560 33016 50564
rect 33032 50620 33096 50624
rect 33032 50564 33036 50620
rect 33036 50564 33092 50620
rect 33092 50564 33096 50620
rect 33032 50560 33096 50564
rect 33112 50620 33176 50624
rect 33112 50564 33116 50620
rect 33116 50564 33172 50620
rect 33172 50564 33176 50620
rect 33112 50560 33176 50564
rect 33192 50620 33256 50624
rect 33192 50564 33196 50620
rect 33196 50564 33252 50620
rect 33252 50564 33256 50620
rect 33192 50560 33256 50564
rect 42952 50620 43016 50624
rect 42952 50564 42956 50620
rect 42956 50564 43012 50620
rect 43012 50564 43016 50620
rect 42952 50560 43016 50564
rect 43032 50620 43096 50624
rect 43032 50564 43036 50620
rect 43036 50564 43092 50620
rect 43092 50564 43096 50620
rect 43032 50560 43096 50564
rect 43112 50620 43176 50624
rect 43112 50564 43116 50620
rect 43116 50564 43172 50620
rect 43172 50564 43176 50620
rect 43112 50560 43176 50564
rect 43192 50620 43256 50624
rect 43192 50564 43196 50620
rect 43196 50564 43252 50620
rect 43252 50564 43256 50620
rect 43192 50560 43256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 27952 50076 28016 50080
rect 27952 50020 27956 50076
rect 27956 50020 28012 50076
rect 28012 50020 28016 50076
rect 27952 50016 28016 50020
rect 28032 50076 28096 50080
rect 28032 50020 28036 50076
rect 28036 50020 28092 50076
rect 28092 50020 28096 50076
rect 28032 50016 28096 50020
rect 28112 50076 28176 50080
rect 28112 50020 28116 50076
rect 28116 50020 28172 50076
rect 28172 50020 28176 50076
rect 28112 50016 28176 50020
rect 28192 50076 28256 50080
rect 28192 50020 28196 50076
rect 28196 50020 28252 50076
rect 28252 50020 28256 50076
rect 28192 50016 28256 50020
rect 37952 50076 38016 50080
rect 37952 50020 37956 50076
rect 37956 50020 38012 50076
rect 38012 50020 38016 50076
rect 37952 50016 38016 50020
rect 38032 50076 38096 50080
rect 38032 50020 38036 50076
rect 38036 50020 38092 50076
rect 38092 50020 38096 50076
rect 38032 50016 38096 50020
rect 38112 50076 38176 50080
rect 38112 50020 38116 50076
rect 38116 50020 38172 50076
rect 38172 50020 38176 50076
rect 38112 50016 38176 50020
rect 38192 50076 38256 50080
rect 38192 50020 38196 50076
rect 38196 50020 38252 50076
rect 38252 50020 38256 50076
rect 38192 50016 38256 50020
rect 47952 50076 48016 50080
rect 47952 50020 47956 50076
rect 47956 50020 48012 50076
rect 48012 50020 48016 50076
rect 47952 50016 48016 50020
rect 48032 50076 48096 50080
rect 48032 50020 48036 50076
rect 48036 50020 48092 50076
rect 48092 50020 48096 50076
rect 48032 50016 48096 50020
rect 48112 50076 48176 50080
rect 48112 50020 48116 50076
rect 48116 50020 48172 50076
rect 48172 50020 48176 50076
rect 48112 50016 48176 50020
rect 48192 50076 48256 50080
rect 48192 50020 48196 50076
rect 48196 50020 48252 50076
rect 48252 50020 48256 50076
rect 48192 50016 48256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 32952 49532 33016 49536
rect 32952 49476 32956 49532
rect 32956 49476 33012 49532
rect 33012 49476 33016 49532
rect 32952 49472 33016 49476
rect 33032 49532 33096 49536
rect 33032 49476 33036 49532
rect 33036 49476 33092 49532
rect 33092 49476 33096 49532
rect 33032 49472 33096 49476
rect 33112 49532 33176 49536
rect 33112 49476 33116 49532
rect 33116 49476 33172 49532
rect 33172 49476 33176 49532
rect 33112 49472 33176 49476
rect 33192 49532 33256 49536
rect 33192 49476 33196 49532
rect 33196 49476 33252 49532
rect 33252 49476 33256 49532
rect 33192 49472 33256 49476
rect 42952 49532 43016 49536
rect 42952 49476 42956 49532
rect 42956 49476 43012 49532
rect 43012 49476 43016 49532
rect 42952 49472 43016 49476
rect 43032 49532 43096 49536
rect 43032 49476 43036 49532
rect 43036 49476 43092 49532
rect 43092 49476 43096 49532
rect 43032 49472 43096 49476
rect 43112 49532 43176 49536
rect 43112 49476 43116 49532
rect 43116 49476 43172 49532
rect 43172 49476 43176 49532
rect 43112 49472 43176 49476
rect 43192 49532 43256 49536
rect 43192 49476 43196 49532
rect 43196 49476 43252 49532
rect 43252 49476 43256 49532
rect 43192 49472 43256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 27952 48988 28016 48992
rect 27952 48932 27956 48988
rect 27956 48932 28012 48988
rect 28012 48932 28016 48988
rect 27952 48928 28016 48932
rect 28032 48988 28096 48992
rect 28032 48932 28036 48988
rect 28036 48932 28092 48988
rect 28092 48932 28096 48988
rect 28032 48928 28096 48932
rect 28112 48988 28176 48992
rect 28112 48932 28116 48988
rect 28116 48932 28172 48988
rect 28172 48932 28176 48988
rect 28112 48928 28176 48932
rect 28192 48988 28256 48992
rect 28192 48932 28196 48988
rect 28196 48932 28252 48988
rect 28252 48932 28256 48988
rect 28192 48928 28256 48932
rect 37952 48988 38016 48992
rect 37952 48932 37956 48988
rect 37956 48932 38012 48988
rect 38012 48932 38016 48988
rect 37952 48928 38016 48932
rect 38032 48988 38096 48992
rect 38032 48932 38036 48988
rect 38036 48932 38092 48988
rect 38092 48932 38096 48988
rect 38032 48928 38096 48932
rect 38112 48988 38176 48992
rect 38112 48932 38116 48988
rect 38116 48932 38172 48988
rect 38172 48932 38176 48988
rect 38112 48928 38176 48932
rect 38192 48988 38256 48992
rect 38192 48932 38196 48988
rect 38196 48932 38252 48988
rect 38252 48932 38256 48988
rect 38192 48928 38256 48932
rect 47952 48988 48016 48992
rect 47952 48932 47956 48988
rect 47956 48932 48012 48988
rect 48012 48932 48016 48988
rect 47952 48928 48016 48932
rect 48032 48988 48096 48992
rect 48032 48932 48036 48988
rect 48036 48932 48092 48988
rect 48092 48932 48096 48988
rect 48032 48928 48096 48932
rect 48112 48988 48176 48992
rect 48112 48932 48116 48988
rect 48116 48932 48172 48988
rect 48172 48932 48176 48988
rect 48112 48928 48176 48932
rect 48192 48988 48256 48992
rect 48192 48932 48196 48988
rect 48196 48932 48252 48988
rect 48252 48932 48256 48988
rect 48192 48928 48256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 32952 48444 33016 48448
rect 32952 48388 32956 48444
rect 32956 48388 33012 48444
rect 33012 48388 33016 48444
rect 32952 48384 33016 48388
rect 33032 48444 33096 48448
rect 33032 48388 33036 48444
rect 33036 48388 33092 48444
rect 33092 48388 33096 48444
rect 33032 48384 33096 48388
rect 33112 48444 33176 48448
rect 33112 48388 33116 48444
rect 33116 48388 33172 48444
rect 33172 48388 33176 48444
rect 33112 48384 33176 48388
rect 33192 48444 33256 48448
rect 33192 48388 33196 48444
rect 33196 48388 33252 48444
rect 33252 48388 33256 48444
rect 33192 48384 33256 48388
rect 42952 48444 43016 48448
rect 42952 48388 42956 48444
rect 42956 48388 43012 48444
rect 43012 48388 43016 48444
rect 42952 48384 43016 48388
rect 43032 48444 43096 48448
rect 43032 48388 43036 48444
rect 43036 48388 43092 48444
rect 43092 48388 43096 48444
rect 43032 48384 43096 48388
rect 43112 48444 43176 48448
rect 43112 48388 43116 48444
rect 43116 48388 43172 48444
rect 43172 48388 43176 48444
rect 43112 48384 43176 48388
rect 43192 48444 43256 48448
rect 43192 48388 43196 48444
rect 43196 48388 43252 48444
rect 43252 48388 43256 48444
rect 43192 48384 43256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 27952 47900 28016 47904
rect 27952 47844 27956 47900
rect 27956 47844 28012 47900
rect 28012 47844 28016 47900
rect 27952 47840 28016 47844
rect 28032 47900 28096 47904
rect 28032 47844 28036 47900
rect 28036 47844 28092 47900
rect 28092 47844 28096 47900
rect 28032 47840 28096 47844
rect 28112 47900 28176 47904
rect 28112 47844 28116 47900
rect 28116 47844 28172 47900
rect 28172 47844 28176 47900
rect 28112 47840 28176 47844
rect 28192 47900 28256 47904
rect 28192 47844 28196 47900
rect 28196 47844 28252 47900
rect 28252 47844 28256 47900
rect 28192 47840 28256 47844
rect 37952 47900 38016 47904
rect 37952 47844 37956 47900
rect 37956 47844 38012 47900
rect 38012 47844 38016 47900
rect 37952 47840 38016 47844
rect 38032 47900 38096 47904
rect 38032 47844 38036 47900
rect 38036 47844 38092 47900
rect 38092 47844 38096 47900
rect 38032 47840 38096 47844
rect 38112 47900 38176 47904
rect 38112 47844 38116 47900
rect 38116 47844 38172 47900
rect 38172 47844 38176 47900
rect 38112 47840 38176 47844
rect 38192 47900 38256 47904
rect 38192 47844 38196 47900
rect 38196 47844 38252 47900
rect 38252 47844 38256 47900
rect 38192 47840 38256 47844
rect 47952 47900 48016 47904
rect 47952 47844 47956 47900
rect 47956 47844 48012 47900
rect 48012 47844 48016 47900
rect 47952 47840 48016 47844
rect 48032 47900 48096 47904
rect 48032 47844 48036 47900
rect 48036 47844 48092 47900
rect 48092 47844 48096 47900
rect 48032 47840 48096 47844
rect 48112 47900 48176 47904
rect 48112 47844 48116 47900
rect 48116 47844 48172 47900
rect 48172 47844 48176 47900
rect 48112 47840 48176 47844
rect 48192 47900 48256 47904
rect 48192 47844 48196 47900
rect 48196 47844 48252 47900
rect 48252 47844 48256 47900
rect 48192 47840 48256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 32952 47356 33016 47360
rect 32952 47300 32956 47356
rect 32956 47300 33012 47356
rect 33012 47300 33016 47356
rect 32952 47296 33016 47300
rect 33032 47356 33096 47360
rect 33032 47300 33036 47356
rect 33036 47300 33092 47356
rect 33092 47300 33096 47356
rect 33032 47296 33096 47300
rect 33112 47356 33176 47360
rect 33112 47300 33116 47356
rect 33116 47300 33172 47356
rect 33172 47300 33176 47356
rect 33112 47296 33176 47300
rect 33192 47356 33256 47360
rect 33192 47300 33196 47356
rect 33196 47300 33252 47356
rect 33252 47300 33256 47356
rect 33192 47296 33256 47300
rect 42952 47356 43016 47360
rect 42952 47300 42956 47356
rect 42956 47300 43012 47356
rect 43012 47300 43016 47356
rect 42952 47296 43016 47300
rect 43032 47356 43096 47360
rect 43032 47300 43036 47356
rect 43036 47300 43092 47356
rect 43092 47300 43096 47356
rect 43032 47296 43096 47300
rect 43112 47356 43176 47360
rect 43112 47300 43116 47356
rect 43116 47300 43172 47356
rect 43172 47300 43176 47356
rect 43112 47296 43176 47300
rect 43192 47356 43256 47360
rect 43192 47300 43196 47356
rect 43196 47300 43252 47356
rect 43252 47300 43256 47356
rect 43192 47296 43256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 27952 46812 28016 46816
rect 27952 46756 27956 46812
rect 27956 46756 28012 46812
rect 28012 46756 28016 46812
rect 27952 46752 28016 46756
rect 28032 46812 28096 46816
rect 28032 46756 28036 46812
rect 28036 46756 28092 46812
rect 28092 46756 28096 46812
rect 28032 46752 28096 46756
rect 28112 46812 28176 46816
rect 28112 46756 28116 46812
rect 28116 46756 28172 46812
rect 28172 46756 28176 46812
rect 28112 46752 28176 46756
rect 28192 46812 28256 46816
rect 28192 46756 28196 46812
rect 28196 46756 28252 46812
rect 28252 46756 28256 46812
rect 28192 46752 28256 46756
rect 37952 46812 38016 46816
rect 37952 46756 37956 46812
rect 37956 46756 38012 46812
rect 38012 46756 38016 46812
rect 37952 46752 38016 46756
rect 38032 46812 38096 46816
rect 38032 46756 38036 46812
rect 38036 46756 38092 46812
rect 38092 46756 38096 46812
rect 38032 46752 38096 46756
rect 38112 46812 38176 46816
rect 38112 46756 38116 46812
rect 38116 46756 38172 46812
rect 38172 46756 38176 46812
rect 38112 46752 38176 46756
rect 38192 46812 38256 46816
rect 38192 46756 38196 46812
rect 38196 46756 38252 46812
rect 38252 46756 38256 46812
rect 38192 46752 38256 46756
rect 47952 46812 48016 46816
rect 47952 46756 47956 46812
rect 47956 46756 48012 46812
rect 48012 46756 48016 46812
rect 47952 46752 48016 46756
rect 48032 46812 48096 46816
rect 48032 46756 48036 46812
rect 48036 46756 48092 46812
rect 48092 46756 48096 46812
rect 48032 46752 48096 46756
rect 48112 46812 48176 46816
rect 48112 46756 48116 46812
rect 48116 46756 48172 46812
rect 48172 46756 48176 46812
rect 48112 46752 48176 46756
rect 48192 46812 48256 46816
rect 48192 46756 48196 46812
rect 48196 46756 48252 46812
rect 48252 46756 48256 46812
rect 48192 46752 48256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 32952 46268 33016 46272
rect 32952 46212 32956 46268
rect 32956 46212 33012 46268
rect 33012 46212 33016 46268
rect 32952 46208 33016 46212
rect 33032 46268 33096 46272
rect 33032 46212 33036 46268
rect 33036 46212 33092 46268
rect 33092 46212 33096 46268
rect 33032 46208 33096 46212
rect 33112 46268 33176 46272
rect 33112 46212 33116 46268
rect 33116 46212 33172 46268
rect 33172 46212 33176 46268
rect 33112 46208 33176 46212
rect 33192 46268 33256 46272
rect 33192 46212 33196 46268
rect 33196 46212 33252 46268
rect 33252 46212 33256 46268
rect 33192 46208 33256 46212
rect 42952 46268 43016 46272
rect 42952 46212 42956 46268
rect 42956 46212 43012 46268
rect 43012 46212 43016 46268
rect 42952 46208 43016 46212
rect 43032 46268 43096 46272
rect 43032 46212 43036 46268
rect 43036 46212 43092 46268
rect 43092 46212 43096 46268
rect 43032 46208 43096 46212
rect 43112 46268 43176 46272
rect 43112 46212 43116 46268
rect 43116 46212 43172 46268
rect 43172 46212 43176 46268
rect 43112 46208 43176 46212
rect 43192 46268 43256 46272
rect 43192 46212 43196 46268
rect 43196 46212 43252 46268
rect 43252 46212 43256 46268
rect 43192 46208 43256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 27952 45724 28016 45728
rect 27952 45668 27956 45724
rect 27956 45668 28012 45724
rect 28012 45668 28016 45724
rect 27952 45664 28016 45668
rect 28032 45724 28096 45728
rect 28032 45668 28036 45724
rect 28036 45668 28092 45724
rect 28092 45668 28096 45724
rect 28032 45664 28096 45668
rect 28112 45724 28176 45728
rect 28112 45668 28116 45724
rect 28116 45668 28172 45724
rect 28172 45668 28176 45724
rect 28112 45664 28176 45668
rect 28192 45724 28256 45728
rect 28192 45668 28196 45724
rect 28196 45668 28252 45724
rect 28252 45668 28256 45724
rect 28192 45664 28256 45668
rect 37952 45724 38016 45728
rect 37952 45668 37956 45724
rect 37956 45668 38012 45724
rect 38012 45668 38016 45724
rect 37952 45664 38016 45668
rect 38032 45724 38096 45728
rect 38032 45668 38036 45724
rect 38036 45668 38092 45724
rect 38092 45668 38096 45724
rect 38032 45664 38096 45668
rect 38112 45724 38176 45728
rect 38112 45668 38116 45724
rect 38116 45668 38172 45724
rect 38172 45668 38176 45724
rect 38112 45664 38176 45668
rect 38192 45724 38256 45728
rect 38192 45668 38196 45724
rect 38196 45668 38252 45724
rect 38252 45668 38256 45724
rect 38192 45664 38256 45668
rect 47952 45724 48016 45728
rect 47952 45668 47956 45724
rect 47956 45668 48012 45724
rect 48012 45668 48016 45724
rect 47952 45664 48016 45668
rect 48032 45724 48096 45728
rect 48032 45668 48036 45724
rect 48036 45668 48092 45724
rect 48092 45668 48096 45724
rect 48032 45664 48096 45668
rect 48112 45724 48176 45728
rect 48112 45668 48116 45724
rect 48116 45668 48172 45724
rect 48172 45668 48176 45724
rect 48112 45664 48176 45668
rect 48192 45724 48256 45728
rect 48192 45668 48196 45724
rect 48196 45668 48252 45724
rect 48252 45668 48256 45724
rect 48192 45664 48256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 32952 45180 33016 45184
rect 32952 45124 32956 45180
rect 32956 45124 33012 45180
rect 33012 45124 33016 45180
rect 32952 45120 33016 45124
rect 33032 45180 33096 45184
rect 33032 45124 33036 45180
rect 33036 45124 33092 45180
rect 33092 45124 33096 45180
rect 33032 45120 33096 45124
rect 33112 45180 33176 45184
rect 33112 45124 33116 45180
rect 33116 45124 33172 45180
rect 33172 45124 33176 45180
rect 33112 45120 33176 45124
rect 33192 45180 33256 45184
rect 33192 45124 33196 45180
rect 33196 45124 33252 45180
rect 33252 45124 33256 45180
rect 33192 45120 33256 45124
rect 42952 45180 43016 45184
rect 42952 45124 42956 45180
rect 42956 45124 43012 45180
rect 43012 45124 43016 45180
rect 42952 45120 43016 45124
rect 43032 45180 43096 45184
rect 43032 45124 43036 45180
rect 43036 45124 43092 45180
rect 43092 45124 43096 45180
rect 43032 45120 43096 45124
rect 43112 45180 43176 45184
rect 43112 45124 43116 45180
rect 43116 45124 43172 45180
rect 43172 45124 43176 45180
rect 43112 45120 43176 45124
rect 43192 45180 43256 45184
rect 43192 45124 43196 45180
rect 43196 45124 43252 45180
rect 43252 45124 43256 45180
rect 43192 45120 43256 45124
rect 35388 44644 35452 44708
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 27952 44636 28016 44640
rect 27952 44580 27956 44636
rect 27956 44580 28012 44636
rect 28012 44580 28016 44636
rect 27952 44576 28016 44580
rect 28032 44636 28096 44640
rect 28032 44580 28036 44636
rect 28036 44580 28092 44636
rect 28092 44580 28096 44636
rect 28032 44576 28096 44580
rect 28112 44636 28176 44640
rect 28112 44580 28116 44636
rect 28116 44580 28172 44636
rect 28172 44580 28176 44636
rect 28112 44576 28176 44580
rect 28192 44636 28256 44640
rect 28192 44580 28196 44636
rect 28196 44580 28252 44636
rect 28252 44580 28256 44636
rect 28192 44576 28256 44580
rect 37952 44636 38016 44640
rect 37952 44580 37956 44636
rect 37956 44580 38012 44636
rect 38012 44580 38016 44636
rect 37952 44576 38016 44580
rect 38032 44636 38096 44640
rect 38032 44580 38036 44636
rect 38036 44580 38092 44636
rect 38092 44580 38096 44636
rect 38032 44576 38096 44580
rect 38112 44636 38176 44640
rect 38112 44580 38116 44636
rect 38116 44580 38172 44636
rect 38172 44580 38176 44636
rect 38112 44576 38176 44580
rect 38192 44636 38256 44640
rect 38192 44580 38196 44636
rect 38196 44580 38252 44636
rect 38252 44580 38256 44636
rect 38192 44576 38256 44580
rect 47952 44636 48016 44640
rect 47952 44580 47956 44636
rect 47956 44580 48012 44636
rect 48012 44580 48016 44636
rect 47952 44576 48016 44580
rect 48032 44636 48096 44640
rect 48032 44580 48036 44636
rect 48036 44580 48092 44636
rect 48092 44580 48096 44636
rect 48032 44576 48096 44580
rect 48112 44636 48176 44640
rect 48112 44580 48116 44636
rect 48116 44580 48172 44636
rect 48172 44580 48176 44636
rect 48112 44576 48176 44580
rect 48192 44636 48256 44640
rect 48192 44580 48196 44636
rect 48196 44580 48252 44636
rect 48252 44580 48256 44636
rect 48192 44576 48256 44580
rect 36676 44236 36740 44300
rect 37228 44236 37292 44300
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 32952 44092 33016 44096
rect 32952 44036 32956 44092
rect 32956 44036 33012 44092
rect 33012 44036 33016 44092
rect 32952 44032 33016 44036
rect 33032 44092 33096 44096
rect 33032 44036 33036 44092
rect 33036 44036 33092 44092
rect 33092 44036 33096 44092
rect 33032 44032 33096 44036
rect 33112 44092 33176 44096
rect 33112 44036 33116 44092
rect 33116 44036 33172 44092
rect 33172 44036 33176 44092
rect 33112 44032 33176 44036
rect 33192 44092 33256 44096
rect 33192 44036 33196 44092
rect 33196 44036 33252 44092
rect 33252 44036 33256 44092
rect 33192 44032 33256 44036
rect 42952 44092 43016 44096
rect 42952 44036 42956 44092
rect 42956 44036 43012 44092
rect 43012 44036 43016 44092
rect 42952 44032 43016 44036
rect 43032 44092 43096 44096
rect 43032 44036 43036 44092
rect 43036 44036 43092 44092
rect 43092 44036 43096 44092
rect 43032 44032 43096 44036
rect 43112 44092 43176 44096
rect 43112 44036 43116 44092
rect 43116 44036 43172 44092
rect 43172 44036 43176 44092
rect 43112 44032 43176 44036
rect 43192 44092 43256 44096
rect 43192 44036 43196 44092
rect 43196 44036 43252 44092
rect 43252 44036 43256 44092
rect 43192 44032 43256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 27952 43548 28016 43552
rect 27952 43492 27956 43548
rect 27956 43492 28012 43548
rect 28012 43492 28016 43548
rect 27952 43488 28016 43492
rect 28032 43548 28096 43552
rect 28032 43492 28036 43548
rect 28036 43492 28092 43548
rect 28092 43492 28096 43548
rect 28032 43488 28096 43492
rect 28112 43548 28176 43552
rect 28112 43492 28116 43548
rect 28116 43492 28172 43548
rect 28172 43492 28176 43548
rect 28112 43488 28176 43492
rect 28192 43548 28256 43552
rect 28192 43492 28196 43548
rect 28196 43492 28252 43548
rect 28252 43492 28256 43548
rect 28192 43488 28256 43492
rect 37952 43548 38016 43552
rect 37952 43492 37956 43548
rect 37956 43492 38012 43548
rect 38012 43492 38016 43548
rect 37952 43488 38016 43492
rect 38032 43548 38096 43552
rect 38032 43492 38036 43548
rect 38036 43492 38092 43548
rect 38092 43492 38096 43548
rect 38032 43488 38096 43492
rect 38112 43548 38176 43552
rect 38112 43492 38116 43548
rect 38116 43492 38172 43548
rect 38172 43492 38176 43548
rect 38112 43488 38176 43492
rect 38192 43548 38256 43552
rect 38192 43492 38196 43548
rect 38196 43492 38252 43548
rect 38252 43492 38256 43548
rect 38192 43488 38256 43492
rect 47952 43548 48016 43552
rect 47952 43492 47956 43548
rect 47956 43492 48012 43548
rect 48012 43492 48016 43548
rect 47952 43488 48016 43492
rect 48032 43548 48096 43552
rect 48032 43492 48036 43548
rect 48036 43492 48092 43548
rect 48092 43492 48096 43548
rect 48032 43488 48096 43492
rect 48112 43548 48176 43552
rect 48112 43492 48116 43548
rect 48116 43492 48172 43548
rect 48172 43492 48176 43548
rect 48112 43488 48176 43492
rect 48192 43548 48256 43552
rect 48192 43492 48196 43548
rect 48196 43492 48252 43548
rect 48252 43492 48256 43548
rect 48192 43488 48256 43492
rect 35940 43420 36004 43484
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 32952 43004 33016 43008
rect 32952 42948 32956 43004
rect 32956 42948 33012 43004
rect 33012 42948 33016 43004
rect 32952 42944 33016 42948
rect 33032 43004 33096 43008
rect 33032 42948 33036 43004
rect 33036 42948 33092 43004
rect 33092 42948 33096 43004
rect 33032 42944 33096 42948
rect 33112 43004 33176 43008
rect 33112 42948 33116 43004
rect 33116 42948 33172 43004
rect 33172 42948 33176 43004
rect 33112 42944 33176 42948
rect 33192 43004 33256 43008
rect 33192 42948 33196 43004
rect 33196 42948 33252 43004
rect 33252 42948 33256 43004
rect 33192 42944 33256 42948
rect 42952 43004 43016 43008
rect 42952 42948 42956 43004
rect 42956 42948 43012 43004
rect 43012 42948 43016 43004
rect 42952 42944 43016 42948
rect 43032 43004 43096 43008
rect 43032 42948 43036 43004
rect 43036 42948 43092 43004
rect 43092 42948 43096 43004
rect 43032 42944 43096 42948
rect 43112 43004 43176 43008
rect 43112 42948 43116 43004
rect 43116 42948 43172 43004
rect 43172 42948 43176 43004
rect 43112 42944 43176 42948
rect 43192 43004 43256 43008
rect 43192 42948 43196 43004
rect 43196 42948 43252 43004
rect 43252 42948 43256 43004
rect 43192 42944 43256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 27952 42460 28016 42464
rect 27952 42404 27956 42460
rect 27956 42404 28012 42460
rect 28012 42404 28016 42460
rect 27952 42400 28016 42404
rect 28032 42460 28096 42464
rect 28032 42404 28036 42460
rect 28036 42404 28092 42460
rect 28092 42404 28096 42460
rect 28032 42400 28096 42404
rect 28112 42460 28176 42464
rect 28112 42404 28116 42460
rect 28116 42404 28172 42460
rect 28172 42404 28176 42460
rect 28112 42400 28176 42404
rect 28192 42460 28256 42464
rect 28192 42404 28196 42460
rect 28196 42404 28252 42460
rect 28252 42404 28256 42460
rect 28192 42400 28256 42404
rect 37952 42460 38016 42464
rect 37952 42404 37956 42460
rect 37956 42404 38012 42460
rect 38012 42404 38016 42460
rect 37952 42400 38016 42404
rect 38032 42460 38096 42464
rect 38032 42404 38036 42460
rect 38036 42404 38092 42460
rect 38092 42404 38096 42460
rect 38032 42400 38096 42404
rect 38112 42460 38176 42464
rect 38112 42404 38116 42460
rect 38116 42404 38172 42460
rect 38172 42404 38176 42460
rect 38112 42400 38176 42404
rect 38192 42460 38256 42464
rect 38192 42404 38196 42460
rect 38196 42404 38252 42460
rect 38252 42404 38256 42460
rect 38192 42400 38256 42404
rect 47952 42460 48016 42464
rect 47952 42404 47956 42460
rect 47956 42404 48012 42460
rect 48012 42404 48016 42460
rect 47952 42400 48016 42404
rect 48032 42460 48096 42464
rect 48032 42404 48036 42460
rect 48036 42404 48092 42460
rect 48092 42404 48096 42460
rect 48032 42400 48096 42404
rect 48112 42460 48176 42464
rect 48112 42404 48116 42460
rect 48116 42404 48172 42460
rect 48172 42404 48176 42460
rect 48112 42400 48176 42404
rect 48192 42460 48256 42464
rect 48192 42404 48196 42460
rect 48196 42404 48252 42460
rect 48252 42404 48256 42460
rect 48192 42400 48256 42404
rect 39988 42060 40052 42124
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 32952 41916 33016 41920
rect 32952 41860 32956 41916
rect 32956 41860 33012 41916
rect 33012 41860 33016 41916
rect 32952 41856 33016 41860
rect 33032 41916 33096 41920
rect 33032 41860 33036 41916
rect 33036 41860 33092 41916
rect 33092 41860 33096 41916
rect 33032 41856 33096 41860
rect 33112 41916 33176 41920
rect 33112 41860 33116 41916
rect 33116 41860 33172 41916
rect 33172 41860 33176 41916
rect 33112 41856 33176 41860
rect 33192 41916 33256 41920
rect 33192 41860 33196 41916
rect 33196 41860 33252 41916
rect 33252 41860 33256 41916
rect 33192 41856 33256 41860
rect 42952 41916 43016 41920
rect 42952 41860 42956 41916
rect 42956 41860 43012 41916
rect 43012 41860 43016 41916
rect 42952 41856 43016 41860
rect 43032 41916 43096 41920
rect 43032 41860 43036 41916
rect 43036 41860 43092 41916
rect 43092 41860 43096 41916
rect 43032 41856 43096 41860
rect 43112 41916 43176 41920
rect 43112 41860 43116 41916
rect 43116 41860 43172 41916
rect 43172 41860 43176 41916
rect 43112 41856 43176 41860
rect 43192 41916 43256 41920
rect 43192 41860 43196 41916
rect 43196 41860 43252 41916
rect 43252 41860 43256 41916
rect 43192 41856 43256 41860
rect 40540 41652 40604 41716
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 27952 41372 28016 41376
rect 27952 41316 27956 41372
rect 27956 41316 28012 41372
rect 28012 41316 28016 41372
rect 27952 41312 28016 41316
rect 28032 41372 28096 41376
rect 28032 41316 28036 41372
rect 28036 41316 28092 41372
rect 28092 41316 28096 41372
rect 28032 41312 28096 41316
rect 28112 41372 28176 41376
rect 28112 41316 28116 41372
rect 28116 41316 28172 41372
rect 28172 41316 28176 41372
rect 28112 41312 28176 41316
rect 28192 41372 28256 41376
rect 28192 41316 28196 41372
rect 28196 41316 28252 41372
rect 28252 41316 28256 41372
rect 28192 41312 28256 41316
rect 37952 41372 38016 41376
rect 37952 41316 37956 41372
rect 37956 41316 38012 41372
rect 38012 41316 38016 41372
rect 37952 41312 38016 41316
rect 38032 41372 38096 41376
rect 38032 41316 38036 41372
rect 38036 41316 38092 41372
rect 38092 41316 38096 41372
rect 38032 41312 38096 41316
rect 38112 41372 38176 41376
rect 38112 41316 38116 41372
rect 38116 41316 38172 41372
rect 38172 41316 38176 41372
rect 38112 41312 38176 41316
rect 38192 41372 38256 41376
rect 38192 41316 38196 41372
rect 38196 41316 38252 41372
rect 38252 41316 38256 41372
rect 38192 41312 38256 41316
rect 47952 41372 48016 41376
rect 47952 41316 47956 41372
rect 47956 41316 48012 41372
rect 48012 41316 48016 41372
rect 47952 41312 48016 41316
rect 48032 41372 48096 41376
rect 48032 41316 48036 41372
rect 48036 41316 48092 41372
rect 48092 41316 48096 41372
rect 48032 41312 48096 41316
rect 48112 41372 48176 41376
rect 48112 41316 48116 41372
rect 48116 41316 48172 41372
rect 48172 41316 48176 41372
rect 48112 41312 48176 41316
rect 48192 41372 48256 41376
rect 48192 41316 48196 41372
rect 48196 41316 48252 41372
rect 48252 41316 48256 41372
rect 48192 41312 48256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 32952 40828 33016 40832
rect 32952 40772 32956 40828
rect 32956 40772 33012 40828
rect 33012 40772 33016 40828
rect 32952 40768 33016 40772
rect 33032 40828 33096 40832
rect 33032 40772 33036 40828
rect 33036 40772 33092 40828
rect 33092 40772 33096 40828
rect 33032 40768 33096 40772
rect 33112 40828 33176 40832
rect 33112 40772 33116 40828
rect 33116 40772 33172 40828
rect 33172 40772 33176 40828
rect 33112 40768 33176 40772
rect 33192 40828 33256 40832
rect 33192 40772 33196 40828
rect 33196 40772 33252 40828
rect 33252 40772 33256 40828
rect 33192 40768 33256 40772
rect 42952 40828 43016 40832
rect 42952 40772 42956 40828
rect 42956 40772 43012 40828
rect 43012 40772 43016 40828
rect 42952 40768 43016 40772
rect 43032 40828 43096 40832
rect 43032 40772 43036 40828
rect 43036 40772 43092 40828
rect 43092 40772 43096 40828
rect 43032 40768 43096 40772
rect 43112 40828 43176 40832
rect 43112 40772 43116 40828
rect 43116 40772 43172 40828
rect 43172 40772 43176 40828
rect 43112 40768 43176 40772
rect 43192 40828 43256 40832
rect 43192 40772 43196 40828
rect 43196 40772 43252 40828
rect 43252 40772 43256 40828
rect 43192 40768 43256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 27952 40284 28016 40288
rect 27952 40228 27956 40284
rect 27956 40228 28012 40284
rect 28012 40228 28016 40284
rect 27952 40224 28016 40228
rect 28032 40284 28096 40288
rect 28032 40228 28036 40284
rect 28036 40228 28092 40284
rect 28092 40228 28096 40284
rect 28032 40224 28096 40228
rect 28112 40284 28176 40288
rect 28112 40228 28116 40284
rect 28116 40228 28172 40284
rect 28172 40228 28176 40284
rect 28112 40224 28176 40228
rect 28192 40284 28256 40288
rect 28192 40228 28196 40284
rect 28196 40228 28252 40284
rect 28252 40228 28256 40284
rect 28192 40224 28256 40228
rect 37952 40284 38016 40288
rect 37952 40228 37956 40284
rect 37956 40228 38012 40284
rect 38012 40228 38016 40284
rect 37952 40224 38016 40228
rect 38032 40284 38096 40288
rect 38032 40228 38036 40284
rect 38036 40228 38092 40284
rect 38092 40228 38096 40284
rect 38032 40224 38096 40228
rect 38112 40284 38176 40288
rect 38112 40228 38116 40284
rect 38116 40228 38172 40284
rect 38172 40228 38176 40284
rect 38112 40224 38176 40228
rect 38192 40284 38256 40288
rect 38192 40228 38196 40284
rect 38196 40228 38252 40284
rect 38252 40228 38256 40284
rect 38192 40224 38256 40228
rect 47952 40284 48016 40288
rect 47952 40228 47956 40284
rect 47956 40228 48012 40284
rect 48012 40228 48016 40284
rect 47952 40224 48016 40228
rect 48032 40284 48096 40288
rect 48032 40228 48036 40284
rect 48036 40228 48092 40284
rect 48092 40228 48096 40284
rect 48032 40224 48096 40228
rect 48112 40284 48176 40288
rect 48112 40228 48116 40284
rect 48116 40228 48172 40284
rect 48172 40228 48176 40284
rect 48112 40224 48176 40228
rect 48192 40284 48256 40288
rect 48192 40228 48196 40284
rect 48196 40228 48252 40284
rect 48252 40228 48256 40284
rect 48192 40224 48256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 32952 39740 33016 39744
rect 32952 39684 32956 39740
rect 32956 39684 33012 39740
rect 33012 39684 33016 39740
rect 32952 39680 33016 39684
rect 33032 39740 33096 39744
rect 33032 39684 33036 39740
rect 33036 39684 33092 39740
rect 33092 39684 33096 39740
rect 33032 39680 33096 39684
rect 33112 39740 33176 39744
rect 33112 39684 33116 39740
rect 33116 39684 33172 39740
rect 33172 39684 33176 39740
rect 33112 39680 33176 39684
rect 33192 39740 33256 39744
rect 33192 39684 33196 39740
rect 33196 39684 33252 39740
rect 33252 39684 33256 39740
rect 33192 39680 33256 39684
rect 42952 39740 43016 39744
rect 42952 39684 42956 39740
rect 42956 39684 43012 39740
rect 43012 39684 43016 39740
rect 42952 39680 43016 39684
rect 43032 39740 43096 39744
rect 43032 39684 43036 39740
rect 43036 39684 43092 39740
rect 43092 39684 43096 39740
rect 43032 39680 43096 39684
rect 43112 39740 43176 39744
rect 43112 39684 43116 39740
rect 43116 39684 43172 39740
rect 43172 39684 43176 39740
rect 43112 39680 43176 39684
rect 43192 39740 43256 39744
rect 43192 39684 43196 39740
rect 43196 39684 43252 39740
rect 43252 39684 43256 39740
rect 43192 39680 43256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 27952 39196 28016 39200
rect 27952 39140 27956 39196
rect 27956 39140 28012 39196
rect 28012 39140 28016 39196
rect 27952 39136 28016 39140
rect 28032 39196 28096 39200
rect 28032 39140 28036 39196
rect 28036 39140 28092 39196
rect 28092 39140 28096 39196
rect 28032 39136 28096 39140
rect 28112 39196 28176 39200
rect 28112 39140 28116 39196
rect 28116 39140 28172 39196
rect 28172 39140 28176 39196
rect 28112 39136 28176 39140
rect 28192 39196 28256 39200
rect 28192 39140 28196 39196
rect 28196 39140 28252 39196
rect 28252 39140 28256 39196
rect 28192 39136 28256 39140
rect 37952 39196 38016 39200
rect 37952 39140 37956 39196
rect 37956 39140 38012 39196
rect 38012 39140 38016 39196
rect 37952 39136 38016 39140
rect 38032 39196 38096 39200
rect 38032 39140 38036 39196
rect 38036 39140 38092 39196
rect 38092 39140 38096 39196
rect 38032 39136 38096 39140
rect 38112 39196 38176 39200
rect 38112 39140 38116 39196
rect 38116 39140 38172 39196
rect 38172 39140 38176 39196
rect 38112 39136 38176 39140
rect 38192 39196 38256 39200
rect 38192 39140 38196 39196
rect 38196 39140 38252 39196
rect 38252 39140 38256 39196
rect 38192 39136 38256 39140
rect 47952 39196 48016 39200
rect 47952 39140 47956 39196
rect 47956 39140 48012 39196
rect 48012 39140 48016 39196
rect 47952 39136 48016 39140
rect 48032 39196 48096 39200
rect 48032 39140 48036 39196
rect 48036 39140 48092 39196
rect 48092 39140 48096 39196
rect 48032 39136 48096 39140
rect 48112 39196 48176 39200
rect 48112 39140 48116 39196
rect 48116 39140 48172 39196
rect 48172 39140 48176 39196
rect 48112 39136 48176 39140
rect 48192 39196 48256 39200
rect 48192 39140 48196 39196
rect 48196 39140 48252 39196
rect 48252 39140 48256 39196
rect 48192 39136 48256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 32952 38652 33016 38656
rect 32952 38596 32956 38652
rect 32956 38596 33012 38652
rect 33012 38596 33016 38652
rect 32952 38592 33016 38596
rect 33032 38652 33096 38656
rect 33032 38596 33036 38652
rect 33036 38596 33092 38652
rect 33092 38596 33096 38652
rect 33032 38592 33096 38596
rect 33112 38652 33176 38656
rect 33112 38596 33116 38652
rect 33116 38596 33172 38652
rect 33172 38596 33176 38652
rect 33112 38592 33176 38596
rect 33192 38652 33256 38656
rect 33192 38596 33196 38652
rect 33196 38596 33252 38652
rect 33252 38596 33256 38652
rect 33192 38592 33256 38596
rect 42952 38652 43016 38656
rect 42952 38596 42956 38652
rect 42956 38596 43012 38652
rect 43012 38596 43016 38652
rect 42952 38592 43016 38596
rect 43032 38652 43096 38656
rect 43032 38596 43036 38652
rect 43036 38596 43092 38652
rect 43092 38596 43096 38652
rect 43032 38592 43096 38596
rect 43112 38652 43176 38656
rect 43112 38596 43116 38652
rect 43116 38596 43172 38652
rect 43172 38596 43176 38652
rect 43112 38592 43176 38596
rect 43192 38652 43256 38656
rect 43192 38596 43196 38652
rect 43196 38596 43252 38652
rect 43252 38596 43256 38652
rect 43192 38592 43256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 27952 38108 28016 38112
rect 27952 38052 27956 38108
rect 27956 38052 28012 38108
rect 28012 38052 28016 38108
rect 27952 38048 28016 38052
rect 28032 38108 28096 38112
rect 28032 38052 28036 38108
rect 28036 38052 28092 38108
rect 28092 38052 28096 38108
rect 28032 38048 28096 38052
rect 28112 38108 28176 38112
rect 28112 38052 28116 38108
rect 28116 38052 28172 38108
rect 28172 38052 28176 38108
rect 28112 38048 28176 38052
rect 28192 38108 28256 38112
rect 28192 38052 28196 38108
rect 28196 38052 28252 38108
rect 28252 38052 28256 38108
rect 28192 38048 28256 38052
rect 37952 38108 38016 38112
rect 37952 38052 37956 38108
rect 37956 38052 38012 38108
rect 38012 38052 38016 38108
rect 37952 38048 38016 38052
rect 38032 38108 38096 38112
rect 38032 38052 38036 38108
rect 38036 38052 38092 38108
rect 38092 38052 38096 38108
rect 38032 38048 38096 38052
rect 38112 38108 38176 38112
rect 38112 38052 38116 38108
rect 38116 38052 38172 38108
rect 38172 38052 38176 38108
rect 38112 38048 38176 38052
rect 38192 38108 38256 38112
rect 38192 38052 38196 38108
rect 38196 38052 38252 38108
rect 38252 38052 38256 38108
rect 38192 38048 38256 38052
rect 47952 38108 48016 38112
rect 47952 38052 47956 38108
rect 47956 38052 48012 38108
rect 48012 38052 48016 38108
rect 47952 38048 48016 38052
rect 48032 38108 48096 38112
rect 48032 38052 48036 38108
rect 48036 38052 48092 38108
rect 48092 38052 48096 38108
rect 48032 38048 48096 38052
rect 48112 38108 48176 38112
rect 48112 38052 48116 38108
rect 48116 38052 48172 38108
rect 48172 38052 48176 38108
rect 48112 38048 48176 38052
rect 48192 38108 48256 38112
rect 48192 38052 48196 38108
rect 48196 38052 48252 38108
rect 48252 38052 48256 38108
rect 48192 38048 48256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 32952 37564 33016 37568
rect 32952 37508 32956 37564
rect 32956 37508 33012 37564
rect 33012 37508 33016 37564
rect 32952 37504 33016 37508
rect 33032 37564 33096 37568
rect 33032 37508 33036 37564
rect 33036 37508 33092 37564
rect 33092 37508 33096 37564
rect 33032 37504 33096 37508
rect 33112 37564 33176 37568
rect 33112 37508 33116 37564
rect 33116 37508 33172 37564
rect 33172 37508 33176 37564
rect 33112 37504 33176 37508
rect 33192 37564 33256 37568
rect 33192 37508 33196 37564
rect 33196 37508 33252 37564
rect 33252 37508 33256 37564
rect 33192 37504 33256 37508
rect 42952 37564 43016 37568
rect 42952 37508 42956 37564
rect 42956 37508 43012 37564
rect 43012 37508 43016 37564
rect 42952 37504 43016 37508
rect 43032 37564 43096 37568
rect 43032 37508 43036 37564
rect 43036 37508 43092 37564
rect 43092 37508 43096 37564
rect 43032 37504 43096 37508
rect 43112 37564 43176 37568
rect 43112 37508 43116 37564
rect 43116 37508 43172 37564
rect 43172 37508 43176 37564
rect 43112 37504 43176 37508
rect 43192 37564 43256 37568
rect 43192 37508 43196 37564
rect 43196 37508 43252 37564
rect 43252 37508 43256 37564
rect 43192 37504 43256 37508
rect 25636 37164 25700 37228
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 27952 37020 28016 37024
rect 27952 36964 27956 37020
rect 27956 36964 28012 37020
rect 28012 36964 28016 37020
rect 27952 36960 28016 36964
rect 28032 37020 28096 37024
rect 28032 36964 28036 37020
rect 28036 36964 28092 37020
rect 28092 36964 28096 37020
rect 28032 36960 28096 36964
rect 28112 37020 28176 37024
rect 28112 36964 28116 37020
rect 28116 36964 28172 37020
rect 28172 36964 28176 37020
rect 28112 36960 28176 36964
rect 28192 37020 28256 37024
rect 28192 36964 28196 37020
rect 28196 36964 28252 37020
rect 28252 36964 28256 37020
rect 28192 36960 28256 36964
rect 37952 37020 38016 37024
rect 37952 36964 37956 37020
rect 37956 36964 38012 37020
rect 38012 36964 38016 37020
rect 37952 36960 38016 36964
rect 38032 37020 38096 37024
rect 38032 36964 38036 37020
rect 38036 36964 38092 37020
rect 38092 36964 38096 37020
rect 38032 36960 38096 36964
rect 38112 37020 38176 37024
rect 38112 36964 38116 37020
rect 38116 36964 38172 37020
rect 38172 36964 38176 37020
rect 38112 36960 38176 36964
rect 38192 37020 38256 37024
rect 38192 36964 38196 37020
rect 38196 36964 38252 37020
rect 38252 36964 38256 37020
rect 38192 36960 38256 36964
rect 47952 37020 48016 37024
rect 47952 36964 47956 37020
rect 47956 36964 48012 37020
rect 48012 36964 48016 37020
rect 47952 36960 48016 36964
rect 48032 37020 48096 37024
rect 48032 36964 48036 37020
rect 48036 36964 48092 37020
rect 48092 36964 48096 37020
rect 48032 36960 48096 36964
rect 48112 37020 48176 37024
rect 48112 36964 48116 37020
rect 48116 36964 48172 37020
rect 48172 36964 48176 37020
rect 48112 36960 48176 36964
rect 48192 37020 48256 37024
rect 48192 36964 48196 37020
rect 48196 36964 48252 37020
rect 48252 36964 48256 37020
rect 48192 36960 48256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 32952 36476 33016 36480
rect 32952 36420 32956 36476
rect 32956 36420 33012 36476
rect 33012 36420 33016 36476
rect 32952 36416 33016 36420
rect 33032 36476 33096 36480
rect 33032 36420 33036 36476
rect 33036 36420 33092 36476
rect 33092 36420 33096 36476
rect 33032 36416 33096 36420
rect 33112 36476 33176 36480
rect 33112 36420 33116 36476
rect 33116 36420 33172 36476
rect 33172 36420 33176 36476
rect 33112 36416 33176 36420
rect 33192 36476 33256 36480
rect 33192 36420 33196 36476
rect 33196 36420 33252 36476
rect 33252 36420 33256 36476
rect 33192 36416 33256 36420
rect 42952 36476 43016 36480
rect 42952 36420 42956 36476
rect 42956 36420 43012 36476
rect 43012 36420 43016 36476
rect 42952 36416 43016 36420
rect 43032 36476 43096 36480
rect 43032 36420 43036 36476
rect 43036 36420 43092 36476
rect 43092 36420 43096 36476
rect 43032 36416 43096 36420
rect 43112 36476 43176 36480
rect 43112 36420 43116 36476
rect 43116 36420 43172 36476
rect 43172 36420 43176 36476
rect 43112 36416 43176 36420
rect 43192 36476 43256 36480
rect 43192 36420 43196 36476
rect 43196 36420 43252 36476
rect 43252 36420 43256 36476
rect 43192 36416 43256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 27952 35932 28016 35936
rect 27952 35876 27956 35932
rect 27956 35876 28012 35932
rect 28012 35876 28016 35932
rect 27952 35872 28016 35876
rect 28032 35932 28096 35936
rect 28032 35876 28036 35932
rect 28036 35876 28092 35932
rect 28092 35876 28096 35932
rect 28032 35872 28096 35876
rect 28112 35932 28176 35936
rect 28112 35876 28116 35932
rect 28116 35876 28172 35932
rect 28172 35876 28176 35932
rect 28112 35872 28176 35876
rect 28192 35932 28256 35936
rect 28192 35876 28196 35932
rect 28196 35876 28252 35932
rect 28252 35876 28256 35932
rect 28192 35872 28256 35876
rect 37952 35932 38016 35936
rect 37952 35876 37956 35932
rect 37956 35876 38012 35932
rect 38012 35876 38016 35932
rect 37952 35872 38016 35876
rect 38032 35932 38096 35936
rect 38032 35876 38036 35932
rect 38036 35876 38092 35932
rect 38092 35876 38096 35932
rect 38032 35872 38096 35876
rect 38112 35932 38176 35936
rect 38112 35876 38116 35932
rect 38116 35876 38172 35932
rect 38172 35876 38176 35932
rect 38112 35872 38176 35876
rect 38192 35932 38256 35936
rect 38192 35876 38196 35932
rect 38196 35876 38252 35932
rect 38252 35876 38256 35932
rect 38192 35872 38256 35876
rect 47952 35932 48016 35936
rect 47952 35876 47956 35932
rect 47956 35876 48012 35932
rect 48012 35876 48016 35932
rect 47952 35872 48016 35876
rect 48032 35932 48096 35936
rect 48032 35876 48036 35932
rect 48036 35876 48092 35932
rect 48092 35876 48096 35932
rect 48032 35872 48096 35876
rect 48112 35932 48176 35936
rect 48112 35876 48116 35932
rect 48116 35876 48172 35932
rect 48172 35876 48176 35932
rect 48112 35872 48176 35876
rect 48192 35932 48256 35936
rect 48192 35876 48196 35932
rect 48196 35876 48252 35932
rect 48252 35876 48256 35932
rect 48192 35872 48256 35876
rect 28396 35668 28460 35732
rect 38332 35728 38396 35732
rect 38332 35672 38382 35728
rect 38382 35672 38396 35728
rect 38332 35668 38396 35672
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 32952 35388 33016 35392
rect 32952 35332 32956 35388
rect 32956 35332 33012 35388
rect 33012 35332 33016 35388
rect 32952 35328 33016 35332
rect 33032 35388 33096 35392
rect 33032 35332 33036 35388
rect 33036 35332 33092 35388
rect 33092 35332 33096 35388
rect 33032 35328 33096 35332
rect 33112 35388 33176 35392
rect 33112 35332 33116 35388
rect 33116 35332 33172 35388
rect 33172 35332 33176 35388
rect 33112 35328 33176 35332
rect 33192 35388 33256 35392
rect 33192 35332 33196 35388
rect 33196 35332 33252 35388
rect 33252 35332 33256 35388
rect 33192 35328 33256 35332
rect 42952 35388 43016 35392
rect 42952 35332 42956 35388
rect 42956 35332 43012 35388
rect 43012 35332 43016 35388
rect 42952 35328 43016 35332
rect 43032 35388 43096 35392
rect 43032 35332 43036 35388
rect 43036 35332 43092 35388
rect 43092 35332 43096 35388
rect 43032 35328 43096 35332
rect 43112 35388 43176 35392
rect 43112 35332 43116 35388
rect 43116 35332 43172 35388
rect 43172 35332 43176 35388
rect 43112 35328 43176 35332
rect 43192 35388 43256 35392
rect 43192 35332 43196 35388
rect 43196 35332 43252 35388
rect 43252 35332 43256 35388
rect 43192 35328 43256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 27952 34844 28016 34848
rect 27952 34788 27956 34844
rect 27956 34788 28012 34844
rect 28012 34788 28016 34844
rect 27952 34784 28016 34788
rect 28032 34844 28096 34848
rect 28032 34788 28036 34844
rect 28036 34788 28092 34844
rect 28092 34788 28096 34844
rect 28032 34784 28096 34788
rect 28112 34844 28176 34848
rect 28112 34788 28116 34844
rect 28116 34788 28172 34844
rect 28172 34788 28176 34844
rect 28112 34784 28176 34788
rect 28192 34844 28256 34848
rect 28192 34788 28196 34844
rect 28196 34788 28252 34844
rect 28252 34788 28256 34844
rect 28192 34784 28256 34788
rect 37952 34844 38016 34848
rect 37952 34788 37956 34844
rect 37956 34788 38012 34844
rect 38012 34788 38016 34844
rect 37952 34784 38016 34788
rect 38032 34844 38096 34848
rect 38032 34788 38036 34844
rect 38036 34788 38092 34844
rect 38092 34788 38096 34844
rect 38032 34784 38096 34788
rect 38112 34844 38176 34848
rect 38112 34788 38116 34844
rect 38116 34788 38172 34844
rect 38172 34788 38176 34844
rect 38112 34784 38176 34788
rect 38192 34844 38256 34848
rect 38192 34788 38196 34844
rect 38196 34788 38252 34844
rect 38252 34788 38256 34844
rect 38192 34784 38256 34788
rect 47952 34844 48016 34848
rect 47952 34788 47956 34844
rect 47956 34788 48012 34844
rect 48012 34788 48016 34844
rect 47952 34784 48016 34788
rect 48032 34844 48096 34848
rect 48032 34788 48036 34844
rect 48036 34788 48092 34844
rect 48092 34788 48096 34844
rect 48032 34784 48096 34788
rect 48112 34844 48176 34848
rect 48112 34788 48116 34844
rect 48116 34788 48172 34844
rect 48172 34788 48176 34844
rect 48112 34784 48176 34788
rect 48192 34844 48256 34848
rect 48192 34788 48196 34844
rect 48196 34788 48252 34844
rect 48252 34788 48256 34844
rect 48192 34784 48256 34788
rect 28580 34580 28644 34644
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 32952 34300 33016 34304
rect 32952 34244 32956 34300
rect 32956 34244 33012 34300
rect 33012 34244 33016 34300
rect 32952 34240 33016 34244
rect 33032 34300 33096 34304
rect 33032 34244 33036 34300
rect 33036 34244 33092 34300
rect 33092 34244 33096 34300
rect 33032 34240 33096 34244
rect 33112 34300 33176 34304
rect 33112 34244 33116 34300
rect 33116 34244 33172 34300
rect 33172 34244 33176 34300
rect 33112 34240 33176 34244
rect 33192 34300 33256 34304
rect 33192 34244 33196 34300
rect 33196 34244 33252 34300
rect 33252 34244 33256 34300
rect 33192 34240 33256 34244
rect 42952 34300 43016 34304
rect 42952 34244 42956 34300
rect 42956 34244 43012 34300
rect 43012 34244 43016 34300
rect 42952 34240 43016 34244
rect 43032 34300 43096 34304
rect 43032 34244 43036 34300
rect 43036 34244 43092 34300
rect 43092 34244 43096 34300
rect 43032 34240 43096 34244
rect 43112 34300 43176 34304
rect 43112 34244 43116 34300
rect 43116 34244 43172 34300
rect 43172 34244 43176 34300
rect 43112 34240 43176 34244
rect 43192 34300 43256 34304
rect 43192 34244 43196 34300
rect 43196 34244 43252 34300
rect 43252 34244 43256 34300
rect 43192 34240 43256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 27952 33756 28016 33760
rect 27952 33700 27956 33756
rect 27956 33700 28012 33756
rect 28012 33700 28016 33756
rect 27952 33696 28016 33700
rect 28032 33756 28096 33760
rect 28032 33700 28036 33756
rect 28036 33700 28092 33756
rect 28092 33700 28096 33756
rect 28032 33696 28096 33700
rect 28112 33756 28176 33760
rect 28112 33700 28116 33756
rect 28116 33700 28172 33756
rect 28172 33700 28176 33756
rect 28112 33696 28176 33700
rect 28192 33756 28256 33760
rect 28192 33700 28196 33756
rect 28196 33700 28252 33756
rect 28252 33700 28256 33756
rect 28192 33696 28256 33700
rect 37952 33756 38016 33760
rect 37952 33700 37956 33756
rect 37956 33700 38012 33756
rect 38012 33700 38016 33756
rect 37952 33696 38016 33700
rect 38032 33756 38096 33760
rect 38032 33700 38036 33756
rect 38036 33700 38092 33756
rect 38092 33700 38096 33756
rect 38032 33696 38096 33700
rect 38112 33756 38176 33760
rect 38112 33700 38116 33756
rect 38116 33700 38172 33756
rect 38172 33700 38176 33756
rect 38112 33696 38176 33700
rect 38192 33756 38256 33760
rect 38192 33700 38196 33756
rect 38196 33700 38252 33756
rect 38252 33700 38256 33756
rect 38192 33696 38256 33700
rect 47952 33756 48016 33760
rect 47952 33700 47956 33756
rect 47956 33700 48012 33756
rect 48012 33700 48016 33756
rect 47952 33696 48016 33700
rect 48032 33756 48096 33760
rect 48032 33700 48036 33756
rect 48036 33700 48092 33756
rect 48092 33700 48096 33756
rect 48032 33696 48096 33700
rect 48112 33756 48176 33760
rect 48112 33700 48116 33756
rect 48116 33700 48172 33756
rect 48172 33700 48176 33756
rect 48112 33696 48176 33700
rect 48192 33756 48256 33760
rect 48192 33700 48196 33756
rect 48196 33700 48252 33756
rect 48252 33700 48256 33756
rect 48192 33696 48256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 32952 33212 33016 33216
rect 32952 33156 32956 33212
rect 32956 33156 33012 33212
rect 33012 33156 33016 33212
rect 32952 33152 33016 33156
rect 33032 33212 33096 33216
rect 33032 33156 33036 33212
rect 33036 33156 33092 33212
rect 33092 33156 33096 33212
rect 33032 33152 33096 33156
rect 33112 33212 33176 33216
rect 33112 33156 33116 33212
rect 33116 33156 33172 33212
rect 33172 33156 33176 33212
rect 33112 33152 33176 33156
rect 33192 33212 33256 33216
rect 33192 33156 33196 33212
rect 33196 33156 33252 33212
rect 33252 33156 33256 33212
rect 33192 33152 33256 33156
rect 42952 33212 43016 33216
rect 42952 33156 42956 33212
rect 42956 33156 43012 33212
rect 43012 33156 43016 33212
rect 42952 33152 43016 33156
rect 43032 33212 43096 33216
rect 43032 33156 43036 33212
rect 43036 33156 43092 33212
rect 43092 33156 43096 33212
rect 43032 33152 43096 33156
rect 43112 33212 43176 33216
rect 43112 33156 43116 33212
rect 43116 33156 43172 33212
rect 43172 33156 43176 33212
rect 43112 33152 43176 33156
rect 43192 33212 43256 33216
rect 43192 33156 43196 33212
rect 43196 33156 43252 33212
rect 43252 33156 43256 33212
rect 43192 33152 43256 33156
rect 35388 32948 35452 33012
rect 27108 32812 27172 32876
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 27952 32668 28016 32672
rect 27952 32612 27956 32668
rect 27956 32612 28012 32668
rect 28012 32612 28016 32668
rect 27952 32608 28016 32612
rect 28032 32668 28096 32672
rect 28032 32612 28036 32668
rect 28036 32612 28092 32668
rect 28092 32612 28096 32668
rect 28032 32608 28096 32612
rect 28112 32668 28176 32672
rect 28112 32612 28116 32668
rect 28116 32612 28172 32668
rect 28172 32612 28176 32668
rect 28112 32608 28176 32612
rect 28192 32668 28256 32672
rect 28192 32612 28196 32668
rect 28196 32612 28252 32668
rect 28252 32612 28256 32668
rect 28192 32608 28256 32612
rect 37952 32668 38016 32672
rect 37952 32612 37956 32668
rect 37956 32612 38012 32668
rect 38012 32612 38016 32668
rect 37952 32608 38016 32612
rect 38032 32668 38096 32672
rect 38032 32612 38036 32668
rect 38036 32612 38092 32668
rect 38092 32612 38096 32668
rect 38032 32608 38096 32612
rect 38112 32668 38176 32672
rect 38112 32612 38116 32668
rect 38116 32612 38172 32668
rect 38172 32612 38176 32668
rect 38112 32608 38176 32612
rect 38192 32668 38256 32672
rect 38192 32612 38196 32668
rect 38196 32612 38252 32668
rect 38252 32612 38256 32668
rect 38192 32608 38256 32612
rect 47952 32668 48016 32672
rect 47952 32612 47956 32668
rect 47956 32612 48012 32668
rect 48012 32612 48016 32668
rect 47952 32608 48016 32612
rect 48032 32668 48096 32672
rect 48032 32612 48036 32668
rect 48036 32612 48092 32668
rect 48092 32612 48096 32668
rect 48032 32608 48096 32612
rect 48112 32668 48176 32672
rect 48112 32612 48116 32668
rect 48116 32612 48172 32668
rect 48172 32612 48176 32668
rect 48112 32608 48176 32612
rect 48192 32668 48256 32672
rect 48192 32612 48196 32668
rect 48196 32612 48252 32668
rect 48252 32612 48256 32668
rect 48192 32608 48256 32612
rect 38332 32464 38396 32468
rect 38332 32408 38346 32464
rect 38346 32408 38396 32464
rect 38332 32404 38396 32408
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 32952 32124 33016 32128
rect 32952 32068 32956 32124
rect 32956 32068 33012 32124
rect 33012 32068 33016 32124
rect 32952 32064 33016 32068
rect 33032 32124 33096 32128
rect 33032 32068 33036 32124
rect 33036 32068 33092 32124
rect 33092 32068 33096 32124
rect 33032 32064 33096 32068
rect 33112 32124 33176 32128
rect 33112 32068 33116 32124
rect 33116 32068 33172 32124
rect 33172 32068 33176 32124
rect 33112 32064 33176 32068
rect 33192 32124 33256 32128
rect 33192 32068 33196 32124
rect 33196 32068 33252 32124
rect 33252 32068 33256 32124
rect 33192 32064 33256 32068
rect 42952 32124 43016 32128
rect 42952 32068 42956 32124
rect 42956 32068 43012 32124
rect 43012 32068 43016 32124
rect 42952 32064 43016 32068
rect 43032 32124 43096 32128
rect 43032 32068 43036 32124
rect 43036 32068 43092 32124
rect 43092 32068 43096 32124
rect 43032 32064 43096 32068
rect 43112 32124 43176 32128
rect 43112 32068 43116 32124
rect 43116 32068 43172 32124
rect 43172 32068 43176 32124
rect 43112 32064 43176 32068
rect 43192 32124 43256 32128
rect 43192 32068 43196 32124
rect 43196 32068 43252 32124
rect 43252 32068 43256 32124
rect 43192 32064 43256 32068
rect 38516 31724 38580 31788
rect 28396 31588 28460 31652
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 27952 31580 28016 31584
rect 27952 31524 27956 31580
rect 27956 31524 28012 31580
rect 28012 31524 28016 31580
rect 27952 31520 28016 31524
rect 28032 31580 28096 31584
rect 28032 31524 28036 31580
rect 28036 31524 28092 31580
rect 28092 31524 28096 31580
rect 28032 31520 28096 31524
rect 28112 31580 28176 31584
rect 28112 31524 28116 31580
rect 28116 31524 28172 31580
rect 28172 31524 28176 31580
rect 28112 31520 28176 31524
rect 28192 31580 28256 31584
rect 28192 31524 28196 31580
rect 28196 31524 28252 31580
rect 28252 31524 28256 31580
rect 28192 31520 28256 31524
rect 37952 31580 38016 31584
rect 37952 31524 37956 31580
rect 37956 31524 38012 31580
rect 38012 31524 38016 31580
rect 37952 31520 38016 31524
rect 38032 31580 38096 31584
rect 38032 31524 38036 31580
rect 38036 31524 38092 31580
rect 38092 31524 38096 31580
rect 38032 31520 38096 31524
rect 38112 31580 38176 31584
rect 38112 31524 38116 31580
rect 38116 31524 38172 31580
rect 38172 31524 38176 31580
rect 38112 31520 38176 31524
rect 38192 31580 38256 31584
rect 38192 31524 38196 31580
rect 38196 31524 38252 31580
rect 38252 31524 38256 31580
rect 38192 31520 38256 31524
rect 47952 31580 48016 31584
rect 47952 31524 47956 31580
rect 47956 31524 48012 31580
rect 48012 31524 48016 31580
rect 47952 31520 48016 31524
rect 48032 31580 48096 31584
rect 48032 31524 48036 31580
rect 48036 31524 48092 31580
rect 48092 31524 48096 31580
rect 48032 31520 48096 31524
rect 48112 31580 48176 31584
rect 48112 31524 48116 31580
rect 48116 31524 48172 31580
rect 48172 31524 48176 31580
rect 48112 31520 48176 31524
rect 48192 31580 48256 31584
rect 48192 31524 48196 31580
rect 48196 31524 48252 31580
rect 48252 31524 48256 31580
rect 48192 31520 48256 31524
rect 28580 31452 28644 31516
rect 22692 31180 22756 31244
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 32952 31036 33016 31040
rect 32952 30980 32956 31036
rect 32956 30980 33012 31036
rect 33012 30980 33016 31036
rect 32952 30976 33016 30980
rect 33032 31036 33096 31040
rect 33032 30980 33036 31036
rect 33036 30980 33092 31036
rect 33092 30980 33096 31036
rect 33032 30976 33096 30980
rect 33112 31036 33176 31040
rect 33112 30980 33116 31036
rect 33116 30980 33172 31036
rect 33172 30980 33176 31036
rect 33112 30976 33176 30980
rect 33192 31036 33256 31040
rect 33192 30980 33196 31036
rect 33196 30980 33252 31036
rect 33252 30980 33256 31036
rect 33192 30976 33256 30980
rect 42952 31036 43016 31040
rect 42952 30980 42956 31036
rect 42956 30980 43012 31036
rect 43012 30980 43016 31036
rect 42952 30976 43016 30980
rect 43032 31036 43096 31040
rect 43032 30980 43036 31036
rect 43036 30980 43092 31036
rect 43092 30980 43096 31036
rect 43032 30976 43096 30980
rect 43112 31036 43176 31040
rect 43112 30980 43116 31036
rect 43116 30980 43172 31036
rect 43172 30980 43176 31036
rect 43112 30976 43176 30980
rect 43192 31036 43256 31040
rect 43192 30980 43196 31036
rect 43196 30980 43252 31036
rect 43252 30980 43256 31036
rect 43192 30976 43256 30980
rect 36676 30908 36740 30972
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 27952 30492 28016 30496
rect 27952 30436 27956 30492
rect 27956 30436 28012 30492
rect 28012 30436 28016 30492
rect 27952 30432 28016 30436
rect 28032 30492 28096 30496
rect 28032 30436 28036 30492
rect 28036 30436 28092 30492
rect 28092 30436 28096 30492
rect 28032 30432 28096 30436
rect 28112 30492 28176 30496
rect 28112 30436 28116 30492
rect 28116 30436 28172 30492
rect 28172 30436 28176 30492
rect 28112 30432 28176 30436
rect 28192 30492 28256 30496
rect 28192 30436 28196 30492
rect 28196 30436 28252 30492
rect 28252 30436 28256 30492
rect 28192 30432 28256 30436
rect 37952 30492 38016 30496
rect 37952 30436 37956 30492
rect 37956 30436 38012 30492
rect 38012 30436 38016 30492
rect 37952 30432 38016 30436
rect 38032 30492 38096 30496
rect 38032 30436 38036 30492
rect 38036 30436 38092 30492
rect 38092 30436 38096 30492
rect 38032 30432 38096 30436
rect 38112 30492 38176 30496
rect 38112 30436 38116 30492
rect 38116 30436 38172 30492
rect 38172 30436 38176 30492
rect 38112 30432 38176 30436
rect 38192 30492 38256 30496
rect 38192 30436 38196 30492
rect 38196 30436 38252 30492
rect 38252 30436 38256 30492
rect 38192 30432 38256 30436
rect 47952 30492 48016 30496
rect 47952 30436 47956 30492
rect 47956 30436 48012 30492
rect 48012 30436 48016 30492
rect 47952 30432 48016 30436
rect 48032 30492 48096 30496
rect 48032 30436 48036 30492
rect 48036 30436 48092 30492
rect 48092 30436 48096 30492
rect 48032 30432 48096 30436
rect 48112 30492 48176 30496
rect 48112 30436 48116 30492
rect 48116 30436 48172 30492
rect 48172 30436 48176 30492
rect 48112 30432 48176 30436
rect 48192 30492 48256 30496
rect 48192 30436 48196 30492
rect 48196 30436 48252 30492
rect 48252 30436 48256 30492
rect 48192 30432 48256 30436
rect 37228 30364 37292 30428
rect 35940 30228 36004 30292
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 32952 29948 33016 29952
rect 32952 29892 32956 29948
rect 32956 29892 33012 29948
rect 33012 29892 33016 29948
rect 32952 29888 33016 29892
rect 33032 29948 33096 29952
rect 33032 29892 33036 29948
rect 33036 29892 33092 29948
rect 33092 29892 33096 29948
rect 33032 29888 33096 29892
rect 33112 29948 33176 29952
rect 33112 29892 33116 29948
rect 33116 29892 33172 29948
rect 33172 29892 33176 29948
rect 33112 29888 33176 29892
rect 33192 29948 33256 29952
rect 33192 29892 33196 29948
rect 33196 29892 33252 29948
rect 33252 29892 33256 29948
rect 33192 29888 33256 29892
rect 42952 29948 43016 29952
rect 42952 29892 42956 29948
rect 42956 29892 43012 29948
rect 43012 29892 43016 29948
rect 42952 29888 43016 29892
rect 43032 29948 43096 29952
rect 43032 29892 43036 29948
rect 43036 29892 43092 29948
rect 43092 29892 43096 29948
rect 43032 29888 43096 29892
rect 43112 29948 43176 29952
rect 43112 29892 43116 29948
rect 43116 29892 43172 29948
rect 43172 29892 43176 29948
rect 43112 29888 43176 29892
rect 43192 29948 43256 29952
rect 43192 29892 43196 29948
rect 43196 29892 43252 29948
rect 43252 29892 43256 29948
rect 43192 29888 43256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 27952 29404 28016 29408
rect 27952 29348 27956 29404
rect 27956 29348 28012 29404
rect 28012 29348 28016 29404
rect 27952 29344 28016 29348
rect 28032 29404 28096 29408
rect 28032 29348 28036 29404
rect 28036 29348 28092 29404
rect 28092 29348 28096 29404
rect 28032 29344 28096 29348
rect 28112 29404 28176 29408
rect 28112 29348 28116 29404
rect 28116 29348 28172 29404
rect 28172 29348 28176 29404
rect 28112 29344 28176 29348
rect 28192 29404 28256 29408
rect 28192 29348 28196 29404
rect 28196 29348 28252 29404
rect 28252 29348 28256 29404
rect 28192 29344 28256 29348
rect 37952 29404 38016 29408
rect 37952 29348 37956 29404
rect 37956 29348 38012 29404
rect 38012 29348 38016 29404
rect 37952 29344 38016 29348
rect 38032 29404 38096 29408
rect 38032 29348 38036 29404
rect 38036 29348 38092 29404
rect 38092 29348 38096 29404
rect 38032 29344 38096 29348
rect 38112 29404 38176 29408
rect 38112 29348 38116 29404
rect 38116 29348 38172 29404
rect 38172 29348 38176 29404
rect 38112 29344 38176 29348
rect 38192 29404 38256 29408
rect 38192 29348 38196 29404
rect 38196 29348 38252 29404
rect 38252 29348 38256 29404
rect 38192 29344 38256 29348
rect 47952 29404 48016 29408
rect 47952 29348 47956 29404
rect 47956 29348 48012 29404
rect 48012 29348 48016 29404
rect 47952 29344 48016 29348
rect 48032 29404 48096 29408
rect 48032 29348 48036 29404
rect 48036 29348 48092 29404
rect 48092 29348 48096 29404
rect 48032 29344 48096 29348
rect 48112 29404 48176 29408
rect 48112 29348 48116 29404
rect 48116 29348 48172 29404
rect 48172 29348 48176 29404
rect 48112 29344 48176 29348
rect 48192 29404 48256 29408
rect 48192 29348 48196 29404
rect 48196 29348 48252 29404
rect 48252 29348 48256 29404
rect 48192 29344 48256 29348
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 32952 28860 33016 28864
rect 32952 28804 32956 28860
rect 32956 28804 33012 28860
rect 33012 28804 33016 28860
rect 32952 28800 33016 28804
rect 33032 28860 33096 28864
rect 33032 28804 33036 28860
rect 33036 28804 33092 28860
rect 33092 28804 33096 28860
rect 33032 28800 33096 28804
rect 33112 28860 33176 28864
rect 33112 28804 33116 28860
rect 33116 28804 33172 28860
rect 33172 28804 33176 28860
rect 33112 28800 33176 28804
rect 33192 28860 33256 28864
rect 33192 28804 33196 28860
rect 33196 28804 33252 28860
rect 33252 28804 33256 28860
rect 33192 28800 33256 28804
rect 42952 28860 43016 28864
rect 42952 28804 42956 28860
rect 42956 28804 43012 28860
rect 43012 28804 43016 28860
rect 42952 28800 43016 28804
rect 43032 28860 43096 28864
rect 43032 28804 43036 28860
rect 43036 28804 43092 28860
rect 43092 28804 43096 28860
rect 43032 28800 43096 28804
rect 43112 28860 43176 28864
rect 43112 28804 43116 28860
rect 43116 28804 43172 28860
rect 43172 28804 43176 28860
rect 43112 28800 43176 28804
rect 43192 28860 43256 28864
rect 43192 28804 43196 28860
rect 43196 28804 43252 28860
rect 43252 28804 43256 28860
rect 43192 28800 43256 28804
rect 40540 28460 40604 28524
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 27952 28316 28016 28320
rect 27952 28260 27956 28316
rect 27956 28260 28012 28316
rect 28012 28260 28016 28316
rect 27952 28256 28016 28260
rect 28032 28316 28096 28320
rect 28032 28260 28036 28316
rect 28036 28260 28092 28316
rect 28092 28260 28096 28316
rect 28032 28256 28096 28260
rect 28112 28316 28176 28320
rect 28112 28260 28116 28316
rect 28116 28260 28172 28316
rect 28172 28260 28176 28316
rect 28112 28256 28176 28260
rect 28192 28316 28256 28320
rect 28192 28260 28196 28316
rect 28196 28260 28252 28316
rect 28252 28260 28256 28316
rect 28192 28256 28256 28260
rect 37952 28316 38016 28320
rect 37952 28260 37956 28316
rect 37956 28260 38012 28316
rect 38012 28260 38016 28316
rect 37952 28256 38016 28260
rect 38032 28316 38096 28320
rect 38032 28260 38036 28316
rect 38036 28260 38092 28316
rect 38092 28260 38096 28316
rect 38032 28256 38096 28260
rect 38112 28316 38176 28320
rect 38112 28260 38116 28316
rect 38116 28260 38172 28316
rect 38172 28260 38176 28316
rect 38112 28256 38176 28260
rect 38192 28316 38256 28320
rect 38192 28260 38196 28316
rect 38196 28260 38252 28316
rect 38252 28260 38256 28316
rect 38192 28256 38256 28260
rect 47952 28316 48016 28320
rect 47952 28260 47956 28316
rect 47956 28260 48012 28316
rect 48012 28260 48016 28316
rect 47952 28256 48016 28260
rect 48032 28316 48096 28320
rect 48032 28260 48036 28316
rect 48036 28260 48092 28316
rect 48092 28260 48096 28316
rect 48032 28256 48096 28260
rect 48112 28316 48176 28320
rect 48112 28260 48116 28316
rect 48116 28260 48172 28316
rect 48172 28260 48176 28316
rect 48112 28256 48176 28260
rect 48192 28316 48256 28320
rect 48192 28260 48196 28316
rect 48196 28260 48252 28316
rect 48252 28260 48256 28316
rect 48192 28256 48256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 32952 27772 33016 27776
rect 32952 27716 32956 27772
rect 32956 27716 33012 27772
rect 33012 27716 33016 27772
rect 32952 27712 33016 27716
rect 33032 27772 33096 27776
rect 33032 27716 33036 27772
rect 33036 27716 33092 27772
rect 33092 27716 33096 27772
rect 33032 27712 33096 27716
rect 33112 27772 33176 27776
rect 33112 27716 33116 27772
rect 33116 27716 33172 27772
rect 33172 27716 33176 27772
rect 33112 27712 33176 27716
rect 33192 27772 33256 27776
rect 33192 27716 33196 27772
rect 33196 27716 33252 27772
rect 33252 27716 33256 27772
rect 33192 27712 33256 27716
rect 42952 27772 43016 27776
rect 42952 27716 42956 27772
rect 42956 27716 43012 27772
rect 43012 27716 43016 27772
rect 42952 27712 43016 27716
rect 43032 27772 43096 27776
rect 43032 27716 43036 27772
rect 43036 27716 43092 27772
rect 43092 27716 43096 27772
rect 43032 27712 43096 27716
rect 43112 27772 43176 27776
rect 43112 27716 43116 27772
rect 43116 27716 43172 27772
rect 43172 27716 43176 27772
rect 43112 27712 43176 27716
rect 43192 27772 43256 27776
rect 43192 27716 43196 27772
rect 43196 27716 43252 27772
rect 43252 27716 43256 27772
rect 43192 27712 43256 27716
rect 38516 27372 38580 27436
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 27952 27228 28016 27232
rect 27952 27172 27956 27228
rect 27956 27172 28012 27228
rect 28012 27172 28016 27228
rect 27952 27168 28016 27172
rect 28032 27228 28096 27232
rect 28032 27172 28036 27228
rect 28036 27172 28092 27228
rect 28092 27172 28096 27228
rect 28032 27168 28096 27172
rect 28112 27228 28176 27232
rect 28112 27172 28116 27228
rect 28116 27172 28172 27228
rect 28172 27172 28176 27228
rect 28112 27168 28176 27172
rect 28192 27228 28256 27232
rect 28192 27172 28196 27228
rect 28196 27172 28252 27228
rect 28252 27172 28256 27228
rect 28192 27168 28256 27172
rect 37952 27228 38016 27232
rect 37952 27172 37956 27228
rect 37956 27172 38012 27228
rect 38012 27172 38016 27228
rect 37952 27168 38016 27172
rect 38032 27228 38096 27232
rect 38032 27172 38036 27228
rect 38036 27172 38092 27228
rect 38092 27172 38096 27228
rect 38032 27168 38096 27172
rect 38112 27228 38176 27232
rect 38112 27172 38116 27228
rect 38116 27172 38172 27228
rect 38172 27172 38176 27228
rect 38112 27168 38176 27172
rect 38192 27228 38256 27232
rect 38192 27172 38196 27228
rect 38196 27172 38252 27228
rect 38252 27172 38256 27228
rect 38192 27168 38256 27172
rect 47952 27228 48016 27232
rect 47952 27172 47956 27228
rect 47956 27172 48012 27228
rect 48012 27172 48016 27228
rect 47952 27168 48016 27172
rect 48032 27228 48096 27232
rect 48032 27172 48036 27228
rect 48036 27172 48092 27228
rect 48092 27172 48096 27228
rect 48032 27168 48096 27172
rect 48112 27228 48176 27232
rect 48112 27172 48116 27228
rect 48116 27172 48172 27228
rect 48172 27172 48176 27228
rect 48112 27168 48176 27172
rect 48192 27228 48256 27232
rect 48192 27172 48196 27228
rect 48196 27172 48252 27228
rect 48252 27172 48256 27228
rect 48192 27168 48256 27172
rect 39988 26964 40052 27028
rect 30604 26828 30668 26892
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 32952 26684 33016 26688
rect 32952 26628 32956 26684
rect 32956 26628 33012 26684
rect 33012 26628 33016 26684
rect 32952 26624 33016 26628
rect 33032 26684 33096 26688
rect 33032 26628 33036 26684
rect 33036 26628 33092 26684
rect 33092 26628 33096 26684
rect 33032 26624 33096 26628
rect 33112 26684 33176 26688
rect 33112 26628 33116 26684
rect 33116 26628 33172 26684
rect 33172 26628 33176 26684
rect 33112 26624 33176 26628
rect 33192 26684 33256 26688
rect 33192 26628 33196 26684
rect 33196 26628 33252 26684
rect 33252 26628 33256 26684
rect 33192 26624 33256 26628
rect 42952 26684 43016 26688
rect 42952 26628 42956 26684
rect 42956 26628 43012 26684
rect 43012 26628 43016 26684
rect 42952 26624 43016 26628
rect 43032 26684 43096 26688
rect 43032 26628 43036 26684
rect 43036 26628 43092 26684
rect 43092 26628 43096 26684
rect 43032 26624 43096 26628
rect 43112 26684 43176 26688
rect 43112 26628 43116 26684
rect 43116 26628 43172 26684
rect 43172 26628 43176 26684
rect 43112 26624 43176 26628
rect 43192 26684 43256 26688
rect 43192 26628 43196 26684
rect 43196 26628 43252 26684
rect 43252 26628 43256 26684
rect 43192 26624 43256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 27952 26140 28016 26144
rect 27952 26084 27956 26140
rect 27956 26084 28012 26140
rect 28012 26084 28016 26140
rect 27952 26080 28016 26084
rect 28032 26140 28096 26144
rect 28032 26084 28036 26140
rect 28036 26084 28092 26140
rect 28092 26084 28096 26140
rect 28032 26080 28096 26084
rect 28112 26140 28176 26144
rect 28112 26084 28116 26140
rect 28116 26084 28172 26140
rect 28172 26084 28176 26140
rect 28112 26080 28176 26084
rect 28192 26140 28256 26144
rect 28192 26084 28196 26140
rect 28196 26084 28252 26140
rect 28252 26084 28256 26140
rect 28192 26080 28256 26084
rect 37952 26140 38016 26144
rect 37952 26084 37956 26140
rect 37956 26084 38012 26140
rect 38012 26084 38016 26140
rect 37952 26080 38016 26084
rect 38032 26140 38096 26144
rect 38032 26084 38036 26140
rect 38036 26084 38092 26140
rect 38092 26084 38096 26140
rect 38032 26080 38096 26084
rect 38112 26140 38176 26144
rect 38112 26084 38116 26140
rect 38116 26084 38172 26140
rect 38172 26084 38176 26140
rect 38112 26080 38176 26084
rect 38192 26140 38256 26144
rect 38192 26084 38196 26140
rect 38196 26084 38252 26140
rect 38252 26084 38256 26140
rect 38192 26080 38256 26084
rect 47952 26140 48016 26144
rect 47952 26084 47956 26140
rect 47956 26084 48012 26140
rect 48012 26084 48016 26140
rect 47952 26080 48016 26084
rect 48032 26140 48096 26144
rect 48032 26084 48036 26140
rect 48036 26084 48092 26140
rect 48092 26084 48096 26140
rect 48032 26080 48096 26084
rect 48112 26140 48176 26144
rect 48112 26084 48116 26140
rect 48116 26084 48172 26140
rect 48172 26084 48176 26140
rect 48112 26080 48176 26084
rect 48192 26140 48256 26144
rect 48192 26084 48196 26140
rect 48196 26084 48252 26140
rect 48252 26084 48256 26140
rect 48192 26080 48256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 32952 25596 33016 25600
rect 32952 25540 32956 25596
rect 32956 25540 33012 25596
rect 33012 25540 33016 25596
rect 32952 25536 33016 25540
rect 33032 25596 33096 25600
rect 33032 25540 33036 25596
rect 33036 25540 33092 25596
rect 33092 25540 33096 25596
rect 33032 25536 33096 25540
rect 33112 25596 33176 25600
rect 33112 25540 33116 25596
rect 33116 25540 33172 25596
rect 33172 25540 33176 25596
rect 33112 25536 33176 25540
rect 33192 25596 33256 25600
rect 33192 25540 33196 25596
rect 33196 25540 33252 25596
rect 33252 25540 33256 25596
rect 33192 25536 33256 25540
rect 42952 25596 43016 25600
rect 42952 25540 42956 25596
rect 42956 25540 43012 25596
rect 43012 25540 43016 25596
rect 42952 25536 43016 25540
rect 43032 25596 43096 25600
rect 43032 25540 43036 25596
rect 43036 25540 43092 25596
rect 43092 25540 43096 25596
rect 43032 25536 43096 25540
rect 43112 25596 43176 25600
rect 43112 25540 43116 25596
rect 43116 25540 43172 25596
rect 43172 25540 43176 25596
rect 43112 25536 43176 25540
rect 43192 25596 43256 25600
rect 43192 25540 43196 25596
rect 43196 25540 43252 25596
rect 43252 25540 43256 25596
rect 43192 25536 43256 25540
rect 30420 25196 30484 25260
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 27952 25052 28016 25056
rect 27952 24996 27956 25052
rect 27956 24996 28012 25052
rect 28012 24996 28016 25052
rect 27952 24992 28016 24996
rect 28032 25052 28096 25056
rect 28032 24996 28036 25052
rect 28036 24996 28092 25052
rect 28092 24996 28096 25052
rect 28032 24992 28096 24996
rect 28112 25052 28176 25056
rect 28112 24996 28116 25052
rect 28116 24996 28172 25052
rect 28172 24996 28176 25052
rect 28112 24992 28176 24996
rect 28192 25052 28256 25056
rect 28192 24996 28196 25052
rect 28196 24996 28252 25052
rect 28252 24996 28256 25052
rect 28192 24992 28256 24996
rect 37952 25052 38016 25056
rect 37952 24996 37956 25052
rect 37956 24996 38012 25052
rect 38012 24996 38016 25052
rect 37952 24992 38016 24996
rect 38032 25052 38096 25056
rect 38032 24996 38036 25052
rect 38036 24996 38092 25052
rect 38092 24996 38096 25052
rect 38032 24992 38096 24996
rect 38112 25052 38176 25056
rect 38112 24996 38116 25052
rect 38116 24996 38172 25052
rect 38172 24996 38176 25052
rect 38112 24992 38176 24996
rect 38192 25052 38256 25056
rect 38192 24996 38196 25052
rect 38196 24996 38252 25052
rect 38252 24996 38256 25052
rect 38192 24992 38256 24996
rect 47952 25052 48016 25056
rect 47952 24996 47956 25052
rect 47956 24996 48012 25052
rect 48012 24996 48016 25052
rect 47952 24992 48016 24996
rect 48032 25052 48096 25056
rect 48032 24996 48036 25052
rect 48036 24996 48092 25052
rect 48092 24996 48096 25052
rect 48032 24992 48096 24996
rect 48112 25052 48176 25056
rect 48112 24996 48116 25052
rect 48116 24996 48172 25052
rect 48172 24996 48176 25052
rect 48112 24992 48176 24996
rect 48192 25052 48256 25056
rect 48192 24996 48196 25052
rect 48196 24996 48252 25052
rect 48252 24996 48256 25052
rect 48192 24992 48256 24996
rect 26004 24712 26068 24716
rect 26004 24656 26018 24712
rect 26018 24656 26068 24712
rect 26004 24652 26068 24656
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 25636 24244 25700 24308
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 22692 22884 22756 22948
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 30420 20632 30484 20636
rect 30420 20576 30470 20632
rect 30470 20576 30484 20632
rect 30420 20572 30484 20576
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 26740 19212 26804 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 27108 18804 27172 18868
rect 27660 18728 27724 18732
rect 27660 18672 27710 18728
rect 27710 18672 27724 18728
rect 27660 18668 27724 18672
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 30604 17988 30668 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 27660 17096 27724 17100
rect 27660 17040 27710 17096
rect 27710 17040 27724 17096
rect 27660 17036 27724 17040
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 30604 12820 30668 12884
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 27108 3028 27172 3092
rect 22692 2892 22756 2956
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 27660 2484 27724 2548
rect 26004 2348 26068 2412
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
rect 26740 1940 26804 2004
rect 25636 1804 25700 1868
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 27944 54432 28264 54448
rect 27944 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28264 54432
rect 27944 53344 28264 54368
rect 27944 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28264 53344
rect 27944 52256 28264 53280
rect 27944 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28264 52256
rect 27944 51168 28264 52192
rect 27944 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28264 51168
rect 27944 50080 28264 51104
rect 27944 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28264 50080
rect 27944 48992 28264 50016
rect 27944 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28264 48992
rect 27944 47904 28264 48928
rect 27944 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28264 47904
rect 27944 46816 28264 47840
rect 27944 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28264 46816
rect 27944 45728 28264 46752
rect 27944 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28264 45728
rect 27944 44640 28264 45664
rect 27944 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28264 44640
rect 27944 43552 28264 44576
rect 27944 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28264 43552
rect 27944 42464 28264 43488
rect 27944 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28264 42464
rect 27944 41376 28264 42400
rect 27944 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28264 41376
rect 27944 40288 28264 41312
rect 27944 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28264 40288
rect 27944 39200 28264 40224
rect 27944 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28264 39200
rect 27944 38112 28264 39136
rect 27944 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28264 38112
rect 25635 37228 25701 37229
rect 25635 37164 25636 37228
rect 25700 37164 25701 37228
rect 25635 37163 25701 37164
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22691 31244 22757 31245
rect 22691 31180 22692 31244
rect 22756 31180 22757 31244
rect 22691 31179 22757 31180
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 22694 22949 22754 31179
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 25638 24309 25698 37163
rect 27944 37024 28264 38048
rect 27944 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28264 37024
rect 27944 35936 28264 36960
rect 27944 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28264 35936
rect 27944 34848 28264 35872
rect 32944 53888 33264 54448
rect 32944 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33264 53888
rect 32944 52800 33264 53824
rect 32944 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33264 52800
rect 32944 51712 33264 52736
rect 32944 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33264 51712
rect 32944 50624 33264 51648
rect 32944 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33264 50624
rect 32944 49536 33264 50560
rect 32944 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33264 49536
rect 32944 48448 33264 49472
rect 32944 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33264 48448
rect 32944 47360 33264 48384
rect 32944 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33264 47360
rect 32944 46272 33264 47296
rect 32944 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33264 46272
rect 32944 45184 33264 46208
rect 32944 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33264 45184
rect 32944 44096 33264 45120
rect 37944 54432 38264 54448
rect 37944 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38264 54432
rect 37944 53344 38264 54368
rect 37944 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38264 53344
rect 37944 52256 38264 53280
rect 37944 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38264 52256
rect 37944 51168 38264 52192
rect 37944 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38264 51168
rect 37944 50080 38264 51104
rect 37944 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38264 50080
rect 37944 48992 38264 50016
rect 37944 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38264 48992
rect 37944 47904 38264 48928
rect 37944 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38264 47904
rect 37944 46816 38264 47840
rect 37944 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38264 46816
rect 37944 45728 38264 46752
rect 37944 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38264 45728
rect 35387 44708 35453 44709
rect 35387 44644 35388 44708
rect 35452 44644 35453 44708
rect 35387 44643 35453 44644
rect 32944 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33264 44096
rect 32944 43008 33264 44032
rect 32944 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33264 43008
rect 32944 41920 33264 42944
rect 32944 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33264 41920
rect 32944 40832 33264 41856
rect 32944 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33264 40832
rect 32944 39744 33264 40768
rect 32944 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33264 39744
rect 32944 38656 33264 39680
rect 32944 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33264 38656
rect 32944 37568 33264 38592
rect 32944 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33264 37568
rect 32944 36480 33264 37504
rect 32944 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33264 36480
rect 28395 35732 28461 35733
rect 28395 35668 28396 35732
rect 28460 35668 28461 35732
rect 28395 35667 28461 35668
rect 27944 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28264 34848
rect 27944 33760 28264 34784
rect 27944 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28264 33760
rect 27107 32876 27173 32877
rect 27107 32812 27108 32876
rect 27172 32812 27173 32876
rect 27107 32811 27173 32812
rect 26003 24716 26069 24717
rect 26003 24652 26004 24716
rect 26068 24652 26069 24716
rect 26003 24651 26069 24652
rect 25635 24308 25701 24309
rect 25635 24244 25636 24308
rect 25700 24244 25701 24308
rect 25635 24243 25701 24244
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22691 22948 22757 22949
rect 22691 22884 22692 22948
rect 22756 22884 22757 22948
rect 22691 22883 22757 22884
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 22694 2957 22754 22883
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22691 2956 22757 2957
rect 22691 2892 22692 2956
rect 22756 2892 22757 2956
rect 22691 2891 22757 2892
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 25638 1869 25698 24243
rect 26006 2413 26066 24651
rect 26739 19276 26805 19277
rect 26739 19212 26740 19276
rect 26804 19212 26805 19276
rect 26739 19211 26805 19212
rect 26003 2412 26069 2413
rect 26003 2348 26004 2412
rect 26068 2348 26069 2412
rect 26003 2347 26069 2348
rect 26742 2005 26802 19211
rect 27110 18869 27170 32811
rect 27944 32672 28264 33696
rect 27944 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28264 32672
rect 27944 31584 28264 32608
rect 28398 31653 28458 35667
rect 32944 35392 33264 36416
rect 32944 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33264 35392
rect 28579 34644 28645 34645
rect 28579 34580 28580 34644
rect 28644 34580 28645 34644
rect 28579 34579 28645 34580
rect 28395 31652 28461 31653
rect 28395 31588 28396 31652
rect 28460 31588 28461 31652
rect 28395 31587 28461 31588
rect 27944 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28264 31584
rect 27944 30496 28264 31520
rect 28582 31517 28642 34579
rect 32944 34304 33264 35328
rect 32944 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33264 34304
rect 32944 33216 33264 34240
rect 32944 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33264 33216
rect 32944 32128 33264 33152
rect 35390 33013 35450 44643
rect 37944 44640 38264 45664
rect 37944 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38264 44640
rect 36675 44300 36741 44301
rect 36675 44236 36676 44300
rect 36740 44236 36741 44300
rect 36675 44235 36741 44236
rect 37227 44300 37293 44301
rect 37227 44236 37228 44300
rect 37292 44236 37293 44300
rect 37227 44235 37293 44236
rect 35939 43484 36005 43485
rect 35939 43420 35940 43484
rect 36004 43420 36005 43484
rect 35939 43419 36005 43420
rect 35387 33012 35453 33013
rect 35387 32948 35388 33012
rect 35452 32948 35453 33012
rect 35387 32947 35453 32948
rect 32944 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33264 32128
rect 28579 31516 28645 31517
rect 28579 31452 28580 31516
rect 28644 31452 28645 31516
rect 28579 31451 28645 31452
rect 27944 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28264 30496
rect 27944 29408 28264 30432
rect 27944 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28264 29408
rect 27944 28320 28264 29344
rect 27944 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28264 28320
rect 27944 27232 28264 28256
rect 27944 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28264 27232
rect 27944 26144 28264 27168
rect 32944 31040 33264 32064
rect 32944 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33264 31040
rect 32944 29952 33264 30976
rect 35942 30293 36002 43419
rect 36678 30973 36738 44235
rect 36675 30972 36741 30973
rect 36675 30908 36676 30972
rect 36740 30908 36741 30972
rect 36675 30907 36741 30908
rect 37230 30429 37290 44235
rect 37944 43552 38264 44576
rect 37944 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38264 43552
rect 37944 42464 38264 43488
rect 37944 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38264 42464
rect 37944 41376 38264 42400
rect 42944 53888 43264 54448
rect 42944 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43264 53888
rect 42944 52800 43264 53824
rect 42944 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43264 52800
rect 42944 51712 43264 52736
rect 42944 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43264 51712
rect 42944 50624 43264 51648
rect 42944 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43264 50624
rect 42944 49536 43264 50560
rect 42944 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43264 49536
rect 42944 48448 43264 49472
rect 42944 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43264 48448
rect 42944 47360 43264 48384
rect 42944 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43264 47360
rect 42944 46272 43264 47296
rect 42944 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43264 46272
rect 42944 45184 43264 46208
rect 42944 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43264 45184
rect 42944 44096 43264 45120
rect 42944 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43264 44096
rect 42944 43008 43264 44032
rect 42944 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43264 43008
rect 39987 42124 40053 42125
rect 39987 42060 39988 42124
rect 40052 42060 40053 42124
rect 39987 42059 40053 42060
rect 37944 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38264 41376
rect 37944 40288 38264 41312
rect 37944 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38264 40288
rect 37944 39200 38264 40224
rect 37944 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38264 39200
rect 37944 38112 38264 39136
rect 37944 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38264 38112
rect 37944 37024 38264 38048
rect 37944 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38264 37024
rect 37944 35936 38264 36960
rect 37944 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38264 35936
rect 37944 34848 38264 35872
rect 38331 35732 38397 35733
rect 38331 35668 38332 35732
rect 38396 35668 38397 35732
rect 38331 35667 38397 35668
rect 37944 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38264 34848
rect 37944 33760 38264 34784
rect 37944 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38264 33760
rect 37944 32672 38264 33696
rect 37944 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38264 32672
rect 37944 31584 38264 32608
rect 38334 32469 38394 35667
rect 38331 32468 38397 32469
rect 38331 32404 38332 32468
rect 38396 32404 38397 32468
rect 38331 32403 38397 32404
rect 38515 31788 38581 31789
rect 38515 31724 38516 31788
rect 38580 31724 38581 31788
rect 38515 31723 38581 31724
rect 37944 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38264 31584
rect 37944 30496 38264 31520
rect 37944 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38264 30496
rect 37227 30428 37293 30429
rect 37227 30364 37228 30428
rect 37292 30364 37293 30428
rect 37227 30363 37293 30364
rect 35939 30292 36005 30293
rect 35939 30228 35940 30292
rect 36004 30228 36005 30292
rect 35939 30227 36005 30228
rect 32944 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33264 29952
rect 32944 28864 33264 29888
rect 32944 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33264 28864
rect 32944 27776 33264 28800
rect 32944 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33264 27776
rect 30603 26892 30669 26893
rect 30603 26828 30604 26892
rect 30668 26828 30669 26892
rect 30603 26827 30669 26828
rect 27944 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28264 26144
rect 27944 25056 28264 26080
rect 30419 25260 30485 25261
rect 30419 25196 30420 25260
rect 30484 25196 30485 25260
rect 30419 25195 30485 25196
rect 27944 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28264 25056
rect 27944 23968 28264 24992
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 30422 20637 30482 25195
rect 30419 20636 30485 20637
rect 30419 20572 30420 20636
rect 30484 20572 30485 20636
rect 30419 20571 30485 20572
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27107 18868 27173 18869
rect 27107 18804 27108 18868
rect 27172 18804 27173 18868
rect 27107 18803 27173 18804
rect 27110 3093 27170 18803
rect 27659 18732 27725 18733
rect 27659 18668 27660 18732
rect 27724 18668 27725 18732
rect 27659 18667 27725 18668
rect 27662 17101 27722 18667
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 30606 18053 30666 26827
rect 32944 26688 33264 27712
rect 32944 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33264 26688
rect 32944 25600 33264 26624
rect 32944 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33264 25600
rect 32944 24512 33264 25536
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 30603 18052 30669 18053
rect 30603 17988 30604 18052
rect 30668 17988 30669 18052
rect 30603 17987 30669 17988
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27659 17100 27725 17101
rect 27659 17036 27660 17100
rect 27724 17036 27725 17100
rect 27659 17035 27725 17036
rect 27107 3092 27173 3093
rect 27107 3028 27108 3092
rect 27172 3028 27173 3092
rect 27107 3027 27173 3028
rect 27662 2549 27722 17035
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 30606 12885 30666 17987
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 30603 12884 30669 12885
rect 30603 12820 30604 12884
rect 30668 12820 30669 12884
rect 30603 12819 30669 12820
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27659 2548 27725 2549
rect 27659 2484 27660 2548
rect 27724 2484 27725 2548
rect 27659 2483 27725 2484
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 29408 38264 30432
rect 37944 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38264 29408
rect 37944 28320 38264 29344
rect 37944 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38264 28320
rect 37944 27232 38264 28256
rect 38518 27437 38578 31723
rect 38515 27436 38581 27437
rect 38515 27372 38516 27436
rect 38580 27372 38581 27436
rect 38515 27371 38581 27372
rect 37944 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38264 27232
rect 37944 26144 38264 27168
rect 39990 27029 40050 42059
rect 42944 41920 43264 42944
rect 42944 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43264 41920
rect 40539 41716 40605 41717
rect 40539 41652 40540 41716
rect 40604 41652 40605 41716
rect 40539 41651 40605 41652
rect 40542 28525 40602 41651
rect 42944 40832 43264 41856
rect 42944 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43264 40832
rect 42944 39744 43264 40768
rect 42944 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43264 39744
rect 42944 38656 43264 39680
rect 42944 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43264 38656
rect 42944 37568 43264 38592
rect 42944 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43264 37568
rect 42944 36480 43264 37504
rect 42944 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43264 36480
rect 42944 35392 43264 36416
rect 42944 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43264 35392
rect 42944 34304 43264 35328
rect 42944 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43264 34304
rect 42944 33216 43264 34240
rect 42944 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43264 33216
rect 42944 32128 43264 33152
rect 42944 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43264 32128
rect 42944 31040 43264 32064
rect 42944 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43264 31040
rect 42944 29952 43264 30976
rect 42944 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43264 29952
rect 42944 28864 43264 29888
rect 42944 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43264 28864
rect 40539 28524 40605 28525
rect 40539 28460 40540 28524
rect 40604 28460 40605 28524
rect 40539 28459 40605 28460
rect 42944 27776 43264 28800
rect 42944 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43264 27776
rect 39987 27028 40053 27029
rect 39987 26964 39988 27028
rect 40052 26964 40053 27028
rect 39987 26963 40053 26964
rect 37944 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38264 26144
rect 37944 25056 38264 26080
rect 37944 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38264 25056
rect 37944 23968 38264 24992
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 26688 43264 27712
rect 42944 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43264 26688
rect 42944 25600 43264 26624
rect 42944 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43264 25600
rect 42944 24512 43264 25536
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 54432 48264 54448
rect 47944 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48264 54432
rect 47944 53344 48264 54368
rect 47944 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48264 53344
rect 47944 52256 48264 53280
rect 47944 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48264 52256
rect 47944 51168 48264 52192
rect 47944 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48264 51168
rect 47944 50080 48264 51104
rect 47944 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48264 50080
rect 47944 48992 48264 50016
rect 47944 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48264 48992
rect 47944 47904 48264 48928
rect 47944 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48264 47904
rect 47944 46816 48264 47840
rect 47944 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48264 46816
rect 47944 45728 48264 46752
rect 47944 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48264 45728
rect 47944 44640 48264 45664
rect 47944 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48264 44640
rect 47944 43552 48264 44576
rect 47944 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48264 43552
rect 47944 42464 48264 43488
rect 47944 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48264 42464
rect 47944 41376 48264 42400
rect 47944 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48264 41376
rect 47944 40288 48264 41312
rect 47944 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48264 40288
rect 47944 39200 48264 40224
rect 47944 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48264 39200
rect 47944 38112 48264 39136
rect 47944 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48264 38112
rect 47944 37024 48264 38048
rect 47944 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48264 37024
rect 47944 35936 48264 36960
rect 47944 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48264 35936
rect 47944 34848 48264 35872
rect 47944 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48264 34848
rect 47944 33760 48264 34784
rect 47944 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48264 33760
rect 47944 32672 48264 33696
rect 47944 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48264 32672
rect 47944 31584 48264 32608
rect 47944 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48264 31584
rect 47944 30496 48264 31520
rect 47944 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48264 30496
rect 47944 29408 48264 30432
rect 47944 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48264 29408
rect 47944 28320 48264 29344
rect 47944 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48264 28320
rect 47944 27232 48264 28256
rect 47944 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48264 27232
rect 47944 26144 48264 27168
rect 47944 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48264 26144
rect 47944 25056 48264 26080
rect 47944 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48264 25056
rect 47944 23968 48264 24992
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
rect 26739 2004 26805 2005
rect 26739 1940 26740 2004
rect 26804 1940 26805 2004
rect 26739 1939 26805 1940
rect 25635 1868 25701 1869
rect 25635 1804 25636 1868
rect 25700 1804 25701 1868
rect 25635 1803 25701 1804
use sky130_fd_sc_hd__clkbuf_2  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 45632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _111_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 46000 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 46092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 46184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 45356 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 29992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 44252 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 43700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 40572 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 42872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 43608 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 43608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 44344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 44068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform 1 0 44068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 43700 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 44160 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform 1 0 44344 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 45172 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 45908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 46736 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 46000 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1676037725
transform 1 0 47104 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 47748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1676037725
transform 1 0 46828 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 47932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 25760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 25576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 24288 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 27140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 27876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 28888 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 28704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 28612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 33028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 33764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 31464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 34040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 36156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 37076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 38180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 35880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 35696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 38916 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 36432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _165_
timestamp 1676037725
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1676037725
transform 1 0 5612 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 6992 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 7728 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 12144 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1676037725
transform 1 0 9108 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform 1 0 10580 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1676037725
transform 1 0 12880 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1676037725
transform 1 0 11960 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform 1 0 12052 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1676037725
transform 1 0 14260 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1676037725
transform 1 0 14168 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform 1 0 16008 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _183_
timestamp 1676037725
transform 1 0 14536 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform 1 0 16744 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform 1 0 17112 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform 1 0 18952 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1676037725
transform 1 0 17940 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform 1 0 20240 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 20148 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1676037725
transform 1 0 21068 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform 1 0 20148 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1676037725
transform 1 0 20056 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1676037725
transform 1 0 22632 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform 1 0 21988 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _195_
timestamp 1676037725
transform 1 0 23000 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 24656 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 23552 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _199_
timestamp 1676037725
transform 1 0 4508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _200_
timestamp 1676037725
transform 1 0 4048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _201_
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _202_
timestamp 1676037725
transform 1 0 5244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _203_
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1676037725
transform 1 0 4968 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1676037725
transform 1 0 4784 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1676037725
transform 1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1676037725
transform 1 0 48576 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1676037725
transform 1 0 46184 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _210_
timestamp 1676037725
transform 1 0 47748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1676037725
transform 1 0 48576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _212_
timestamp 1676037725
transform 1 0 48576 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 47932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 47932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 25024 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 26496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 27232 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 31464 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 34868 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 12420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 22724 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 28428 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 29440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 33488 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 23184 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 27784 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 36156 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 21620 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 21160 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 20884 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 25024 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 26036 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 27692 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 41216 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 39192 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 39376 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 23184 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 35328 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 30912 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 22264 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 21160 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 21068 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 37628 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 32936 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 15456 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 33488 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1676037725
transform 1 0 19688 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1676037725
transform 1 0 35696 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1676037725
transform 1 0 29900 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1676037725
transform 1 0 36156 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1676037725
transform 1 0 30912 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1676037725
transform 1 0 36064 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1676037725
transform 1 0 38640 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24564 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21804 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 19596 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23000 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24748 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26496 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27324 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 25852 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__265 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 19320 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28796 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28428 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28244 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 27140 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 23000 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25760 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__266
timestamp 1676037725
transform 1 0 25760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 24564 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29992 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28244 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28428 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 27232 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 23276 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25944 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 20700 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__267
timestamp 1676037725
transform 1 0 23552 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 22816 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24012 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27324 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 26772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 25024 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 20516 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 22264 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__268
timestamp 1676037725
transform 1 0 22724 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7636 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 7544 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 7728 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 10672 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 8832 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12328 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 7820 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 8372 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 12604 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 7544 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 9568 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27048 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21712 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 28244 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 20516 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 21160 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 23644 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 34868 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 32936 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 36892 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 37720 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 31832 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 30636 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 37076 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 35972 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43
timestamp 1676037725
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 1676037725
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123
timestamp 1676037725
transform 1 0 12420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1676037725
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1676037725
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1676037725
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1676037725
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1676037725
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1676037725
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1676037725
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1676037725
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1676037725
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1676037725
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1676037725
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_467
timestamp 1676037725
transform 1 0 44068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_481
timestamp 1676037725
transform 1 0 45356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1676037725
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_523
timestamp 1676037725
transform 1 0 49220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_16 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_28
timestamp 1676037725
transform 1 0 3680 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1676037725
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1676037725
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_77
timestamp 1676037725
transform 1 0 8188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_129
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1676037725
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_185
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_257
timestamp 1676037725
transform 1 0 24748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1676037725
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1676037725
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_321
timestamp 1676037725
transform 1 0 30636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1676037725
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_355
timestamp 1676037725
transform 1 0 33764 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_375
timestamp 1676037725
transform 1 0 35604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1676037725
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_411
timestamp 1676037725
transform 1 0 38916 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_431
timestamp 1676037725
transform 1 0 40756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1676037725
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_467
timestamp 1676037725
transform 1 0 44068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1676037725
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_491
timestamp 1676037725
transform 1 0 46276 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1676037725
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1676037725
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1676037725
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_271
timestamp 1676037725
transform 1 0 26036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_283
timestamp 1676037725
transform 1 0 27140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_295
timestamp 1676037725
transform 1 0 28244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_327
timestamp 1676037725
transform 1 0 31188 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_347
timestamp 1676037725
transform 1 0 33028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1676037725
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1676037725
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1676037725
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1676037725
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_439
timestamp 1676037725
transform 1 0 41492 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_459
timestamp 1676037725
transform 1 0 43332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_471
timestamp 1676037725
transform 1 0 44436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_495
timestamp 1676037725
transform 1 0 46644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_507
timestamp 1676037725
transform 1 0 47748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_477
timestamp 1676037725
transform 1 0 44988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_489
timestamp 1676037725
transform 1 0 46092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_501
timestamp 1676037725
transform 1 0 47196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_513
timestamp 1676037725
transform 1 0 48300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_310
timestamp 1676037725
transform 1 0 29624 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_318
timestamp 1676037725
transform 1 0 30360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_330
timestamp 1676037725
transform 1 0 31464 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_521
timestamp 1676037725
transform 1 0 49036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1676037725
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_520
timestamp 1676037725
transform 1 0 48944 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_526
timestamp 1676037725
transform 1 0 49496 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_399
timestamp 1676037725
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_407
timestamp 1676037725
transform 1 0 38548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_504
timestamp 1676037725
transform 1 0 47472 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_508
timestamp 1676037725
transform 1 0 47840 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_380
timestamp 1676037725
transform 1 0 36064 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_399
timestamp 1676037725
transform 1 0 37812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_411
timestamp 1676037725
transform 1 0 38916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_423
timestamp 1676037725
transform 1 0 40020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_435
timestamp 1676037725
transform 1 0 41124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_381
timestamp 1676037725
transform 1 0 36156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1676037725
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_403
timestamp 1676037725
transform 1 0 38180 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_415
timestamp 1676037725
transform 1 0 39284 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_427
timestamp 1676037725
transform 1 0 40388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_439
timestamp 1676037725
transform 1 0 41492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_481
timestamp 1676037725
transform 1 0 45356 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_488
timestamp 1676037725
transform 1 0 46000 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_500
timestamp 1676037725
transform 1 0 47104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_485
timestamp 1676037725
transform 1 0 45724 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_491
timestamp 1676037725
transform 1 0 46276 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_503
timestamp 1676037725
transform 1 0 47380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_515
timestamp 1676037725
transform 1 0 48484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_343
timestamp 1676037725
transform 1 0 32660 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_355
timestamp 1676037725
transform 1 0 33764 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_367
timestamp 1676037725
transform 1 0 34868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_375
timestamp 1676037725
transform 1 0 35604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_382
timestamp 1676037725
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_491
timestamp 1676037725
transform 1 0 46276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1676037725
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1676037725
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_337
timestamp 1676037725
transform 1 0 32108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_349
timestamp 1676037725
transform 1 0 33212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1676037725
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1676037725
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_256
timestamp 1676037725
transform 1 0 24656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_268
timestamp 1676037725
transform 1 0 25760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_429
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_433
timestamp 1676037725
transform 1 0 40940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_445
timestamp 1676037725
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_146
timestamp 1676037725
transform 1 0 14536 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_158
timestamp 1676037725
transform 1 0 15640 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_182
timestamp 1676037725
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1676037725
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1676037725
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1676037725
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1676037725
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1676037725
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_494
timestamp 1676037725
transform 1 0 46552 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_506
timestamp 1676037725
transform 1 0 47656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1676037725
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1676037725
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_437
timestamp 1676037725
transform 1 0 41308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_442
timestamp 1676037725
transform 1 0 41768 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_477
timestamp 1676037725
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1676037725
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1676037725
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1676037725
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_297
timestamp 1676037725
transform 1 0 28428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1676037725
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_386
timestamp 1676037725
transform 1 0 36616 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_398
timestamp 1676037725
transform 1 0 37720 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_410
timestamp 1676037725
transform 1 0 38824 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_415
timestamp 1676037725
transform 1 0 39284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_439
timestamp 1676037725
transform 1 0 41492 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_451
timestamp 1676037725
transform 1 0 42596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_463
timestamp 1676037725
transform 1 0 43700 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_472
timestamp 1676037725
transform 1 0 44528 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1676037725
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_287
timestamp 1676037725
transform 1 0 27508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_295
timestamp 1676037725
transform 1 0 28244 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_310
timestamp 1676037725
transform 1 0 29624 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_323
timestamp 1676037725
transform 1 0 30820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_353
timestamp 1676037725
transform 1 0 33580 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_374
timestamp 1676037725
transform 1 0 35512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1676037725
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_467
timestamp 1676037725
transform 1 0 44068 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_479
timestamp 1676037725
transform 1 0 45172 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_491
timestamp 1676037725
transform 1 0 46276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_270
timestamp 1676037725
transform 1 0 25944 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_282
timestamp 1676037725
transform 1 0 27048 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_294
timestamp 1676037725
transform 1 0 28152 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1676037725
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1676037725
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_387
timestamp 1676037725
transform 1 0 36708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_395
timestamp 1676037725
transform 1 0 37444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_399
timestamp 1676037725
transform 1 0 37812 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_403
timestamp 1676037725
transform 1 0 38180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_415
timestamp 1676037725
transform 1 0 39284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1676037725
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1676037725
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1676037725
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1676037725
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_301
timestamp 1676037725
transform 1 0 28796 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_306
timestamp 1676037725
transform 1 0 29256 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_321
timestamp 1676037725
transform 1 0 30636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1676037725
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_349
timestamp 1676037725
transform 1 0 33212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_355
timestamp 1676037725
transform 1 0 33764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_376
timestamp 1676037725
transform 1 0 35696 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_384
timestamp 1676037725
transform 1 0 36432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1676037725
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_399
timestamp 1676037725
transform 1 0 37812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_407
timestamp 1676037725
transform 1 0 38548 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_414
timestamp 1676037725
transform 1 0 39192 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_426
timestamp 1676037725
transform 1 0 40296 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_438
timestamp 1676037725
transform 1 0 41400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1676037725
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1676037725
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_339
timestamp 1676037725
transform 1 0 32292 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_352
timestamp 1676037725
transform 1 0 33488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_371
timestamp 1676037725
transform 1 0 35236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_383
timestamp 1676037725
transform 1 0 36340 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_391
timestamp 1676037725
transform 1 0 37076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_401
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_408
timestamp 1676037725
transform 1 0 38640 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_426
timestamp 1676037725
transform 1 0 40296 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_438
timestamp 1676037725
transform 1 0 41400 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_450
timestamp 1676037725
transform 1 0 42504 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_462
timestamp 1676037725
transform 1 0 43608 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1676037725
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_231
timestamp 1676037725
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_252
timestamp 1676037725
transform 1 0 24288 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_268
timestamp 1676037725
transform 1 0 25760 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_309
timestamp 1676037725
transform 1 0 29532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_317
timestamp 1676037725
transform 1 0 30268 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_324
timestamp 1676037725
transform 1 0 30912 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_348
timestamp 1676037725
transform 1 0 33120 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_360
timestamp 1676037725
transform 1 0 34224 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_372
timestamp 1676037725
transform 1 0 35328 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_384
timestamp 1676037725
transform 1 0 36432 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_404
timestamp 1676037725
transform 1 0 38272 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_416
timestamp 1676037725
transform 1 0 39376 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_428
timestamp 1676037725
transform 1 0 40480 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_440
timestamp 1676037725
transform 1 0 41584 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_445
timestamp 1676037725
transform 1 0 42044 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_259
timestamp 1676037725
transform 1 0 24932 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_267
timestamp 1676037725
transform 1 0 25668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_272
timestamp 1676037725
transform 1 0 26128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_285
timestamp 1676037725
transform 1 0 27324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_298
timestamp 1676037725
transform 1 0 28520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_331
timestamp 1676037725
transform 1 0 31556 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_339
timestamp 1676037725
transform 1 0 32292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_343
timestamp 1676037725
transform 1 0 32660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1676037725
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_397
timestamp 1676037725
transform 1 0 37628 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_409
timestamp 1676037725
transform 1 0 38732 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_417
timestamp 1676037725
transform 1 0 39468 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_258
timestamp 1676037725
transform 1 0 24840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_262
timestamp 1676037725
transform 1 0 25208 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_272
timestamp 1676037725
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_292
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_300
timestamp 1676037725
transform 1 0 28704 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_321
timestamp 1676037725
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1676037725
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_345
timestamp 1676037725
transform 1 0 32844 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1676037725
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_362
timestamp 1676037725
transform 1 0 34408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_369
timestamp 1676037725
transform 1 0 35052 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_377
timestamp 1676037725
transform 1 0 35788 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_383
timestamp 1676037725
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_398
timestamp 1676037725
transform 1 0 37720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_406
timestamp 1676037725
transform 1 0 38456 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_412
timestamp 1676037725
transform 1 0 39008 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_424
timestamp 1676037725
transform 1 0 40112 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_436
timestamp 1676037725
transform 1 0 41216 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_51
timestamp 1676037725
transform 1 0 5796 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_63
timestamp 1676037725
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1676037725
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1676037725
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1676037725
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_278
timestamp 1676037725
transform 1 0 26680 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_282
timestamp 1676037725
transform 1 0 27048 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_292
timestamp 1676037725
transform 1 0 27968 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1676037725
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_387
timestamp 1676037725
transform 1 0 36708 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_404
timestamp 1676037725
transform 1 0 38272 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1676037725
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1676037725
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_201
timestamp 1676037725
transform 1 0 19596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_233
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1676037725
transform 1 0 23644 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_258
timestamp 1676037725
transform 1 0 24840 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1676037725
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_306
timestamp 1676037725
transform 1 0 29256 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_342
timestamp 1676037725
transform 1 0 32568 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_350
timestamp 1676037725
transform 1 0 33304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_362
timestamp 1676037725
transform 1 0 34408 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1676037725
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_382
timestamp 1676037725
transform 1 0 36248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1676037725
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_399
timestamp 1676037725
transform 1 0 37812 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_403
timestamp 1676037725
transform 1 0 38180 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_415
timestamp 1676037725
transform 1 0 39284 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_427
timestamp 1676037725
transform 1 0 40388 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_439
timestamp 1676037725
transform 1 0 41492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_466
timestamp 1676037725
transform 1 0 43976 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_478
timestamp 1676037725
transform 1 0 45080 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_490
timestamp 1676037725
transform 1 0 46184 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_502
timestamp 1676037725
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_203
timestamp 1676037725
transform 1 0 19780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_213
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_240
timestamp 1676037725
transform 1 0 23184 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1676037725
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_277
timestamp 1676037725
transform 1 0 26588 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_294
timestamp 1676037725
transform 1 0 28152 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_317
timestamp 1676037725
transform 1 0 30268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_341
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_349
timestamp 1676037725
transform 1 0 33212 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1676037725
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_373
timestamp 1676037725
transform 1 0 35420 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_394
timestamp 1676037725
transform 1 0 37352 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1676037725
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_445
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_453
timestamp 1676037725
transform 1 0 42780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_458
timestamp 1676037725
transform 1 0 43240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_466
timestamp 1676037725
transform 1 0 43976 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1676037725
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1676037725
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_212
timestamp 1676037725
transform 1 0 20608 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1676037725
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1676037725
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1676037725
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_294
timestamp 1676037725
transform 1 0 28152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_306
timestamp 1676037725
transform 1 0 29256 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_321
timestamp 1676037725
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1676037725
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_359
timestamp 1676037725
transform 1 0 34132 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_383
timestamp 1676037725
transform 1 0 36340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_404
timestamp 1676037725
transform 1 0 38272 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_416
timestamp 1676037725
transform 1 0 39376 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_428
timestamp 1676037725
transform 1 0 40480 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_440
timestamp 1676037725
transform 1 0 41584 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_220
timestamp 1676037725
transform 1 0 21344 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_235
timestamp 1676037725
transform 1 0 22724 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_279
timestamp 1676037725
transform 1 0 26772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_305
timestamp 1676037725
transform 1 0 29164 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_321
timestamp 1676037725
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_334
timestamp 1676037725
transform 1 0 31832 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_346
timestamp 1676037725
transform 1 0 32936 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1676037725
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_385
timestamp 1676037725
transform 1 0 36524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_409
timestamp 1676037725
transform 1 0 38732 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_417
timestamp 1676037725
transform 1 0 39468 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1676037725
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_457
timestamp 1676037725
transform 1 0 43148 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_465
timestamp 1676037725
transform 1 0 43884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1676037725
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1676037725
transform 1 0 19412 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_209
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_251
timestamp 1676037725
transform 1 0 24196 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1676037725
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_321
timestamp 1676037725
transform 1 0 30636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1676037725
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_353
timestamp 1676037725
transform 1 0 33580 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_375
timestamp 1676037725
transform 1 0 35604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_415
timestamp 1676037725
transform 1 0 39284 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_427
timestamp 1676037725
transform 1 0 40388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_439
timestamp 1676037725
transform 1 0 41492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_158
timestamp 1676037725
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_182
timestamp 1676037725
transform 1 0 17848 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1676037725
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_261
timestamp 1676037725
transform 1 0 25116 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_271
timestamp 1676037725
transform 1 0 26036 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_288
timestamp 1676037725
transform 1 0 27600 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1676037725
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_337
timestamp 1676037725
transform 1 0 32108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_342
timestamp 1676037725
transform 1 0 32568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_346
timestamp 1676037725
transform 1 0 32936 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_351
timestamp 1676037725
transform 1 0 33396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1676037725
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_371
timestamp 1676037725
transform 1 0 35236 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_378
timestamp 1676037725
transform 1 0 35880 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_390
timestamp 1676037725
transform 1 0 36984 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_402
timestamp 1676037725
transform 1 0 38088 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_414
timestamp 1676037725
transform 1 0 39192 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_465
timestamp 1676037725
transform 1 0 43884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_471
timestamp 1676037725
transform 1 0 44436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_33
timestamp 1676037725
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_45
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1676037725
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_260
timestamp 1676037725
transform 1 0 25024 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1676037725
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1676037725
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1676037725
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_313
timestamp 1676037725
transform 1 0 29900 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_323
timestamp 1676037725
transform 1 0 30820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1676037725
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1676037725
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_385
timestamp 1676037725
transform 1 0 36524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1676037725
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1676037725
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_36
timestamp 1676037725
transform 1 0 4416 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_48
timestamp 1676037725
transform 1 0 5520 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_60
timestamp 1676037725
transform 1 0 6624 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_72
timestamp 1676037725
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_95
timestamp 1676037725
transform 1 0 9844 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_107
timestamp 1676037725
transform 1 0 10948 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1676037725
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1676037725
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_208
timestamp 1676037725
transform 1 0 20240 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_220
timestamp 1676037725
transform 1 0 21344 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_232
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1676037725
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1676037725
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1676037725
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1676037725
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_326
timestamp 1676037725
transform 1 0 31096 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_340
timestamp 1676037725
transform 1 0 32384 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_352
timestamp 1676037725
transform 1 0 33488 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_385
timestamp 1676037725
transform 1 0 36524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_397
timestamp 1676037725
transform 1 0 37628 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_408
timestamp 1676037725
transform 1 0 38640 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_467
timestamp 1676037725
transform 1 0 44068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_89
timestamp 1676037725
transform 1 0 9292 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1676037725
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_146
timestamp 1676037725
transform 1 0 14536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_158
timestamp 1676037725
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1676037725
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_289
timestamp 1676037725
transform 1 0 27692 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1676037725
transform 1 0 28244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_308
timestamp 1676037725
transform 1 0 29440 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1676037725
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_372
timestamp 1676037725
transform 1 0 35328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_376
timestamp 1676037725
transform 1 0 35696 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_380
timestamp 1676037725
transform 1 0 36064 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_426
timestamp 1676037725
transform 1 0 40296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_438
timestamp 1676037725
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1676037725
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_49
timestamp 1676037725
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1676037725
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1676037725
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_131
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_181
timestamp 1676037725
transform 1 0 17756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_224
timestamp 1676037725
transform 1 0 21712 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1676037725
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_259
timestamp 1676037725
transform 1 0 24932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_262
timestamp 1676037725
transform 1 0 25208 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_275
timestamp 1676037725
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_287
timestamp 1676037725
transform 1 0 27508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_295
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_314
timestamp 1676037725
transform 1 0 29992 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_326
timestamp 1676037725
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_338
timestamp 1676037725
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_350
timestamp 1676037725
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1676037725
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_371
timestamp 1676037725
transform 1 0 35236 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_393
timestamp 1676037725
transform 1 0 37260 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_400
timestamp 1676037725
transform 1 0 37904 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_412
timestamp 1676037725
transform 1 0 39008 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_186
timestamp 1676037725
transform 1 0 18216 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_198
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1676037725
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_212
timestamp 1676037725
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_250
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_254
timestamp 1676037725
transform 1 0 24472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_264
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_271
timestamp 1676037725
transform 1 0 26036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_303
timestamp 1676037725
transform 1 0 28980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_309
timestamp 1676037725
transform 1 0 29532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_319
timestamp 1676037725
transform 1 0 30452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1676037725
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_342
timestamp 1676037725
transform 1 0 32568 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_363
timestamp 1676037725
transform 1 0 34500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_375
timestamp 1676037725
transform 1 0 35604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1676037725
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_419
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_431
timestamp 1676037725
transform 1 0 40756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_443
timestamp 1676037725
transform 1 0 41860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_467
timestamp 1676037725
transform 1 0 44068 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_472
timestamp 1676037725
transform 1 0 44528 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_484
timestamp 1676037725
transform 1 0 45632 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_496
timestamp 1676037725
transform 1 0 46736 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_36
timestamp 1676037725
transform 1 0 4416 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_46
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_58
timestamp 1676037725
transform 1 0 6440 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_70
timestamp 1676037725
transform 1 0 7544 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_90
timestamp 1676037725
transform 1 0 9384 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_102
timestamp 1676037725
transform 1 0 10488 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_114
timestamp 1676037725
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_126
timestamp 1676037725
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_173
timestamp 1676037725
transform 1 0 17020 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_219
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_231
timestamp 1676037725
transform 1 0 22356 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_237
timestamp 1676037725
transform 1 0 22908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1676037725
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_276
timestamp 1676037725
transform 1 0 26496 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_282
timestamp 1676037725
transform 1 0 27048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1676037725
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_335
timestamp 1676037725
transform 1 0 31924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1676037725
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_387
timestamp 1676037725
transform 1 0 36708 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_398
timestamp 1676037725
transform 1 0 37720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_402
timestamp 1676037725
transform 1 0 38088 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_412
timestamp 1676037725
transform 1 0 39008 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_426
timestamp 1676037725
transform 1 0 40296 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_438
timestamp 1676037725
transform 1 0 41400 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_450
timestamp 1676037725
transform 1 0 42504 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_462
timestamp 1676037725
transform 1 0 43608 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1676037725
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_92
timestamp 1676037725
transform 1 0 9568 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1676037725
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_121
timestamp 1676037725
transform 1 0 12236 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1676037725
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_197
timestamp 1676037725
transform 1 0 19228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_207
timestamp 1676037725
transform 1 0 20148 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_254
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_258
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_265
timestamp 1676037725
transform 1 0 25484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_291
timestamp 1676037725
transform 1 0 27876 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_304
timestamp 1676037725
transform 1 0 29072 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_316
timestamp 1676037725
transform 1 0 30176 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_328
timestamp 1676037725
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_359
timestamp 1676037725
transform 1 0 34132 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_372
timestamp 1676037725
transform 1 0 35328 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_384
timestamp 1676037725
transform 1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1676037725
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1676037725
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_103
timestamp 1676037725
transform 1 0 10580 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_122
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1676037725
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1676037725
transform 1 0 20700 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_234
timestamp 1676037725
transform 1 0 22632 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_259
timestamp 1676037725
transform 1 0 24932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_269
timestamp 1676037725
transform 1 0 25852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_282
timestamp 1676037725
transform 1 0 27048 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_297
timestamp 1676037725
transform 1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1676037725
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_320
timestamp 1676037725
transform 1 0 30544 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_332
timestamp 1676037725
transform 1 0 31648 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_344
timestamp 1676037725
transform 1 0 32752 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_352
timestamp 1676037725
transform 1 0 33488 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_388
timestamp 1676037725
transform 1 0 36800 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1676037725
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1676037725
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_432
timestamp 1676037725
transform 1 0 40848 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_444
timestamp 1676037725
transform 1 0 41952 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_456
timestamp 1676037725
transform 1 0 43056 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_468
timestamp 1676037725
transform 1 0 44160 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_501
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_77
timestamp 1676037725
transform 1 0 8188 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_82
timestamp 1676037725
transform 1 0 8648 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_94
timestamp 1676037725
transform 1 0 9752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1676037725
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_201
timestamp 1676037725
transform 1 0 19596 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_233
timestamp 1676037725
transform 1 0 22540 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_238
timestamp 1676037725
transform 1 0 23000 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_250
timestamp 1676037725
transform 1 0 24104 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_262
timestamp 1676037725
transform 1 0 25208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1676037725
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_303
timestamp 1676037725
transform 1 0 28980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1676037725
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_350
timestamp 1676037725
transform 1 0 33304 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_356
timestamp 1676037725
transform 1 0 33856 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_380
timestamp 1676037725
transform 1 0 36064 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_386
timestamp 1676037725
transform 1 0 36616 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1676037725
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_404
timestamp 1676037725
transform 1 0 38272 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_416
timestamp 1676037725
transform 1 0 39376 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_422
timestamp 1676037725
transform 1 0 39928 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_426
timestamp 1676037725
transform 1 0 40296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_438
timestamp 1676037725
transform 1 0 41400 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1676037725
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_525
timestamp 1676037725
transform 1 0 49404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1676037725
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_45
timestamp 1676037725
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_57
timestamp 1676037725
transform 1 0 6348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_69
timestamp 1676037725
transform 1 0 7452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1676037725
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_146
timestamp 1676037725
transform 1 0 14536 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_158
timestamp 1676037725
transform 1 0 15640 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_170
timestamp 1676037725
transform 1 0 16744 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_229
timestamp 1676037725
transform 1 0 22172 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_239
timestamp 1676037725
transform 1 0 23092 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_264
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_290
timestamp 1676037725
transform 1 0 27784 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1676037725
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_314
timestamp 1676037725
transform 1 0 29992 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_322
timestamp 1676037725
transform 1 0 30728 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_332
timestamp 1676037725
transform 1 0 31648 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_345
timestamp 1676037725
transform 1 0 32844 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_351
timestamp 1676037725
transform 1 0 33396 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1676037725
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_369
timestamp 1676037725
transform 1 0 35052 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_379
timestamp 1676037725
transform 1 0 35972 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_394
timestamp 1676037725
transform 1 0 37352 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_418
timestamp 1676037725
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_432
timestamp 1676037725
transform 1 0 40848 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_444
timestamp 1676037725
transform 1 0 41952 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_456
timestamp 1676037725
transform 1 0 43056 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_468
timestamp 1676037725
transform 1 0 44160 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_474
timestamp 1676037725
transform 1 0 44712 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_483
timestamp 1676037725
transform 1 0 45540 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_491
timestamp 1676037725
transform 1 0 46276 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_503
timestamp 1676037725
transform 1 0 47380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_515
timestamp 1676037725
transform 1 0 48484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_91
timestamp 1676037725
transform 1 0 9476 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_103
timestamp 1676037725
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_245
timestamp 1676037725
transform 1 0 23644 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_255
timestamp 1676037725
transform 1 0 24564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_262
timestamp 1676037725
transform 1 0 25208 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_268
timestamp 1676037725
transform 1 0 25760 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_272
timestamp 1676037725
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_317
timestamp 1676037725
transform 1 0 30268 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1676037725
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_348
timestamp 1676037725
transform 1 0 33120 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_360
timestamp 1676037725
transform 1 0 34224 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_366
timestamp 1676037725
transform 1 0 34776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_376
timestamp 1676037725
transform 1 0 35696 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_384
timestamp 1676037725
transform 1 0 36432 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1676037725
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_404
timestamp 1676037725
transform 1 0 38272 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_417
timestamp 1676037725
transform 1 0 39468 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_425
timestamp 1676037725
transform 1 0 40204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_446
timestamp 1676037725
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1676037725
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1676037725
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_485
timestamp 1676037725
transform 1 0 45724 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_492
timestamp 1676037725
transform 1 0 46368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1676037725
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_521
timestamp 1676037725
transform 1 0 49036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_525
timestamp 1676037725
transform 1 0 49404 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_71
timestamp 1676037725
transform 1 0 7636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_75
timestamp 1676037725
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_95
timestamp 1676037725
transform 1 0 9844 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_107
timestamp 1676037725
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_119
timestamp 1676037725
transform 1 0 12052 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_131
timestamp 1676037725
transform 1 0 13156 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_227
timestamp 1676037725
transform 1 0 21988 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1676037725
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_264
timestamp 1676037725
transform 1 0 25392 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_276
timestamp 1676037725
transform 1 0 26496 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_286
timestamp 1676037725
transform 1 0 27416 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1676037725
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_321
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_331
timestamp 1676037725
transform 1 0 31556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_337
timestamp 1676037725
transform 1 0 32108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_358
timestamp 1676037725
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_378
timestamp 1676037725
transform 1 0 35880 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_386
timestamp 1676037725
transform 1 0 36616 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_400
timestamp 1676037725
transform 1 0 37904 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_408
timestamp 1676037725
transform 1 0 38640 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_418
timestamp 1676037725
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_444
timestamp 1676037725
transform 1 0 41952 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_456
timestamp 1676037725
transform 1 0 43056 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_468
timestamp 1676037725
transform 1 0 44160 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_504
timestamp 1676037725
transform 1 0 47472 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_508
timestamp 1676037725
transform 1 0 47840 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_511
timestamp 1676037725
transform 1 0 48116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_94
timestamp 1676037725
transform 1 0 9752 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 1676037725
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_233
timestamp 1676037725
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_244
timestamp 1676037725
transform 1 0 23552 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_248
timestamp 1676037725
transform 1 0 23920 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_253
timestamp 1676037725
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_265
timestamp 1676037725
transform 1 0 25484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1676037725
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_286
timestamp 1676037725
transform 1 0 27416 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_318
timestamp 1676037725
transform 1 0 30360 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1676037725
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1676037725
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_345
timestamp 1676037725
transform 1 0 32844 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_356
timestamp 1676037725
transform 1 0 33856 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_381
timestamp 1676037725
transform 1 0 36156 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1676037725
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_397
timestamp 1676037725
transform 1 0 37628 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_409
timestamp 1676037725
transform 1 0 38732 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_421
timestamp 1676037725
transform 1 0 39836 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_425
timestamp 1676037725
transform 1 0 40204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_446
timestamp 1676037725
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1676037725
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1676037725
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_500
timestamp 1676037725
transform 1 0 47104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_511
timestamp 1676037725
transform 1 0 48116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_525
timestamp 1676037725
transform 1 0 49404 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1676037725
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_74
timestamp 1676037725
transform 1 0 7912 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1676037725
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_239
timestamp 1676037725
transform 1 0 23092 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1676037725
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_279
timestamp 1676037725
transform 1 0 26772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_287
timestamp 1676037725
transform 1 0 27508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_297
timestamp 1676037725
transform 1 0 28428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1676037725
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_315
timestamp 1676037725
transform 1 0 30084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_325
timestamp 1676037725
transform 1 0 31004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_342
timestamp 1676037725
transform 1 0 32568 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1676037725
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_376
timestamp 1676037725
transform 1 0 35696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_388
timestamp 1676037725
transform 1 0 36800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_410
timestamp 1676037725
transform 1 0 38824 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1676037725
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_444
timestamp 1676037725
transform 1 0 41952 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_456
timestamp 1676037725
transform 1 0 43056 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_464
timestamp 1676037725
transform 1 0 43792 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1676037725
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_497
timestamp 1676037725
transform 1 0 46828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_504
timestamp 1676037725
transform 1 0 47472 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_512
timestamp 1676037725
transform 1 0 48208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1676037725
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_91
timestamp 1676037725
transform 1 0 9476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_103
timestamp 1676037725
transform 1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_231
timestamp 1676037725
transform 1 0 22356 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1676037725
transform 1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1676037725
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_289
timestamp 1676037725
transform 1 0 27692 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_312
timestamp 1676037725
transform 1 0 29808 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_320
timestamp 1676037725
transform 1 0 30544 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1676037725
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_359
timestamp 1676037725
transform 1 0 34132 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_371
timestamp 1676037725
transform 1 0 35236 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1676037725
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_404
timestamp 1676037725
transform 1 0 38272 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1676037725
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1676037725
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1676037725
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1676037725
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1676037725
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1676037725
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_513
timestamp 1676037725
transform 1 0 48300 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_525
timestamp 1676037725
transform 1 0 49404 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_225
timestamp 1676037725
transform 1 0 21804 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_238
timestamp 1676037725
transform 1 0 23000 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_276
timestamp 1676037725
transform 1 0 26496 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1676037725
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_314
timestamp 1676037725
transform 1 0 29992 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_331
timestamp 1676037725
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_343
timestamp 1676037725
transform 1 0 32660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_351
timestamp 1676037725
transform 1 0 33396 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1676037725
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_376
timestamp 1676037725
transform 1 0 35696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_389
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_402
timestamp 1676037725
transform 1 0 38088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_409
timestamp 1676037725
transform 1 0 38732 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_417
timestamp 1676037725
transform 1 0 39468 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_432
timestamp 1676037725
transform 1 0 40848 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_444
timestamp 1676037725
transform 1 0 41952 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_456
timestamp 1676037725
transform 1 0 43056 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_468
timestamp 1676037725
transform 1 0 44160 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_521
timestamp 1676037725
transform 1 0 49036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1676037725
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1676037725
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_236
timestamp 1676037725
transform 1 0 22816 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_242
timestamp 1676037725
transform 1 0 23368 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_254
timestamp 1676037725
transform 1 0 24472 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_266
timestamp 1676037725
transform 1 0 25576 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1676037725
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_309
timestamp 1676037725
transform 1 0 29532 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_322
timestamp 1676037725
transform 1 0 30728 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1676037725
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_377
timestamp 1676037725
transform 1 0 35788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1676037725
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1676037725
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_429
timestamp 1676037725
transform 1 0 40572 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_440
timestamp 1676037725
transform 1 0 41584 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_521
timestamp 1676037725
transform 1 0 49036 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_525
timestamp 1676037725
transform 1 0 49404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1676037725
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_217
timestamp 1676037725
transform 1 0 21068 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_229
timestamp 1676037725
transform 1 0 22172 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1676037725
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1676037725
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_261
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_272
timestamp 1676037725
transform 1 0 26128 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_279
timestamp 1676037725
transform 1 0 26772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_291
timestamp 1676037725
transform 1 0 27876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_303
timestamp 1676037725
transform 1 0 28980 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_320
timestamp 1676037725
transform 1 0 30544 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_332
timestamp 1676037725
transform 1 0 31648 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_344
timestamp 1676037725
transform 1 0 32752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_356
timestamp 1676037725
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_383
timestamp 1676037725
transform 1 0 36340 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_404
timestamp 1676037725
transform 1 0 38272 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_408
timestamp 1676037725
transform 1 0 38640 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_418
timestamp 1676037725
transform 1 0 39560 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_453
timestamp 1676037725
transform 1 0 42780 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_465
timestamp 1676037725
transform 1 0 43884 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_473
timestamp 1676037725
transform 1 0 44620 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_65
timestamp 1676037725
transform 1 0 7084 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_89
timestamp 1676037725
transform 1 0 9292 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_101
timestamp 1676037725
transform 1 0 10396 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_109
timestamp 1676037725
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1676037725
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1676037725
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_241
timestamp 1676037725
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_256
timestamp 1676037725
transform 1 0 24656 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_262
timestamp 1676037725
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1676037725
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1676037725
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_289
timestamp 1676037725
transform 1 0 27692 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_292
timestamp 1676037725
transform 1 0 27968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_315
timestamp 1676037725
transform 1 0 30084 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_328
timestamp 1676037725
transform 1 0 31280 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_353
timestamp 1676037725
transform 1 0 33580 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_363
timestamp 1676037725
transform 1 0 34500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_371
timestamp 1676037725
transform 1 0 35236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_383
timestamp 1676037725
transform 1 0 36340 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_404
timestamp 1676037725
transform 1 0 38272 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_408
timestamp 1676037725
transform 1 0 38640 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_429
timestamp 1676037725
transform 1 0 40572 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_442
timestamp 1676037725
transform 1 0 41768 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_521
timestamp 1676037725
transform 1 0 49036 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_525
timestamp 1676037725
transform 1 0 49404 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_217
timestamp 1676037725
transform 1 0 21068 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_230
timestamp 1676037725
transform 1 0 22264 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_237
timestamp 1676037725
transform 1 0 22908 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1676037725
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_257
timestamp 1676037725
transform 1 0 24748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_278
timestamp 1676037725
transform 1 0 26680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_302
timestamp 1676037725
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_320
timestamp 1676037725
transform 1 0 30544 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_326
timestamp 1676037725
transform 1 0 31096 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_348
timestamp 1676037725
transform 1 0 33120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1676037725
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_392
timestamp 1676037725
transform 1 0 37168 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1676037725
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_407
timestamp 1676037725
transform 1 0 38548 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_417
timestamp 1676037725
transform 1 0 39468 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_432
timestamp 1676037725
transform 1 0 40848 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_436
timestamp 1676037725
transform 1 0 41216 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_440
timestamp 1676037725
transform 1 0 41584 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_447
timestamp 1676037725
transform 1 0 42228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_455
timestamp 1676037725
transform 1 0 42964 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_459
timestamp 1676037725
transform 1 0 43332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_471
timestamp 1676037725
transform 1 0 44436 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1676037725
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1676037725
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_520
timestamp 1676037725
transform 1 0 48944 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_526
timestamp 1676037725
transform 1 0 49496 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_217
timestamp 1676037725
transform 1 0 21068 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_236
timestamp 1676037725
transform 1 0 22816 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_242
timestamp 1676037725
transform 1 0 23368 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_252
timestamp 1676037725
transform 1 0 24288 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1676037725
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_345
timestamp 1676037725
transform 1 0 32844 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_355
timestamp 1676037725
transform 1 0 33764 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_383
timestamp 1676037725
transform 1 0 36340 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1676037725
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_399
timestamp 1676037725
transform 1 0 37812 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_412
timestamp 1676037725
transform 1 0 39008 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_424
timestamp 1676037725
transform 1 0 40112 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_433
timestamp 1676037725
transform 1 0 40940 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_445
timestamp 1676037725
transform 1 0 42044 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_460
timestamp 1676037725
transform 1 0 43424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_472
timestamp 1676037725
transform 1 0 44528 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_480
timestamp 1676037725
transform 1 0 45264 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1676037725
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1676037725
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1676037725
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_511
timestamp 1676037725
transform 1 0 48116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_525
timestamp 1676037725
transform 1 0 49404 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_229
timestamp 1676037725
transform 1 0 22172 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1676037725
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_258
timestamp 1676037725
transform 1 0 24840 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_266
timestamp 1676037725
transform 1 0 25576 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_289
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1676037725
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_348
timestamp 1676037725
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1676037725
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_382
timestamp 1676037725
transform 1 0 36248 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_394
timestamp 1676037725
transform 1 0 37352 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_409
timestamp 1676037725
transform 1 0 38732 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1676037725
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_441
timestamp 1676037725
transform 1 0 41676 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_464
timestamp 1676037725
transform 1 0 43792 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_511
timestamp 1676037725
transform 1 0 48116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_8
timestamp 1676037725
transform 1 0 1840 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_20
timestamp 1676037725
transform 1 0 2944 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_32
timestamp 1676037725
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_44
timestamp 1676037725
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_184
timestamp 1676037725
transform 1 0 18032 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_191
timestamp 1676037725
transform 1 0 18676 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_203
timestamp 1676037725
transform 1 0 19780 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_215
timestamp 1676037725
transform 1 0 20884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_245
timestamp 1676037725
transform 1 0 23644 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_267
timestamp 1676037725
transform 1 0 25668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_302
timestamp 1676037725
transform 1 0 28888 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_314
timestamp 1676037725
transform 1 0 29992 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_326
timestamp 1676037725
transform 1 0 31096 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1676037725
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 1676037725
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1676037725
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_413
timestamp 1676037725
transform 1 0 39100 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_435
timestamp 1676037725
transform 1 0 41124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1676037725
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_454
timestamp 1676037725
transform 1 0 42872 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_466
timestamp 1676037725
transform 1 0 43976 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_474
timestamp 1676037725
transform 1 0 44712 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_478
timestamp 1676037725
transform 1 0 45080 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_490
timestamp 1676037725
transform 1 0 46184 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_502
timestamp 1676037725
transform 1 0 47288 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_513
timestamp 1676037725
transform 1 0 48300 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_525
timestamp 1676037725
transform 1 0 49404 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_237
timestamp 1676037725
transform 1 0 22908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1676037725
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_273
timestamp 1676037725
transform 1 0 26220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_286
timestamp 1676037725
transform 1 0 27416 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_294
timestamp 1676037725
transform 1 0 28152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1676037725
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_320
timestamp 1676037725
transform 1 0 30544 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_376
timestamp 1676037725
transform 1 0 35696 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_402
timestamp 1676037725
transform 1 0 38088 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_414
timestamp 1676037725
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_436
timestamp 1676037725
transform 1 0 41216 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_449
timestamp 1676037725
transform 1 0 42412 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_461
timestamp 1676037725
transform 1 0 43516 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_465
timestamp 1676037725
transform 1 0 43884 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_473
timestamp 1676037725
transform 1 0 44620 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_521
timestamp 1676037725
transform 1 0 49036 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1676037725
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1676037725
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_233
timestamp 1676037725
transform 1 0 22540 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_256
timestamp 1676037725
transform 1 0 24656 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_269
timestamp 1676037725
transform 1 0 25852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1676037725
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_299
timestamp 1676037725
transform 1 0 28612 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_309
timestamp 1676037725
transform 1 0 29532 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_322
timestamp 1676037725
transform 1 0 30728 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1676037725
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_377
timestamp 1676037725
transform 1 0 35788 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_383
timestamp 1676037725
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_404
timestamp 1676037725
transform 1 0 38272 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_419
timestamp 1676037725
transform 1 0 39652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_425
timestamp 1676037725
transform 1 0 40204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_446
timestamp 1676037725
transform 1 0 42136 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_525
timestamp 1676037725
transform 1 0 49404 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1676037725
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_233
timestamp 1676037725
transform 1 0 22540 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1676037725
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_264
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_272
timestamp 1676037725
transform 1 0 26128 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_293
timestamp 1676037725
transform 1 0 28060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1676037725
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_314
timestamp 1676037725
transform 1 0 29992 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_331
timestamp 1676037725
transform 1 0 31556 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_338
timestamp 1676037725
transform 1 0 32200 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_350
timestamp 1676037725
transform 1 0 33304 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1676037725
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_373
timestamp 1676037725
transform 1 0 35420 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_378
timestamp 1676037725
transform 1 0 35880 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_391
timestamp 1676037725
transform 1 0 37076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_399
timestamp 1676037725
transform 1 0 37812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_412
timestamp 1676037725
transform 1 0 39008 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_418
timestamp 1676037725
transform 1 0 39560 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_450
timestamp 1676037725
transform 1 0 42504 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_462
timestamp 1676037725
transform 1 0 43608 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_474
timestamp 1676037725
transform 1 0 44712 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_521
timestamp 1676037725
transform 1 0 49036 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_8
timestamp 1676037725
transform 1 0 1840 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_20
timestamp 1676037725
transform 1 0 2944 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_32
timestamp 1676037725
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_44
timestamp 1676037725
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_259
timestamp 1676037725
transform 1 0 24932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1676037725
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_315
timestamp 1676037725
transform 1 0 30084 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_323
timestamp 1676037725
transform 1 0 30820 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1676037725
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_348
timestamp 1676037725
transform 1 0 33120 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_354
timestamp 1676037725
transform 1 0 33672 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_378
timestamp 1676037725
transform 1 0 35880 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1676037725
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_420
timestamp 1676037725
transform 1 0 39744 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_433
timestamp 1676037725
transform 1 0 40940 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_446
timestamp 1676037725
transform 1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_464
timestamp 1676037725
transform 1 0 43792 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_476
timestamp 1676037725
transform 1 0 44896 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_488
timestamp 1676037725
transform 1 0 46000 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_500
timestamp 1676037725
transform 1 0 47104 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_521
timestamp 1676037725
transform 1 0 49036 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_525
timestamp 1676037725
transform 1 0 49404 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1676037725
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_270
timestamp 1676037725
transform 1 0 25944 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_280
timestamp 1676037725
transform 1 0 26864 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1676037725
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_320
timestamp 1676037725
transform 1 0 30544 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_324
timestamp 1676037725
transform 1 0 30912 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_334
timestamp 1676037725
transform 1 0 31832 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 1676037725
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_388
timestamp 1676037725
transform 1 0 36800 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1676037725
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_416
timestamp 1676037725
transform 1 0 39376 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_433
timestamp 1676037725
transform 1 0 40940 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_441
timestamp 1676037725
transform 1 0 41676 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_445
timestamp 1676037725
transform 1 0 42044 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_451
timestamp 1676037725
transform 1 0 42596 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_472
timestamp 1676037725
transform 1 0 44528 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_521
timestamp 1676037725
transform 1 0 49036 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 1676037725
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1676037725
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1676037725
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_249
timestamp 1676037725
transform 1 0 24012 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_255
timestamp 1676037725
transform 1 0 24564 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1676037725
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_286
timestamp 1676037725
transform 1 0 27416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_298
timestamp 1676037725
transform 1 0 28520 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_324
timestamp 1676037725
transform 1 0 30912 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_330
timestamp 1676037725
transform 1 0 31464 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1676037725
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_348
timestamp 1676037725
transform 1 0 33120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_357
timestamp 1676037725
transform 1 0 33948 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_361
timestamp 1676037725
transform 1 0 34316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_371
timestamp 1676037725
transform 1 0 35236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_384
timestamp 1676037725
transform 1 0 36432 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_401
timestamp 1676037725
transform 1 0 37996 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_422
timestamp 1676037725
transform 1 0 39928 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_435
timestamp 1676037725
transform 1 0 41124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1676037725
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_471
timestamp 1676037725
transform 1 0 44436 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_483
timestamp 1676037725
transform 1 0 45540 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_495
timestamp 1676037725
transform 1 0 46644 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_521
timestamp 1676037725
transform 1 0 49036 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_525
timestamp 1676037725
transform 1 0 49404 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_209
timestamp 1676037725
transform 1 0 20332 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_231
timestamp 1676037725
transform 1 0 22356 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1676037725
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1676037725
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_277
timestamp 1676037725
transform 1 0 26588 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_283
timestamp 1676037725
transform 1 0 27140 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_289
timestamp 1676037725
transform 1 0 27692 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_299
timestamp 1676037725
transform 1 0 28612 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1676037725
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_378
timestamp 1676037725
transform 1 0 35880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_391
timestamp 1676037725
transform 1 0 37076 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_404
timestamp 1676037725
transform 1 0 38272 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_416
timestamp 1676037725
transform 1 0 39376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_441
timestamp 1676037725
transform 1 0 41676 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_452
timestamp 1676037725
transform 1 0 42688 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_464
timestamp 1676037725
transform 1 0 43792 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_8
timestamp 1676037725
transform 1 0 1840 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_20
timestamp 1676037725
transform 1 0 2944 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_32
timestamp 1676037725
transform 1 0 4048 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_44
timestamp 1676037725
transform 1 0 5152 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_208
timestamp 1676037725
transform 1 0 20240 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1676037725
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_233
timestamp 1676037725
transform 1 0 22540 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_238
timestamp 1676037725
transform 1 0 23000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_265
timestamp 1676037725
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1676037725
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_292
timestamp 1676037725
transform 1 0 27968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_304
timestamp 1676037725
transform 1 0 29072 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_312
timestamp 1676037725
transform 1 0 29808 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_322
timestamp 1676037725
transform 1 0 30728 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_330
timestamp 1676037725
transform 1 0 31464 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1676037725
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_348
timestamp 1676037725
transform 1 0 33120 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_360
timestamp 1676037725
transform 1 0 34224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_382
timestamp 1676037725
transform 1 0 36248 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1676037725
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_404
timestamp 1676037725
transform 1 0 38272 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_415
timestamp 1676037725
transform 1 0 39284 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_419
timestamp 1676037725
transform 1 0 39652 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_460
timestamp 1676037725
transform 1 0 43424 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_472
timestamp 1676037725
transform 1 0 44528 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_484
timestamp 1676037725
transform 1 0 45632 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_496
timestamp 1676037725
transform 1 0 46736 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_521
timestamp 1676037725
transform 1 0 49036 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_525
timestamp 1676037725
transform 1 0 49404 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_224
timestamp 1676037725
transform 1 0 21712 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1676037725
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1676037725
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_258
timestamp 1676037725
transform 1 0 24840 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_264
timestamp 1676037725
transform 1 0 25392 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_274
timestamp 1676037725
transform 1 0 26312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_278
timestamp 1676037725
transform 1 0 26680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_299
timestamp 1676037725
transform 1 0 28612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1676037725
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_320
timestamp 1676037725
transform 1 0 30544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_346
timestamp 1676037725
transform 1 0 32936 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_358
timestamp 1676037725
transform 1 0 34040 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1676037725
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_416
timestamp 1676037725
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_432
timestamp 1676037725
transform 1 0 40848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_439
timestamp 1676037725
transform 1 0 41492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_466
timestamp 1676037725
transform 1 0 43976 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_474
timestamp 1676037725
transform 1 0 44712 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_511
timestamp 1676037725
transform 1 0 48116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_231
timestamp 1676037725
transform 1 0 22356 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_235
timestamp 1676037725
transform 1 0 22724 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_259
timestamp 1676037725
transform 1 0 24932 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_271
timestamp 1676037725
transform 1 0 26036 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1676037725
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_306
timestamp 1676037725
transform 1 0 29256 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_317
timestamp 1676037725
transform 1 0 30268 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_332
timestamp 1676037725
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_345
timestamp 1676037725
transform 1 0 32844 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_348
timestamp 1676037725
transform 1 0 33120 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_373
timestamp 1676037725
transform 1 0 35420 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_390
timestamp 1676037725
transform 1 0 36984 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_405
timestamp 1676037725
transform 1 0 38364 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_427
timestamp 1676037725
transform 1 0 40388 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_440
timestamp 1676037725
transform 1 0 41584 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_460
timestamp 1676037725
transform 1 0 43424 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_472
timestamp 1676037725
transform 1 0 44528 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_484
timestamp 1676037725
transform 1 0 45632 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_496
timestamp 1676037725
transform 1 0 46736 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_521
timestamp 1676037725
transform 1 0 49036 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_525
timestamp 1676037725
transform 1 0 49404 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_237
timestamp 1676037725
transform 1 0 22908 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1676037725
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_273
timestamp 1676037725
transform 1 0 26220 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_278
timestamp 1676037725
transform 1 0 26680 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_291
timestamp 1676037725
transform 1 0 27876 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1676037725
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1676037725
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_387
timestamp 1676037725
transform 1 0 36708 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_402
timestamp 1676037725
transform 1 0 38088 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_416
timestamp 1676037725
transform 1 0 39376 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_432
timestamp 1676037725
transform 1 0 40848 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_438
timestamp 1676037725
transform 1 0 41400 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_459
timestamp 1676037725
transform 1 0 43332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_471
timestamp 1676037725
transform 1 0 44436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_521
timestamp 1676037725
transform 1 0 49036 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_8
timestamp 1676037725
transform 1 0 1840 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_20
timestamp 1676037725
transform 1 0 2944 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_32
timestamp 1676037725
transform 1 0 4048 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_44
timestamp 1676037725
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_229
timestamp 1676037725
transform 1 0 22172 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_232
timestamp 1676037725
transform 1 0 22448 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_245
timestamp 1676037725
transform 1 0 23644 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_253
timestamp 1676037725
transform 1 0 24380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_263
timestamp 1676037725
transform 1 0 25300 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1676037725
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_294
timestamp 1676037725
transform 1 0 28152 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_307
timestamp 1676037725
transform 1 0 29348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_319
timestamp 1676037725
transform 1 0 30452 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_323
timestamp 1676037725
transform 1 0 30820 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_326
timestamp 1676037725
transform 1 0 31096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_332
timestamp 1676037725
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_353
timestamp 1676037725
transform 1 0 33580 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_363
timestamp 1676037725
transform 1 0 34500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_369
timestamp 1676037725
transform 1 0 35052 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_373
timestamp 1676037725
transform 1 0 35420 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_404
timestamp 1676037725
transform 1 0 38272 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_424
timestamp 1676037725
transform 1 0 40112 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_446
timestamp 1676037725
transform 1 0 42136 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_525
timestamp 1676037725
transform 1 0 49404 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_223
timestamp 1676037725
transform 1 0 21620 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_236
timestamp 1676037725
transform 1 0 22816 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1676037725
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_275
timestamp 1676037725
transform 1 0 26404 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_287
timestamp 1676037725
transform 1 0 27508 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_299
timestamp 1676037725
transform 1 0 28612 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_315
timestamp 1676037725
transform 1 0 30084 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_336
timestamp 1676037725
transform 1 0 32016 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_342
timestamp 1676037725
transform 1 0 32568 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_352
timestamp 1676037725
transform 1 0 33488 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_362
timestamp 1676037725
transform 1 0 34408 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_371
timestamp 1676037725
transform 1 0 35236 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_374
timestamp 1676037725
transform 1 0 35512 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_378
timestamp 1676037725
transform 1 0 35880 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_399
timestamp 1676037725
transform 1 0 37812 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_407
timestamp 1676037725
transform 1 0 38548 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_418
timestamp 1676037725
transform 1 0 39560 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_454
timestamp 1676037725
transform 1 0 42872 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_466
timestamp 1676037725
transform 1 0 43976 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_474
timestamp 1676037725
transform 1 0 44712 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_260
timestamp 1676037725
transform 1 0 25024 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_272
timestamp 1676037725
transform 1 0 26128 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_314
timestamp 1676037725
transform 1 0 29992 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_326
timestamp 1676037725
transform 1 0 31096 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_334
timestamp 1676037725
transform 1 0 31832 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_359
timestamp 1676037725
transform 1 0 34132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1676037725
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_427
timestamp 1676037725
transform 1 0 40388 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_440
timestamp 1676037725
transform 1 0 41584 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_513
timestamp 1676037725
transform 1 0 48300 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_525
timestamp 1676037725
transform 1 0 49404 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_239
timestamp 1676037725
transform 1 0 23092 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_249
timestamp 1676037725
transform 1 0 24012 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_274
timestamp 1676037725
transform 1 0 26312 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_287
timestamp 1676037725
transform 1 0 27508 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 1676037725
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1676037725
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_331
timestamp 1676037725
transform 1 0 31556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_337
timestamp 1676037725
transform 1 0 32108 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_347
timestamp 1676037725
transform 1 0 33028 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_362
timestamp 1676037725
transform 1 0 34408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_380
timestamp 1676037725
transform 1 0 36064 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_392
timestamp 1676037725
transform 1 0 37168 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_404
timestamp 1676037725
transform 1 0 38272 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_408
timestamp 1676037725
transform 1 0 38640 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_418
timestamp 1676037725
transform 1 0 39560 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1676037725
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1676037725
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1676037725
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_47
timestamp 1676037725
transform 1 0 5428 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_97
timestamp 1676037725
transform 1 0 10028 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_107
timestamp 1676037725
transform 1 0 10948 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1676037725
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_236
timestamp 1676037725
transform 1 0 22816 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_242
timestamp 1676037725
transform 1 0 23368 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_254
timestamp 1676037725
transform 1 0 24472 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_277
timestamp 1676037725
transform 1 0 26588 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_304
timestamp 1676037725
transform 1 0 29072 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1676037725
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1676037725
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_345
timestamp 1676037725
transform 1 0 32844 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_368
timestamp 1676037725
transform 1 0 34960 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_380
timestamp 1676037725
transform 1 0 36064 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_401
timestamp 1676037725
transform 1 0 37996 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_423
timestamp 1676037725
transform 1 0 40020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_435
timestamp 1676037725
transform 1 0 41124 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_513
timestamp 1676037725
transform 1 0 48300 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_525
timestamp 1676037725
transform 1 0 49404 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_9
timestamp 1676037725
transform 1 0 1932 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1676037725
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_219
timestamp 1676037725
transform 1 0 21252 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_246
timestamp 1676037725
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1676037725
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_277
timestamp 1676037725
transform 1 0 26588 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_290
timestamp 1676037725
transform 1 0 27784 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_302
timestamp 1676037725
transform 1 0 28888 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_321
timestamp 1676037725
transform 1 0 30636 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_349
timestamp 1676037725
transform 1 0 33212 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 1676037725
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_387
timestamp 1676037725
transform 1 0 36708 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_411
timestamp 1676037725
transform 1 0 38916 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_525
timestamp 1676037725
transform 1 0 49404 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_63
timestamp 1676037725
transform 1 0 6900 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_68
timestamp 1676037725
transform 1 0 7360 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_76
timestamp 1676037725
transform 1 0 8096 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_88
timestamp 1676037725
transform 1 0 9200 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_100
timestamp 1676037725
transform 1 0 10304 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_216
timestamp 1676037725
transform 1 0 20976 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_231
timestamp 1676037725
transform 1 0 22356 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_243
timestamp 1676037725
transform 1 0 23460 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_270
timestamp 1676037725
transform 1 0 25944 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1676037725
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_310
timestamp 1676037725
transform 1 0 29624 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1676037725
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_355
timestamp 1676037725
transform 1 0 33764 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_376
timestamp 1676037725
transform 1 0 35696 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_388
timestamp 1676037725
transform 1 0 36800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_401
timestamp 1676037725
transform 1 0 37996 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_424
timestamp 1676037725
transform 1 0 40112 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_445
timestamp 1676037725
transform 1 0 42044 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_513
timestamp 1676037725
transform 1 0 48300 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_525
timestamp 1676037725
transform 1 0 49404 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_91
timestamp 1676037725
transform 1 0 9476 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_103
timestamp 1676037725
transform 1 0 10580 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_115
timestamp 1676037725
transform 1 0 11684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_127
timestamp 1676037725
transform 1 0 12788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_173
timestamp 1676037725
transform 1 0 17020 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_178
timestamp 1676037725
transform 1 0 17480 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_190
timestamp 1676037725
transform 1 0 18584 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_286
timestamp 1676037725
transform 1 0 27416 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_298
timestamp 1676037725
transform 1 0 28520 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1676037725
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1676037725
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1676037725
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1676037725
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1676037725
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1676037725
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_373
timestamp 1676037725
transform 1 0 35420 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_395
timestamp 1676037725
transform 1 0 37444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_407
timestamp 1676037725
transform 1 0 38548 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1676037725
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_432
timestamp 1676037725
transform 1 0 40848 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_444
timestamp 1676037725
transform 1 0 41952 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_456
timestamp 1676037725
transform 1 0 43056 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_468
timestamp 1676037725
transform 1 0 44160 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1676037725
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1676037725
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_117
timestamp 1676037725
transform 1 0 11868 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_122
timestamp 1676037725
transform 1 0 12328 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_134
timestamp 1676037725
transform 1 0 13432 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_146
timestamp 1676037725
transform 1 0 14536 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_158
timestamp 1676037725
transform 1 0 15640 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1676037725
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_174
timestamp 1676037725
transform 1 0 17112 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_186
timestamp 1676037725
transform 1 0 18216 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_198
timestamp 1676037725
transform 1 0 19320 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_206
timestamp 1676037725
transform 1 0 20056 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_211
timestamp 1676037725
transform 1 0 20516 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_218
timestamp 1676037725
transform 1 0 21160 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_261
timestamp 1676037725
transform 1 0 25116 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_278
timestamp 1676037725
transform 1 0 26680 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_293
timestamp 1676037725
transform 1 0 28060 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_321
timestamp 1676037725
transform 1 0 30636 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_333
timestamp 1676037725
transform 1 0 31740 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_359
timestamp 1676037725
transform 1 0 34132 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_383
timestamp 1676037725
transform 1 0 36340 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1676037725
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_430
timestamp 1676037725
transform 1 0 40664 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_442
timestamp 1676037725
transform 1 0 41768 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_513
timestamp 1676037725
transform 1 0 48300 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_525
timestamp 1676037725
transform 1 0 49404 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_117
timestamp 1676037725
transform 1 0 11868 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_123
timestamp 1676037725
transform 1 0 12420 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_131
timestamp 1676037725
transform 1 0 13156 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_137
timestamp 1676037725
transform 1 0 13708 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_158
timestamp 1676037725
transform 1 0 15640 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_166
timestamp 1676037725
transform 1 0 16376 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_174
timestamp 1676037725
transform 1 0 17112 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_186
timestamp 1676037725
transform 1 0 18216 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_194
timestamp 1676037725
transform 1 0 18952 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_201
timestamp 1676037725
transform 1 0 19596 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_204
timestamp 1676037725
transform 1 0 19872 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_212
timestamp 1676037725
transform 1 0 20608 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_216
timestamp 1676037725
transform 1 0 20976 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_228
timestamp 1676037725
transform 1 0 22080 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_238
timestamp 1676037725
transform 1 0 23000 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1676037725
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1676037725
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1676037725
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_289
timestamp 1676037725
transform 1 0 27692 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1676037725
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_313
timestamp 1676037725
transform 1 0 29900 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_334
timestamp 1676037725
transform 1 0 31832 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_358
timestamp 1676037725
transform 1 0 34040 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1676037725
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_389
timestamp 1676037725
transform 1 0 36892 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_402
timestamp 1676037725
transform 1 0 38088 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_414
timestamp 1676037725
transform 1 0 39192 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1676037725
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1676037725
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1676037725
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1676037725
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1676037725
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1676037725
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_141
timestamp 1676037725
transform 1 0 14076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_146
timestamp 1676037725
transform 1 0 14536 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_158
timestamp 1676037725
transform 1 0 15640 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_166
timestamp 1676037725
transform 1 0 16376 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1676037725
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1676037725
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1676037725
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1676037725
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1676037725
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1676037725
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1676037725
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1676037725
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1676037725
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_373
timestamp 1676037725
transform 1 0 35420 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_390
timestamp 1676037725
transform 1 0 36984 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_405
timestamp 1676037725
transform 1 0 38364 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_418
timestamp 1676037725
transform 1 0 39560 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_430
timestamp 1676037725
transform 1 0 40664 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_442
timestamp 1676037725
transform 1 0 41768 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_525
timestamp 1676037725
transform 1 0 49404 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_240
timestamp 1676037725
transform 1 0 23184 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_259
timestamp 1676037725
transform 1 0 24932 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_263
timestamp 1676037725
transform 1 0 25300 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_275
timestamp 1676037725
transform 1 0 26404 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_287
timestamp 1676037725
transform 1 0 27508 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_299
timestamp 1676037725
transform 1 0 28612 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1676037725
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1676037725
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1676037725
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1676037725
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1676037725
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_376
timestamp 1676037725
transform 1 0 35696 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_388
timestamp 1676037725
transform 1 0 36800 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_400
timestamp 1676037725
transform 1 0 37904 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_412
timestamp 1676037725
transform 1 0 39008 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_525
timestamp 1676037725
transform 1 0 49404 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_153
timestamp 1676037725
transform 1 0 15180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1676037725
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1676037725
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1676037725
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1676037725
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1676037725
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1676037725
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1676037725
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1676037725
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_348
timestamp 1676037725
transform 1 0 33120 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1676037725
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1676037725
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1676037725
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1676037725
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1676037725
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1676037725
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1676037725
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1676037725
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1676037725
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1676037725
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_519
timestamp 1676037725
transform 1 0 48852 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_9
timestamp 1676037725
transform 1 0 1932 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1676037725
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_177
timestamp 1676037725
transform 1 0 17388 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_185
timestamp 1676037725
transform 1 0 18124 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_191
timestamp 1676037725
transform 1 0 18676 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1676037725
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_203
timestamp 1676037725
transform 1 0 19780 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_215
timestamp 1676037725
transform 1 0 20884 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_227
timestamp 1676037725
transform 1 0 21988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_239
timestamp 1676037725
transform 1 0 23092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1676037725
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_277
timestamp 1676037725
transform 1 0 26588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_281
timestamp 1676037725
transform 1 0 26956 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_293
timestamp 1676037725
transform 1 0 28060 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_305
timestamp 1676037725
transform 1 0 29164 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1676037725
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1676037725
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1676037725
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1676037725
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1676037725
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1676037725
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1676037725
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1676037725
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1676037725
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1676037725
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1676037725
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1676037725
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1676037725
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1676037725
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1676037725
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1676037725
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1676037725
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1676037725
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1676037725
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1676037725
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1676037725
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1676037725
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1676037725
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_525
timestamp 1676037725
transform 1 0 49404 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1676037725
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1676037725
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1676037725
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1676037725
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1676037725
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1676037725
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1676037725
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1676037725
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1676037725
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1676037725
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1676037725
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_525
timestamp 1676037725
transform 1 0 49404 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_258
timestamp 1676037725
transform 1 0 24840 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_270
timestamp 1676037725
transform 1 0 25944 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_278
timestamp 1676037725
transform 1 0 26680 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1676037725
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1676037725
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1676037725
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1676037725
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1676037725
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1676037725
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1676037725
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1676037725
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1676037725
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1676037725
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1676037725
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1676037725
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1676037725
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1676037725
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_525
timestamp 1676037725
transform 1 0 49404 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1676037725
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1676037725
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1676037725
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1676037725
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1676037725
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1676037725
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1676037725
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1676037725
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1676037725
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1676037725
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1676037725
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1676037725
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1676037725
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1676037725
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_513
timestamp 1676037725
transform 1 0 48300 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_525
timestamp 1676037725
transform 1 0 49404 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1676037725
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1676037725
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1676037725
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1676037725
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1676037725
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1676037725
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1676037725
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1676037725
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_525
timestamp 1676037725
transform 1 0 49404 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1676037725
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_86_187
timestamp 1676037725
transform 1 0 18308 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_205
timestamp 1676037725
transform 1 0 19964 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_211
timestamp 1676037725
transform 1 0 20516 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_223
timestamp 1676037725
transform 1 0 21620 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_235
timestamp 1676037725
transform 1 0 22724 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_247
timestamp 1676037725
transform 1 0 23828 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1676037725
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1676037725
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1676037725
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1676037725
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1676037725
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1676037725
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1676037725
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1676037725
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1676037725
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1676037725
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1676037725
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1676037725
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1676037725
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1676037725
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1676037725
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1676037725
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1676037725
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1676037725
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1676037725
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_119
timestamp 1676037725
transform 1 0 12052 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_124
timestamp 1676037725
transform 1 0 12512 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_136
timestamp 1676037725
transform 1 0 13616 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_144
timestamp 1676037725
transform 1 0 14352 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_150
timestamp 1676037725
transform 1 0 14904 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_162
timestamp 1676037725
transform 1 0 16008 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1676037725
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1676037725
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1676037725
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1676037725
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1676037725
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1676037725
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1676037725
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1676037725
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1676037725
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1676037725
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1676037725
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1676037725
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1676037725
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1676037725
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1676037725
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_525
timestamp 1676037725
transform 1 0 49404 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1676037725
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1676037725
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_205
timestamp 1676037725
transform 1 0 19964 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_210
timestamp 1676037725
transform 1 0 20424 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_222
timestamp 1676037725
transform 1 0 21528 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_234
timestamp 1676037725
transform 1 0 22632 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_246
timestamp 1676037725
transform 1 0 23736 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1676037725
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1676037725
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1676037725
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1676037725
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1676037725
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_513
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_525
timestamp 1676037725
transform 1 0 49404 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_9
timestamp 1676037725
transform 1 0 1932 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_21
timestamp 1676037725
transform 1 0 3036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_33
timestamp 1676037725
transform 1 0 4140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_45
timestamp 1676037725
transform 1 0 5244 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_53
timestamp 1676037725
transform 1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_89_231
timestamp 1676037725
transform 1 0 22356 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_242
timestamp 1676037725
transform 1 0 23368 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_254
timestamp 1676037725
transform 1 0 24472 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_266
timestamp 1676037725
transform 1 0 25576 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_278
timestamp 1676037725
transform 1 0 26680 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1676037725
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1676037725
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1676037725
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1676037725
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1676037725
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1676037725
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1676037725
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1676037725
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1676037725
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_517
timestamp 1676037725
transform 1 0 48668 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_525
timestamp 1676037725
transform 1 0 49404 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1676037725
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1676037725
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_127
timestamp 1676037725
transform 1 0 12788 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_132
timestamp 1676037725
transform 1 0 13248 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_147
timestamp 1676037725
transform 1 0 14628 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_159
timestamp 1676037725
transform 1 0 15732 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_171
timestamp 1676037725
transform 1 0 16836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_183
timestamp 1676037725
transform 1 0 17940 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_259
timestamp 1676037725
transform 1 0 24932 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_271
timestamp 1676037725
transform 1 0 26036 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_283
timestamp 1676037725
transform 1 0 27140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_295
timestamp 1676037725
transform 1 0 28244 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1676037725
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1676037725
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1676037725
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1676037725
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1676037725
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1676037725
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1676037725
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1676037725
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_513
timestamp 1676037725
transform 1 0 48300 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_525
timestamp 1676037725
transform 1 0 49404 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_21
timestamp 1676037725
transform 1 0 3036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_33
timestamp 1676037725
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1676037725
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1676037725
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1676037725
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1676037725
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_243
timestamp 1676037725
transform 1 0 23460 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_247
timestamp 1676037725
transform 1 0 23828 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_259
timestamp 1676037725
transform 1 0 24932 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_271
timestamp 1676037725
transform 1 0 26036 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_517
timestamp 1676037725
transform 1 0 48668 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_525
timestamp 1676037725
transform 1 0 49404 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_21
timestamp 1676037725
transform 1 0 3036 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_49
timestamp 1676037725
transform 1 0 5612 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_61
timestamp 1676037725
transform 1 0 6716 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_73
timestamp 1676037725
transform 1 0 7820 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_81
timestamp 1676037725
transform 1 0 8556 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_105
timestamp 1676037725
transform 1 0 10764 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_117
timestamp 1676037725
transform 1 0 11868 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_129
timestamp 1676037725
transform 1 0 12972 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_137
timestamp 1676037725
transform 1 0 13708 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_161
timestamp 1676037725
transform 1 0 15916 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_173
timestamp 1676037725
transform 1 0 17020 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_185
timestamp 1676037725
transform 1 0 18124 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_193
timestamp 1676037725
transform 1 0 18860 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1676037725
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1676037725
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1676037725
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1676037725
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1676037725
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1676037725
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1676037725
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1676037725
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1676037725
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1676037725
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_525
timestamp 1676037725
transform 1 0 49404 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_9
timestamp 1676037725
transform 1 0 1932 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_33
timestamp 1676037725
transform 1 0 4140 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_37
timestamp 1676037725
transform 1 0 4508 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1676037725
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_89
timestamp 1676037725
transform 1 0 9292 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1676037725
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_145
timestamp 1676037725
transform 1 0 14444 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_166
timestamp 1676037725
transform 1 0 16376 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1676037725
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1676037725
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1676037725
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1676037725
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_489
timestamp 1676037725
transform 1 0 46092 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_493
timestamp 1676037725
transform 1 0 46460 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_501
timestamp 1676037725
transform 1 0 47196 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_525
timestamp 1676037725
transform 1 0 49404 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_94_25
timestamp 1676037725
transform 1 0 3404 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_61
timestamp 1676037725
transform 1 0 6716 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_81
timestamp 1676037725
transform 1 0 8556 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_117
timestamp 1676037725
transform 1 0 11868 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_137
timestamp 1676037725
transform 1 0 13708 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_157
timestamp 1676037725
transform 1 0 15548 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_174
timestamp 1676037725
transform 1 0 17112 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_194
timestamp 1676037725
transform 1 0 18952 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_241
timestamp 1676037725
transform 1 0 23276 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_248
timestamp 1676037725
transform 1 0 23920 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_259
timestamp 1676037725
transform 1 0 24932 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_271
timestamp 1676037725
transform 1 0 26036 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_283
timestamp 1676037725
transform 1 0 27140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_295
timestamp 1676037725
transform 1 0 28244 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1676037725
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_314
timestamp 1676037725
transform 1 0 29992 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_326
timestamp 1676037725
transform 1 0 31096 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_334
timestamp 1676037725
transform 1 0 31832 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_340
timestamp 1676037725
transform 1 0 32384 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_352
timestamp 1676037725
transform 1 0 33488 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_372
timestamp 1676037725
transform 1 0 35328 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_384
timestamp 1676037725
transform 1 0 36432 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_396
timestamp 1676037725
transform 1 0 37536 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_400
timestamp 1676037725
transform 1 0 37904 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_404
timestamp 1676037725
transform 1 0 38272 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_416
timestamp 1676037725
transform 1 0 39376 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_433
timestamp 1676037725
transform 1 0 40940 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_444
timestamp 1676037725
transform 1 0 41952 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_456
timestamp 1676037725
transform 1 0 43056 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_468
timestamp 1676037725
transform 1 0 44160 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_525
timestamp 1676037725
transform 1 0 49404 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_34
timestamp 1676037725
transform 1 0 4232 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1676037725
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_121
timestamp 1676037725
transform 1 0 12236 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1676037725
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_149
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_166
timestamp 1676037725
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_177
timestamp 1676037725
transform 1 0 17388 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_194
timestamp 1676037725
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_222
timestamp 1676037725
transform 1 0 21528 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_249
timestamp 1676037725
transform 1 0 24012 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_261
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_269
timestamp 1676037725
transform 1 0 25852 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_276
timestamp 1676037725
transform 1 0 26496 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_287
timestamp 1676037725
transform 1 0 27508 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_295
timestamp 1676037725
transform 1 0 28244 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_303
timestamp 1676037725
transform 1 0 28980 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_307
timestamp 1676037725
transform 1 0 29348 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_309
timestamp 1676037725
transform 1 0 29532 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_317
timestamp 1676037725
transform 1 0 30268 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_325
timestamp 1676037725
transform 1 0 31004 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_333
timestamp 1676037725
transform 1 0 31740 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_349
timestamp 1676037725
transform 1 0 33212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_357
timestamp 1676037725
transform 1 0 33948 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_363
timestamp 1676037725
transform 1 0 34500 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_365
timestamp 1676037725
transform 1 0 34684 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_371
timestamp 1676037725
transform 1 0 35236 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_381
timestamp 1676037725
transform 1 0 36156 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_389
timestamp 1676037725
transform 1 0 36892 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_399
timestamp 1676037725
transform 1 0 37812 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_407
timestamp 1676037725
transform 1 0 38548 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_413
timestamp 1676037725
transform 1 0 39100 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_419
timestamp 1676037725
transform 1 0 39652 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_421
timestamp 1676037725
transform 1 0 39836 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_427
timestamp 1676037725
transform 1 0 40388 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_435
timestamp 1676037725
transform 1 0 41124 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_442
timestamp 1676037725
transform 1 0 41768 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_457
timestamp 1676037725
transform 1 0 43148 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_464
timestamp 1676037725
transform 1 0 43792 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_471
timestamp 1676037725
transform 1 0 44436 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_475
timestamp 1676037725
transform 1 0 44804 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_477
timestamp 1676037725
transform 1 0 44988 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_482
timestamp 1676037725
transform 1 0 45448 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_494
timestamp 1676037725
transform 1 0 46552 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_502
timestamp 1676037725
transform 1 0 47288 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_525
timestamp 1676037725
transform 1 0 49404 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 3956 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 49128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 48484 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 49128 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 49128 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 49128 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 49128 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 49128 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 49128 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1676037725
transform 1 0 48484 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 49128 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 49128 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1676037725
transform 1 0 48484 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 48484 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform 1 0 48484 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1676037725
transform 1 0 48484 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 48484 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1676037725
transform 1 0 48484 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform 1 0 48484 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform 1 0 48484 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1676037725
transform 1 0 48484 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1676037725
transform 1 0 48484 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 47932 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1676037725
transform 1 0 48484 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1676037725
transform 1 0 48484 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 49128 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 49128 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1676037725
transform 1 0 48484 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 49128 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform 1 0 48484 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform 1 0 48484 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input35
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1676037725
transform 1 0 10672 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input39
timestamp 1676037725
transform 1 0 11868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input41
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1676037725
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input46
timestamp 1676037725
transform 1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input47
timestamp 1676037725
transform 1 0 17020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1676037725
transform 1 0 19228 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input51
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1676037725
transform 1 0 20608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1676037725
transform 1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1676037725
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1676037725
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input60
timestamp 1676037725
transform 1 0 5520 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1676037725
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1676037725
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 23644 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1676037725
transform 1 0 30636 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1676037725
transform 1 0 31372 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 32108 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 32844 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 33580 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1676037725
transform 1 0 34868 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 35052 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 35788 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 36524 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 37444 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 24564 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1676037725
transform 1 0 37996 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 38732 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 40020 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 40756 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 41492 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 41676 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input81
timestamp 1676037725
transform 1 0 42596 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 43516 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 44160 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 45172 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1676037725
transform 1 0 24748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1676037725
transform 1 0 25484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 26220 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1676037725
transform 1 0 27140 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1676037725
transform 1 0 27876 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1676037725
transform 1 0 28612 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 29716 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1676037725
transform 1 0 29900 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 1564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 1564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 1564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1676037725
transform 1 0 45448 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1676037725
transform 1 0 46368 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1676037725
transform 1 0 49036 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1676037725
transform 1 0 49036 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1676037725
transform 1 0 49036 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform 1 0 49036 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1676037725
transform 1 0 49036 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input105
timestamp 1676037725
transform 1 0 48852 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform 1 0 49036 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input107
timestamp 1676037725
transform 1 0 49036 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input108
timestamp 1676037725
transform 1 0 48484 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input111
timestamp 1676037725
transform 1 0 1564 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1676037725
transform 1 0 1564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  left_tile_264
timestamp 1676037725
transform 1 0 49128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output113 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 1564 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 47932 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 47932 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 47932 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 47932 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 47932 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 47932 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 47932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 47932 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 47932 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 47932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 47932 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 47932 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 47932 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 47932 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 31556 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 34132 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 33948 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 34868 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 36708 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 23276 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 39284 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 39100 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 40020 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 41860 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 42596 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 44436 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 25208 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 27324 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 29716 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 1564 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform 1 0 9292 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 10396 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform 1 0 12972 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 14444 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform 1 0 14904 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform 1 0 1932 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 15640 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform 1 0 14904 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform 1 0 17388 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform 1 0 17480 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 17480 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 19596 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform 1 0 19964 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 20056 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform 1 0 21804 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 22540 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 2668 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 4140 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 5244 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 7084 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform 1 0 7820 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output211
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output212
timestamp 1676037725
transform 1 0 47748 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output213
timestamp 1676037725
transform 1 0 47932 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output214
timestamp 1676037725
transform 1 0 46828 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output215
timestamp 1676037725
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output216
timestamp 1676037725
transform 1 0 47932 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output217
timestamp 1676037725
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output218
timestamp 1676037725
transform 1 0 47932 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 49864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 49864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 49864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 49864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 49864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 49864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 49864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 49864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 49864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 49864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 49864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 49864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 49864 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 49864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 49864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 49864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 49864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 49864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 49864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 49864 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 49864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 49864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 49864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 49864 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 49864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 49864 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 49864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 49864 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 49864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 49864 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 49864 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 49864 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 49864 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 49864 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 49864 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 49864 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 49864 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 49864 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 49864 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 49864 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 49864 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 49864 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 49864 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 49864 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 49864 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 49864 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 49864 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 49864 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 49864 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 49864 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 49864 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 49864 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 49864 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 49864 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 49864 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33672 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30084 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29808 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32476 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35328 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38732 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 38456 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37536 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34960 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33948 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32200 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34224 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 36984 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37720 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40296 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 40296 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 36432 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33948 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34500 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32476 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 31280 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 36248 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40296 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 39284 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34040 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21620 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33948 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38732 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 41860 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 42596 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 42688 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 42136 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38548 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 38088 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 39744 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40296 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 41492 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38180 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 38548 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 38272 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35972 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37076 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35604 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34684 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34868 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33856 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33120 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34500 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 31372 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32200 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29992 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28796 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28152 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 28244 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27232 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26220 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 27048 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27692 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27968 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28520 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28428 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29348 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27140 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25944 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24932 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24656 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22448 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19228 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22448 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25852 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28796 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30636 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34500 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35512 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37720 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33672 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33856 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10120 0 1 47872
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24104 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 25576 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27692 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30176 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29716 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29072 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 26772 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24656 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23092 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23368 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21712 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20516 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23000 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23828 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22264 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22816 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21068 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19504 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24564 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23184 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24748 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27232 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34408 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32200 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31740 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35512 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 25576 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32016 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__269
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28612 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30268 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33028 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 37444 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33488 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__219
timestamp 1676037725
transform 1 0 31464 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 29992 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32384 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 35972 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40940 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38732 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__222
timestamp 1676037725
transform 1 0 40020 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38180 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37812 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36064 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38640 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__224
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1676037725
transform 1 0 31004 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35144 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33672 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32936 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38364 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 32292 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__270
timestamp 1676037725
transform 1 0 29716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 27600 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 31004 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32476 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33672 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40388 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 34868 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__271
timestamp 1676037725
transform 1 0 36708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36524 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 34868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34960 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41584 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 37444 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__272
timestamp 1676037725
transform 1 0 40020 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40112 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 37444 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35420 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__273
timestamp 1676037725
transform 1 0 36156 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36064 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38180 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34684 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 29716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27600 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30820 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27968 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40756 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 41676 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 42596 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 42596 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 38732 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 35604 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__223
timestamp 1676037725
transform 1 0 31556 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32016 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37904 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38180 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__225
timestamp 1676037725
transform 1 0 38456 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38640 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 40756 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 43976 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 41216 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40296 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 37444 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 41860 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__231
timestamp 1676037725
transform 1 0 41768 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 41308 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 42964 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 45448 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38548 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__242
timestamp 1676037725
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34868 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 38916 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 43056 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 39836 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 36248 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40756 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__251
timestamp 1676037725
transform 1 0 41216 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 40112 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 44804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 38732 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 39284 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1676037725
transform 1 0 34408 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38732 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38456 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__252
timestamp 1676037725
transform 1 0 39008 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 38732 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 43608 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37260 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 36984 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__226
timestamp 1676037725
transform 1 0 31924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30728 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41308 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 36156 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36340 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__227
timestamp 1676037725
transform 1 0 31556 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36248 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41952 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35512 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__228
timestamp 1676037725
transform 1 0 33672 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35052 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40664 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__229
timestamp 1676037725
transform 1 0 28980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33672 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39284 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32200 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27140 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__230
timestamp 1676037725
transform 1 0 27416 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33672 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37536 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28428 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32108 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 28612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27232 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 26680 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29900 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 26496 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25300 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__234
timestamp 1676037725
transform 1 0 27140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30728 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37444 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31924 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__235
timestamp 1676037725
transform 1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25484 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30820 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37628 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__236
timestamp 1676037725
transform 1 0 24564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29624 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30176 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26220 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__237
timestamp 1676037725
transform 1 0 25208 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29900 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__238
timestamp 1676037725
transform 1 0 24932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23736 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28336 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 35788 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__239
timestamp 1676037725
transform 1 0 23184 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22724 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27784 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 35052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__240
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 30360 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25300 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 30636 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29808 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__243
timestamp 1676037725
transform 1 0 32016 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29808 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__244
timestamp 1676037725
transform 1 0 34776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33028 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31004 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__245
timestamp 1676037725
transform 1 0 35972 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34776 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33304 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__246
timestamp 1676037725
transform 1 0 37904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41768 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 38640 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__247
timestamp 1676037725
transform 1 0 34132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__248
timestamp 1676037725
transform 1 0 38364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37168 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41492 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32660 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__249
timestamp 1676037725
transform 1 0 36340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40664 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33580 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__250
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35236 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 31004 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__253
timestamp 1676037725
transform 1 0 22724 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 23276 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 26956 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25852 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38548 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32660 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__256
timestamp 1676037725
transform 1 0 29992 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30912 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29440 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 26680 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32384 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38824 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 25576 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__260
timestamp 1676037725
transform 1 0 27140 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 26036 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 27324 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 25024 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 37444 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 30452 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1676037725
transform 1 0 21988 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__263
timestamp 1676037725
transform 1 0 22632 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27048 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25300 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24472 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22908 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35604 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28336 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__254
timestamp 1676037725
transform 1 0 21252 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25024 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21804 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 36340 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28428 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__255
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23460 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22080 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31004 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 37352 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 22172 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__257
timestamp 1676037725
transform 1 0 23368 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20700 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27784 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28428 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__258
timestamp 1676037725
transform 1 0 18400 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17204 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28520 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28428 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__259
timestamp 1676037725
transform 1 0 22448 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22080 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23184 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18400 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__261
timestamp 1676037725
transform 1 0 24564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19504 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37352 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__262
timestamp 1676037725
transform 1 0 29716 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28704 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29900 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20884 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 29440 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 34592 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 39744 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 44896 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 54952 800 55072 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 386 56200 442 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 50200 25304 51000 25424 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 50200 32104 51000 32224 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 50200 32784 51000 32904 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 50200 33464 51000 33584 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 50200 34144 51000 34264 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 50200 34824 51000 34944 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 50200 35504 51000 35624 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 50200 36184 51000 36304 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 50200 36864 51000 36984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 50200 37544 51000 37664 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 50200 38224 51000 38344 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 50200 25984 51000 26104 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 50200 38904 51000 39024 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 50200 39584 51000 39704 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 50200 40264 51000 40384 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 50200 40944 51000 41064 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 50200 41624 51000 41744 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 50200 42304 51000 42424 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 50200 42984 51000 43104 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 50200 43664 51000 43784 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 50200 44344 51000 44464 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 50200 45024 51000 45144 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 50200 26664 51000 26784 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 50200 27344 51000 27464 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 50200 28024 51000 28144 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 50200 28704 51000 28824 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 50200 29384 51000 29504 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 50200 30064 51000 30184 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 50200 30744 51000 30864 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 50200 31424 51000 31544 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 50200 4904 51000 5024 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 50200 11704 51000 11824 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 50200 13064 51000 13184 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 50200 13744 51000 13864 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 50200 15104 51000 15224 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 50200 15784 51000 15904 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 50200 17144 51000 17264 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 50200 17824 51000 17944 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 50200 5584 51000 5704 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 50200 19184 51000 19304 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 50200 19864 51000 19984 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 50200 21224 51000 21344 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 50200 23264 51000 23384 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 50200 23944 51000 24064 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 50200 6944 51000 7064 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 50200 7624 51000 7744 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 50200 8984 51000 9104 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 50200 9664 51000 9784 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 50200 11024 51000 11144 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 23202 56200 23258 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 30562 56200 30618 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 31298 56200 31354 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 32034 56200 32090 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 32770 56200 32826 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 33506 56200 33562 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 34242 56200 34298 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 34978 56200 35034 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 35714 56200 35770 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 36450 56200 36506 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 37186 56200 37242 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 23938 56200 23994 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 37922 56200 37978 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 38658 56200 38714 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 39394 56200 39450 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 40130 56200 40186 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 40866 56200 40922 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 41602 56200 41658 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 42338 56200 42394 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 43074 56200 43130 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 43810 56200 43866 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 44546 56200 44602 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 24674 56200 24730 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 25410 56200 25466 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 26146 56200 26202 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 26882 56200 26938 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 27618 56200 27674 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 28354 56200 28410 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 29090 56200 29146 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 29826 56200 29882 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1122 56200 1178 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 8482 56200 8538 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 9218 56200 9274 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 11426 56200 11482 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 12162 56200 12218 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 12898 56200 12954 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 13634 56200 13690 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 14370 56200 14426 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 1858 56200 1914 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 15842 56200 15898 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 16578 56200 16634 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 17314 56200 17370 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 18050 56200 18106 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 18786 56200 18842 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 19522 56200 19578 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 20994 56200 21050 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 22466 56200 22522 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2594 56200 2650 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 3330 56200 3386 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 4066 56200 4122 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 5538 56200 5594 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 6274 56200 6330 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 7010 56200 7066 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 7746 56200 7802 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 31832 800 31952 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 36456 800 36576 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 24896 800 25016 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 prog_reset_bottom_in
port 200 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 prog_reset_bottom_out
port 201 nsew signal tristate
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 prog_reset_left_in
port 202 nsew signal input
flabel metal3 s 50200 45704 51000 45824 0 FreeSans 480 0 0 0 prog_reset_right_out
port 203 nsew signal tristate
flabel metal2 s 47490 56200 47546 57000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 204 nsew signal input
flabel metal2 s 46754 56200 46810 57000 0 FreeSans 224 90 0 0 prog_reset_top_out
port 205 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 reset_bottom_in
port 206 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 reset_bottom_out
port 207 nsew signal tristate
flabel metal3 s 50200 46384 51000 46504 0 FreeSans 480 0 0 0 reset_right_in
port 208 nsew signal input
flabel metal2 s 48962 56200 49018 57000 0 FreeSans 224 90 0 0 reset_top_in
port 209 nsew signal input
flabel metal2 s 48226 56200 48282 57000 0 FreeSans 224 90 0 0 reset_top_out
port 210 nsew signal tristate
flabel metal3 s 50200 47064 51000 47184 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 211 nsew signal input
flabel metal3 s 50200 47744 51000 47864 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 212 nsew signal input
flabel metal3 s 50200 48424 51000 48544 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 213 nsew signal input
flabel metal3 s 50200 49104 51000 49224 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 214 nsew signal input
flabel metal3 s 50200 49784 51000 49904 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 215 nsew signal input
flabel metal3 s 50200 50464 51000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 216 nsew signal input
flabel metal3 s 50200 51144 51000 51264 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 217 nsew signal input
flabel metal3 s 50200 51824 51000 51944 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 218 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 219 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 220 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 221 nsew signal tristate
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 222 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 test_enable_bottom_in
port 223 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 test_enable_bottom_out
port 224 nsew signal tristate
flabel metal3 s 50200 52504 51000 52624 0 FreeSans 480 0 0 0 test_enable_right_in
port 225 nsew signal input
flabel metal2 s 50434 56200 50490 57000 0 FreeSans 224 90 0 0 test_enable_top_in
port 226 nsew signal input
flabel metal2 s 49698 56200 49754 57000 0 FreeSans 224 90 0 0 test_enable_top_out
port 227 nsew signal tristate
flabel metal3 s 0 45704 800 45824 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 228 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 229 nsew signal input
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 230 nsew signal input
flabel metal3 s 0 52640 800 52760 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 231 nsew signal input
rlabel metal1 25484 54400 25484 54400 0 VGND
rlabel metal1 25484 53856 25484 53856 0 VPWR
rlabel metal1 17986 22576 17986 22576 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal1 10028 26418 10028 26418 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 13248 21658 13248 21658 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 12650 20026 12650 20026 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 11592 21522 11592 21522 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20010 23596 20010 23596 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal2 21574 13838 21574 13838 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal2 21114 23120 21114 23120 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal2 21298 24174 21298 24174 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 21436 19686 21436 19686 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 29026 17136 29026 17136 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal2 20562 18870 20562 18870 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal2 21298 19482 21298 19482 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 21206 17714 21206 17714 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal2 25070 17476 25070 17476 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal2 21942 18496 21942 18496 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 21298 18156 21298 18156 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 27738 18190 27738 18190 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 24978 18802 24978 18802 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 20010 22610 20010 22610 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal2 26542 17680 26542 17680 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20240 23834 20240 23834 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 17940 23834 17940 23834 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 27370 18802 27370 18802 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28382 18632 28382 18632 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25714 21658 25714 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23414 19278 23414 19278 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 25116 20026 25116 20026 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24380 21658 24380 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21068 23630 21068 23630 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 23322 24480 23322 24480 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 19826 23562 19826 23562 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 28796 12954 28796 12954 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20332 19482 20332 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 16054 20468 16054 20468 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 28014 16558 28014 16558 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26220 20570 26220 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 26680 18938 26680 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22770 19584 22770 19584 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 26772 16422 26772 16422 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24288 18734 24288 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 20010 17850 20010 17850 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 21252 19482 21252 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 21022 19142 21022 19142 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 29532 12682 29532 12682 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20286 18394 20286 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 15686 18938 15686 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 27968 13498 27968 13498 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27462 21862 27462 21862 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 26818 17306 26818 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21206 21488 21206 21488 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 25898 16014 25898 16014 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 25208 17306 25208 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 21206 19312 21206 19312 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 22862 17782 22862 17782 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 21298 17680 21298 17680 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 27186 17442 27186 17442 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18630 22746 18630 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 15134 22066 15134 22066 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 26174 18394 26174 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 26818 20978 26818 20978 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23782 21930 23782 21930 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20240 18938 20240 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24012 18938 24012 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 23322 22406 23322 22406 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 19688 21114 19688 21114 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 22310 23936 22310 23936 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 19320 22474 19320 22474 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 10810 25398 10810 25398 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 4554 23086 4554 23086 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 5957 28050 5957 28050 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 7751 27574 7751 27574 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 14122 23970 14122 23970 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 8464 23630 8464 23630 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 6026 24548 6026 24548 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 7843 26554 7843 26554 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 16606 19006 16606 19006 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 9338 19822 9338 19822 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 9706 22066 9706 22066 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 8441 24718 8441 24718 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 9798 20162 9798 20162 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 10258 21794 10258 21794 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 9177 23154 9177 23154 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal3 1740 55012 1740 55012 0 ccff_head
rlabel metal3 1740 1836 1740 1836 0 ccff_head_0
rlabel metal3 49734 4284 49734 4284 0 ccff_tail
rlabel metal1 1656 55726 1656 55726 0 ccff_tail_0
rlabel metal2 49358 25619 49358 25619 0 chanx_right_in[0]
rlabel metal2 48530 32249 48530 32249 0 chanx_right_in[10]
rlabel via2 49358 32861 49358 32861 0 chanx_right_in[11]
rlabel metal2 49358 33745 49358 33745 0 chanx_right_in[12]
rlabel metal2 49358 34391 49358 34391 0 chanx_right_in[13]
rlabel metal2 49358 34969 49358 34969 0 chanx_right_in[14]
rlabel metal2 49358 35615 49358 35615 0 chanx_right_in[15]
rlabel metal2 49358 36499 49358 36499 0 chanx_right_in[16]
rlabel metal2 48530 37111 48530 37111 0 chanx_right_in[17]
rlabel metal2 49358 37723 49358 37723 0 chanx_right_in[18]
rlabel via2 49358 38301 49358 38301 0 chanx_right_in[19]
rlabel metal2 48392 26044 48392 26044 0 chanx_right_in[1]
rlabel metal2 48530 39185 48530 39185 0 chanx_right_in[20]
rlabel metal2 48530 39797 48530 39797 0 chanx_right_in[21]
rlabel metal2 48530 40409 48530 40409 0 chanx_right_in[22]
rlabel via2 48530 41021 48530 41021 0 chanx_right_in[23]
rlabel metal2 48530 41905 48530 41905 0 chanx_right_in[24]
rlabel metal2 48530 42517 48530 42517 0 chanx_right_in[25]
rlabel metal2 48530 43129 48530 43129 0 chanx_right_in[26]
rlabel via2 48530 43741 48530 43741 0 chanx_right_in[27]
rlabel metal2 48530 44625 48530 44625 0 chanx_right_in[28]
rlabel metal1 48254 45458 48254 45458 0 chanx_right_in[29]
rlabel metal2 48530 26809 48530 26809 0 chanx_right_in[2]
rlabel via2 48530 27421 48530 27421 0 chanx_right_in[3]
rlabel metal2 49358 28305 49358 28305 0 chanx_right_in[4]
rlabel metal2 49358 28951 49358 28951 0 chanx_right_in[5]
rlabel metal2 48530 29529 48530 29529 0 chanx_right_in[6]
rlabel metal2 49358 30175 49358 30175 0 chanx_right_in[7]
rlabel metal2 48530 31025 48530 31025 0 chanx_right_in[8]
rlabel metal2 48530 31637 48530 31637 0 chanx_right_in[9]
rlabel metal3 49734 11764 49734 11764 0 chanx_right_out[10]
rlabel metal2 49174 12597 49174 12597 0 chanx_right_out[11]
rlabel metal3 49734 13124 49734 13124 0 chanx_right_out[12]
rlabel via2 49174 13821 49174 13821 0 chanx_right_out[13]
rlabel metal2 49174 14705 49174 14705 0 chanx_right_out[14]
rlabel metal3 49734 15164 49734 15164 0 chanx_right_out[15]
rlabel metal2 49174 15929 49174 15929 0 chanx_right_out[16]
rlabel via2 49174 16507 49174 16507 0 chanx_right_out[17]
rlabel metal3 49734 17204 49734 17204 0 chanx_right_out[18]
rlabel metal2 49174 18037 49174 18037 0 chanx_right_out[19]
rlabel metal3 49734 5644 49734 5644 0 chanx_right_out[1]
rlabel metal3 49734 18564 49734 18564 0 chanx_right_out[20]
rlabel metal2 49174 19295 49174 19295 0 chanx_right_out[21]
rlabel metal2 49174 20145 49174 20145 0 chanx_right_out[22]
rlabel metal3 49734 20604 49734 20604 0 chanx_right_out[23]
rlabel metal2 49174 21369 49174 21369 0 chanx_right_out[24]
rlabel metal3 49734 21964 49734 21964 0 chanx_right_out[25]
rlabel metal3 49734 22644 49734 22644 0 chanx_right_out[26]
rlabel metal2 49174 23477 49174 23477 0 chanx_right_out[27]
rlabel metal3 49734 24004 49734 24004 0 chanx_right_out[28]
rlabel via2 49174 24701 49174 24701 0 chanx_right_out[29]
rlabel metal3 49734 6324 49734 6324 0 chanx_right_out[2]
rlabel metal2 49174 7157 49174 7157 0 chanx_right_out[3]
rlabel metal3 49734 7684 49734 7684 0 chanx_right_out[4]
rlabel via2 49174 8381 49174 8381 0 chanx_right_out[5]
rlabel metal2 49174 9265 49174 9265 0 chanx_right_out[6]
rlabel metal3 49734 9724 49734 9724 0 chanx_right_out[7]
rlabel metal2 49174 10489 49174 10489 0 chanx_right_out[8]
rlabel metal3 49734 11084 49734 11084 0 chanx_right_out[9]
rlabel metal2 782 1860 782 1860 0 chany_bottom_in[0]
rlabel metal2 8142 823 8142 823 0 chany_bottom_in[10]
rlabel metal2 8878 1554 8878 1554 0 chany_bottom_in[11]
rlabel metal2 9614 1588 9614 1588 0 chany_bottom_in[12]
rlabel metal2 10350 1894 10350 1894 0 chany_bottom_in[13]
rlabel metal2 11086 1554 11086 1554 0 chany_bottom_in[14]
rlabel metal2 11822 1554 11822 1554 0 chany_bottom_in[15]
rlabel metal1 12650 3026 12650 3026 0 chany_bottom_in[16]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_in[17]
rlabel metal1 14076 3026 14076 3026 0 chany_bottom_in[18]
rlabel metal2 14766 1588 14766 1588 0 chany_bottom_in[19]
rlabel metal2 1518 1894 1518 1894 0 chany_bottom_in[1]
rlabel metal2 15502 1554 15502 1554 0 chany_bottom_in[20]
rlabel metal2 16238 1554 16238 1554 0 chany_bottom_in[21]
rlabel metal2 16974 1554 16974 1554 0 chany_bottom_in[22]
rlabel metal1 17756 3026 17756 3026 0 chany_bottom_in[23]
rlabel metal2 18446 1622 18446 1622 0 chany_bottom_in[24]
rlabel metal1 19228 2958 19228 2958 0 chany_bottom_in[25]
rlabel metal2 19918 1588 19918 1588 0 chany_bottom_in[26]
rlabel metal2 20654 1860 20654 1860 0 chany_bottom_in[27]
rlabel metal2 21390 1622 21390 1622 0 chany_bottom_in[28]
rlabel metal1 22080 2958 22080 2958 0 chany_bottom_in[29]
rlabel metal2 2254 1588 2254 1588 0 chany_bottom_in[2]
rlabel metal2 2990 1554 2990 1554 0 chany_bottom_in[3]
rlabel metal2 3726 1894 3726 1894 0 chany_bottom_in[4]
rlabel metal2 4462 1554 4462 1554 0 chany_bottom_in[5]
rlabel metal2 5198 1894 5198 1894 0 chany_bottom_in[6]
rlabel metal2 5934 1554 5934 1554 0 chany_bottom_in[7]
rlabel metal2 6670 1894 6670 1894 0 chany_bottom_in[8]
rlabel metal2 7406 1588 7406 1588 0 chany_bottom_in[9]
rlabel metal2 22862 1622 22862 1622 0 chany_bottom_out[0]
rlabel metal2 30222 1622 30222 1622 0 chany_bottom_out[10]
rlabel metal2 30958 2166 30958 2166 0 chany_bottom_out[11]
rlabel metal2 31694 1860 31694 1860 0 chany_bottom_out[12]
rlabel metal2 32430 1826 32430 1826 0 chany_bottom_out[13]
rlabel metal2 33166 1520 33166 1520 0 chany_bottom_out[14]
rlabel metal2 33902 2404 33902 2404 0 chany_bottom_out[15]
rlabel metal2 34638 2166 34638 2166 0 chany_bottom_out[16]
rlabel metal2 35374 1622 35374 1622 0 chany_bottom_out[17]
rlabel metal2 36110 2166 36110 2166 0 chany_bottom_out[18]
rlabel metal2 36846 1860 36846 1860 0 chany_bottom_out[19]
rlabel metal1 23690 2958 23690 2958 0 chany_bottom_out[1]
rlabel metal2 37582 1826 37582 1826 0 chany_bottom_out[20]
rlabel metal2 38318 1622 38318 1622 0 chany_bottom_out[21]
rlabel metal2 39054 2404 39054 2404 0 chany_bottom_out[22]
rlabel metal2 39790 2166 39790 2166 0 chany_bottom_out[23]
rlabel metal2 40526 1622 40526 1622 0 chany_bottom_out[24]
rlabel metal2 41262 2166 41262 2166 0 chany_bottom_out[25]
rlabel metal2 41998 1860 41998 1860 0 chany_bottom_out[26]
rlabel metal2 42734 1826 42734 1826 0 chany_bottom_out[27]
rlabel metal2 43470 2404 43470 2404 0 chany_bottom_out[28]
rlabel metal2 44206 2166 44206 2166 0 chany_bottom_out[29]
rlabel metal1 24702 3570 24702 3570 0 chany_bottom_out[2]
rlabel metal1 25346 2958 25346 2958 0 chany_bottom_out[3]
rlabel metal2 25806 1622 25806 1622 0 chany_bottom_out[4]
rlabel metal2 26542 1622 26542 1622 0 chany_bottom_out[5]
rlabel metal1 27554 2958 27554 2958 0 chany_bottom_out[6]
rlabel metal2 28014 823 28014 823 0 chany_bottom_out[7]
rlabel metal1 29210 2958 29210 2958 0 chany_bottom_out[8]
rlabel metal1 29854 3570 29854 3570 0 chany_bottom_out[9]
rlabel metal2 23230 55711 23230 55711 0 chany_top_in_0[0]
rlabel metal1 30636 54162 30636 54162 0 chany_top_in_0[10]
rlabel metal1 31372 54162 31372 54162 0 chany_top_in_0[11]
rlabel metal1 32200 53550 32200 53550 0 chany_top_in_0[12]
rlabel metal1 32890 54230 32890 54230 0 chany_top_in_0[13]
rlabel metal1 33626 54230 33626 54230 0 chany_top_in_0[14]
rlabel metal1 34592 54162 34592 54162 0 chany_top_in_0[15]
rlabel metal1 35144 53550 35144 53550 0 chany_top_in_0[16]
rlabel metal1 35788 54162 35788 54162 0 chany_top_in_0[17]
rlabel metal1 36524 54162 36524 54162 0 chany_top_in_0[18]
rlabel metal1 37398 54230 37398 54230 0 chany_top_in_0[19]
rlabel metal1 24334 53550 24334 53550 0 chany_top_in_0[1]
rlabel metal2 37950 55711 37950 55711 0 chany_top_in_0[20]
rlabel metal1 38732 54162 38732 54162 0 chany_top_in_0[21]
rlabel metal1 39744 54162 39744 54162 0 chany_top_in_0[22]
rlabel metal1 40480 54162 40480 54162 0 chany_top_in_0[23]
rlabel metal1 41308 54162 41308 54162 0 chany_top_in_0[24]
rlabel metal1 41768 53550 41768 53550 0 chany_top_in_0[25]
rlabel metal1 42550 54230 42550 54230 0 chany_top_in_0[26]
rlabel metal1 43424 54162 43424 54162 0 chany_top_in_0[27]
rlabel metal2 44022 56236 44022 56236 0 chany_top_in_0[28]
rlabel metal1 44988 54162 44988 54162 0 chany_top_in_0[29]
rlabel metal1 24794 54230 24794 54230 0 chany_top_in_0[2]
rlabel metal1 25484 54162 25484 54162 0 chany_top_in_0[3]
rlabel metal2 26174 55209 26174 55209 0 chany_top_in_0[4]
rlabel metal1 27048 54162 27048 54162 0 chany_top_in_0[5]
rlabel metal1 27784 54162 27784 54162 0 chany_top_in_0[6]
rlabel metal1 28566 54230 28566 54230 0 chany_top_in_0[7]
rlabel metal1 29532 53550 29532 53550 0 chany_top_in_0[8]
rlabel metal1 29900 54162 29900 54162 0 chany_top_in_0[9]
rlabel metal1 1610 52530 1610 52530 0 chany_top_out_0[0]
rlabel metal1 8464 54230 8464 54230 0 chany_top_out_0[10]
rlabel metal1 9522 52530 9522 52530 0 chany_top_out_0[11]
rlabel metal1 10120 53006 10120 53006 0 chany_top_out_0[12]
rlabel metal1 10810 53618 10810 53618 0 chany_top_out_0[13]
rlabel metal1 11224 54230 11224 54230 0 chany_top_out_0[14]
rlabel metal1 12466 53618 12466 53618 0 chany_top_out_0[15]
rlabel metal2 12926 55711 12926 55711 0 chany_top_out_0[16]
rlabel metal1 13616 54230 13616 54230 0 chany_top_out_0[17]
rlabel metal1 14674 52530 14674 52530 0 chany_top_out_0[18]
rlabel metal1 15272 53006 15272 53006 0 chany_top_out_0[19]
rlabel metal1 2162 53618 2162 53618 0 chany_top_out_0[1]
rlabel metal1 15870 53652 15870 53652 0 chany_top_out_0[20]
rlabel metal2 16606 55226 16606 55226 0 chany_top_out_0[21]
rlabel metal1 17618 53006 17618 53006 0 chany_top_out_0[22]
rlabel metal2 18262 56236 18262 56236 0 chany_top_out_0[23]
rlabel metal1 18768 54230 18768 54230 0 chany_top_out_0[24]
rlabel metal1 19826 53006 19826 53006 0 chany_top_out_0[25]
rlabel metal1 20378 53618 20378 53618 0 chany_top_out_0[26]
rlabel metal2 21022 55226 21022 55226 0 chany_top_out_0[27]
rlabel metal1 22034 53618 22034 53618 0 chany_top_out_0[28]
rlabel metal1 22770 54094 22770 54094 0 chany_top_out_0[29]
rlabel metal1 2898 53006 2898 53006 0 chany_top_out_0[2]
rlabel metal1 3312 54230 3312 54230 0 chany_top_out_0[3]
rlabel metal1 4370 52530 4370 52530 0 chany_top_out_0[4]
rlabel metal2 4830 55711 4830 55711 0 chany_top_out_0[5]
rlabel metal1 5658 53618 5658 53618 0 chany_top_out_0[6]
rlabel metal1 6072 54230 6072 54230 0 chany_top_out_0[7]
rlabel metal1 7314 53618 7314 53618 0 chany_top_out_0[8]
rlabel metal1 8050 53006 8050 53006 0 chany_top_out_0[9]
rlabel metal1 22034 19448 22034 19448 0 clknet_0_prog_clk
rlabel metal1 19044 16626 19044 16626 0 clknet_4_0_0_prog_clk
rlabel metal2 38548 21522 38548 21522 0 clknet_4_10_0_prog_clk
rlabel metal1 37812 32402 37812 32402 0 clknet_4_11_0_prog_clk
rlabel metal2 32614 38930 32614 38930 0 clknet_4_12_0_prog_clk
rlabel metal1 24150 42228 24150 42228 0 clknet_4_13_0_prog_clk
rlabel metal1 42366 37298 42366 37298 0 clknet_4_14_0_prog_clk
rlabel metal1 37490 41650 37490 41650 0 clknet_4_15_0_prog_clk
rlabel metal2 19642 20740 19642 20740 0 clknet_4_1_0_prog_clk
rlabel metal1 32039 18190 32039 18190 0 clknet_4_2_0_prog_clk
rlabel metal2 32522 21318 32522 21318 0 clknet_4_3_0_prog_clk
rlabel metal1 12374 23664 12374 23664 0 clknet_4_4_0_prog_clk
rlabel metal2 21114 33150 21114 33150 0 clknet_4_5_0_prog_clk
rlabel metal2 28474 25364 28474 25364 0 clknet_4_6_0_prog_clk
rlabel metal1 22172 41650 22172 41650 0 clknet_4_7_0_prog_clk
rlabel metal2 34914 14790 34914 14790 0 clknet_4_8_0_prog_clk
rlabel metal1 32338 32334 32338 32334 0 clknet_4_9_0_prog_clk
rlabel metal3 1740 13396 1740 13396 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 15708 1004 15708 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18020 1004 18020 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 20332 1004 20332 0 gfpga_pad_io_soc_dir[3]
rlabel metal3 820 31892 820 31892 0 gfpga_pad_io_soc_in[0]
rlabel metal3 1234 34204 1234 34204 0 gfpga_pad_io_soc_in[1]
rlabel metal3 820 36516 820 36516 0 gfpga_pad_io_soc_in[2]
rlabel metal3 820 38828 820 38828 0 gfpga_pad_io_soc_in[3]
rlabel metal3 1004 22644 1004 22644 0 gfpga_pad_io_soc_out[0]
rlabel metal3 1004 24956 1004 24956 0 gfpga_pad_io_soc_out[1]
rlabel metal3 1004 27268 1004 27268 0 gfpga_pad_io_soc_out[2]
rlabel metal3 1004 29580 1004 29580 0 gfpga_pad_io_soc_out[3]
rlabel metal3 1188 41140 1188 41140 0 isol_n
rlabel metal2 4002 51000 4002 51000 0 net1
rlabel metal2 44574 34748 44574 34748 0 net10
rlabel metal1 48990 47430 48990 47430 0 net100
rlabel metal1 44712 47974 44712 47974 0 net101
rlabel metal2 41630 36992 41630 36992 0 net102
rlabel metal1 49082 49062 49082 49062 0 net103
rlabel metal2 43930 39236 43930 39236 0 net104
rlabel metal1 49358 50694 49358 50694 0 net105
rlabel metal2 48990 35025 48990 35025 0 net106
rlabel metal2 49266 42840 49266 42840 0 net107
rlabel metal1 48760 6290 48760 6290 0 net108
rlabel metal2 1794 45696 1794 45696 0 net109
rlabel metal1 41814 36312 41814 36312 0 net11
rlabel metal1 21482 39304 21482 39304 0 net110
rlabel metal2 1748 42228 1748 42228 0 net111
rlabel metal1 1932 52938 1932 52938 0 net112
rlabel metal1 18998 18938 18998 18938 0 net113
rlabel metal2 23690 41718 23690 41718 0 net114
rlabel metal2 44758 12444 44758 12444 0 net115
rlabel metal2 46782 12988 46782 12988 0 net116
rlabel metal1 43838 17510 43838 17510 0 net117
rlabel metal1 44666 17578 44666 17578 0 net118
rlabel metal1 45356 17034 45356 17034 0 net119
rlabel metal1 42504 37910 42504 37910 0 net12
rlabel metal1 45034 17646 45034 17646 0 net120
rlabel metal1 46138 18666 46138 18666 0 net121
rlabel metal1 45310 19754 45310 19754 0 net122
rlabel metal2 45218 19244 45218 19244 0 net123
rlabel metal2 46782 20366 46782 20366 0 net124
rlabel metal1 47104 5678 47104 5678 0 net125
rlabel metal2 44666 21964 44666 21964 0 net126
rlabel metal2 45494 22270 45494 22270 0 net127
rlabel metal1 47932 20434 47932 20434 0 net128
rlabel metal1 47518 20910 47518 20910 0 net129
rlabel metal1 37628 37978 37628 37978 0 net13
rlabel metal1 47150 21522 47150 21522 0 net130
rlabel metal1 47794 21998 47794 21998 0 net131
rlabel metal1 47840 23086 47840 23086 0 net132
rlabel metal1 47380 23698 47380 23698 0 net133
rlabel metal1 47886 24174 47886 24174 0 net134
rlabel metal2 47242 25500 47242 25500 0 net135
rlabel metal1 46966 6834 46966 6834 0 net136
rlabel metal1 47932 7378 47932 7378 0 net137
rlabel metal1 47150 7854 47150 7854 0 net138
rlabel metal1 47242 8466 47242 8466 0 net139
rlabel via2 42182 27115 42182 27115 0 net14
rlabel metal1 47334 9554 47334 9554 0 net140
rlabel metal2 46782 10846 46782 10846 0 net141
rlabel metal2 47886 5949 47886 5949 0 net142
rlabel metal2 44298 11594 44298 11594 0 net143
rlabel metal1 23736 15334 23736 15334 0 net144
rlabel metal1 31694 2414 31694 2414 0 net145
rlabel metal1 30866 3502 30866 3502 0 net146
rlabel metal1 32936 3026 32936 3026 0 net147
rlabel metal1 34224 19754 34224 19754 0 net148
rlabel metal1 34362 2414 34362 2414 0 net149
rlabel via2 48806 39491 48806 39491 0 net15
rlabel metal1 33304 9418 33304 9418 0 net150
rlabel metal1 34592 3502 34592 3502 0 net151
rlabel metal1 36386 2414 36386 2414 0 net152
rlabel metal1 36616 18666 36616 18666 0 net153
rlabel metal1 37904 8330 37904 8330 0 net154
rlabel metal1 25116 15538 25116 15538 0 net155
rlabel metal1 38318 3094 38318 3094 0 net156
rlabel metal1 38916 13974 38916 13974 0 net157
rlabel metal1 38778 4114 38778 4114 0 net158
rlabel metal1 38732 3502 38732 3502 0 net159
rlabel metal1 48806 39882 48806 39882 0 net16
rlabel metal1 42044 2414 42044 2414 0 net160
rlabel metal1 40572 12138 40572 12138 0 net161
rlabel metal1 39698 8398 39698 8398 0 net162
rlabel metal1 41492 6698 41492 6698 0 net163
rlabel metal1 38962 6766 38962 6766 0 net164
rlabel metal1 41492 7242 41492 7242 0 net165
rlabel metal1 25208 13158 25208 13158 0 net166
rlabel metal2 25162 6766 25162 6766 0 net167
rlabel metal1 26312 12614 26312 12614 0 net168
rlabel metal1 27692 12682 27692 12682 0 net169
rlabel metal1 44482 34986 44482 34986 0 net17
rlabel metal1 28244 15334 28244 15334 0 net170
rlabel metal2 29946 6154 29946 6154 0 net171
rlabel metal2 29210 7582 29210 7582 0 net172
rlabel metal1 29486 13838 29486 13838 0 net173
rlabel metal1 2760 52462 2760 52462 0 net174
rlabel metal1 12650 43962 12650 43962 0 net175
rlabel metal1 12006 52462 12006 52462 0 net176
rlabel metal1 12098 44506 12098 44506 0 net177
rlabel metal1 12788 45526 12788 45526 0 net178
rlabel metal1 15456 43962 15456 43962 0 net179
rlabel metal1 48714 41038 48714 41038 0 net18
rlabel metal1 13570 53550 13570 53550 0 net180
rlabel metal2 16974 48552 16974 48552 0 net181
rlabel metal1 16008 42738 16008 42738 0 net182
rlabel metal2 19182 47940 19182 47940 0 net183
rlabel metal1 15134 53074 15134 53074 0 net184
rlabel metal1 2162 53516 2162 53516 0 net185
rlabel metal2 20470 48688 20470 48688 0 net186
rlabel metal2 20378 44479 20378 44479 0 net187
rlabel metal1 17618 53108 17618 53108 0 net188
rlabel metal1 18078 53550 18078 53550 0 net189
rlabel metal1 48806 42092 48806 42092 0 net19
rlabel metal2 17710 52326 17710 52326 0 net190
rlabel metal1 21298 43894 21298 43894 0 net191
rlabel metal1 20194 53516 20194 53516 0 net192
rlabel metal1 20332 54162 20332 54162 0 net193
rlabel metal1 23782 51578 23782 51578 0 net194
rlabel metal1 23184 52122 23184 52122 0 net195
rlabel metal1 2898 53108 2898 53108 0 net196
rlabel metal1 2254 54128 2254 54128 0 net197
rlabel metal1 9292 42738 9292 42738 0 net198
rlabel metal1 5865 53074 5865 53074 0 net199
rlabel metal1 3588 3706 3588 3706 0 net2
rlabel metal1 48806 42602 48806 42602 0 net20
rlabel metal1 6187 53550 6187 53550 0 net200
rlabel metal1 4830 54230 4830 54230 0 net201
rlabel metal1 10626 43214 10626 43214 0 net202
rlabel metal1 10718 43894 10718 43894 0 net203
rlabel metal1 3726 13906 3726 13906 0 net204
rlabel metal1 3772 18598 3772 18598 0 net205
rlabel metal1 2346 18258 2346 18258 0 net206
rlabel metal1 2300 20434 2300 20434 0 net207
rlabel metal1 2668 23086 2668 23086 0 net208
rlabel metal1 2990 25262 2990 25262 0 net209
rlabel metal2 41676 37196 41676 37196 0 net21
rlabel metal1 3404 27438 3404 27438 0 net210
rlabel metal2 4830 28900 4830 28900 0 net211
rlabel metal2 47794 3162 47794 3162 0 net212
rlabel metal2 48622 45764 48622 45764 0 net213
rlabel metal2 46230 53380 46230 53380 0 net214
rlabel metal1 47380 6630 47380 6630 0 net215
rlabel metal1 47932 31450 47932 31450 0 net216
rlabel metal1 48254 3502 48254 3502 0 net217
rlabel metal1 48254 30906 48254 30906 0 net218
rlabel metal1 30590 20502 30590 20502 0 net219
rlabel metal1 43171 43758 43171 43758 0 net22
rlabel metal1 28980 27438 28980 27438 0 net220
rlabel metal1 42918 31450 42918 31450 0 net221
rlabel metal1 39422 23086 39422 23086 0 net222
rlabel metal1 32430 36176 32430 36176 0 net223
rlabel metal1 31970 22610 31970 22610 0 net224
rlabel metal2 39054 28356 39054 28356 0 net225
rlabel metal1 31648 33966 31648 33966 0 net226
rlabel metal1 32246 34714 32246 34714 0 net227
rlabel metal1 33304 35666 33304 35666 0 net228
rlabel metal1 29670 37230 29670 37230 0 net229
rlabel metal1 41975 44846 41975 44846 0 net23
rlabel metal1 27600 36346 27600 36346 0 net230
rlabel metal2 41722 34884 41722 34884 0 net231
rlabel metal1 28244 32402 28244 32402 0 net232
rlabel metal1 26220 29614 26220 29614 0 net233
rlabel metal2 27002 26554 27002 26554 0 net234
rlabel metal2 25898 25262 25898 25262 0 net235
rlabel metal2 24978 23290 24978 23290 0 net236
rlabel metal1 25438 23732 25438 23732 0 net237
rlabel metal1 24656 25874 24656 25874 0 net238
rlabel metal2 23138 27268 23138 27268 0 net239
rlabel metal1 43102 37740 43102 37740 0 net24
rlabel metal1 13938 11118 13938 11118 0 net240
rlabel metal2 30222 14586 30222 14586 0 net241
rlabel metal1 34914 32878 34914 32878 0 net242
rlabel metal2 32246 14790 32246 14790 0 net243
rlabel metal2 33442 15674 33442 15674 0 net244
rlabel metal1 35696 17170 35696 17170 0 net245
rlabel metal1 37996 16558 37996 16558 0 net246
rlabel metal1 33856 16082 33856 16082 0 net247
rlabel metal1 38088 14382 38088 14382 0 net248
rlabel metal1 36432 12410 36432 12410 0 net249
rlabel metal1 41630 27404 41630 27404 0 net25
rlabel metal1 37766 15130 37766 15130 0 net250
rlabel metal2 41446 36686 41446 36686 0 net251
rlabel metal1 39054 36754 39054 36754 0 net252
rlabel metal2 23690 36346 23690 36346 0 net253
rlabel metal2 21850 30906 21850 30906 0 net254
rlabel metal1 24334 31790 24334 31790 0 net255
rlabel metal2 31326 37434 31326 37434 0 net256
rlabel metal2 23598 30362 23598 30362 0 net257
rlabel metal1 18124 32402 18124 32402 0 net258
rlabel metal2 22494 37434 22494 37434 0 net259
rlabel metal1 41630 26826 41630 26826 0 net26
rlabel metal1 26450 35122 26450 35122 0 net260
rlabel metal1 24242 37230 24242 37230 0 net261
rlabel metal2 29118 33796 29118 33796 0 net262
rlabel metal2 22862 31076 22862 31076 0 net263
rlabel via2 49358 4981 49358 4981 0 net264
rlabel metal1 24518 25262 24518 25262 0 net265
rlabel metal1 25484 22610 25484 22610 0 net266
rlabel metal2 23230 17476 23230 17476 0 net267
rlabel metal1 22816 24786 22816 24786 0 net268
rlabel metal1 29486 21658 29486 21658 0 net269
rlabel metal2 39514 28356 39514 28356 0 net27
rlabel metal1 28566 24106 28566 24106 0 net270
rlabel metal2 36938 25432 36938 25432 0 net271
rlabel metal1 40342 24786 40342 24786 0 net272
rlabel metal1 36432 28526 36432 28526 0 net273
rlabel metal1 45540 29070 45540 29070 0 net28
rlabel metal1 37214 33830 37214 33830 0 net29
rlabel metal2 49174 25568 49174 25568 0 net3
rlabel metal1 42780 31382 42780 31382 0 net30
rlabel metal2 42274 37536 42274 37536 0 net31
rlabel metal1 45540 31926 45540 31926 0 net32
rlabel metal1 4646 2856 4646 2856 0 net33
rlabel metal2 21942 39814 21942 39814 0 net34
rlabel metal2 13478 38080 13478 38080 0 net35
rlabel metal2 10074 3740 10074 3740 0 net36
rlabel metal1 12558 2890 12558 2890 0 net37
rlabel metal2 21574 41446 21574 41446 0 net38
rlabel metal2 21206 35632 21206 35632 0 net39
rlabel metal2 48806 32708 48806 32708 0 net4
rlabel metal2 12834 3264 12834 3264 0 net40
rlabel metal3 19320 35088 19320 35088 0 net41
rlabel metal1 17342 42602 17342 42602 0 net42
rlabel metal1 16652 2618 16652 2618 0 net43
rlabel metal1 1794 2924 1794 2924 0 net44
rlabel metal2 15318 2125 15318 2125 0 net45
rlabel metal1 20378 43792 20378 43792 0 net46
rlabel metal2 20286 37740 20286 37740 0 net47
rlabel metal2 17986 3111 17986 3111 0 net48
rlabel metal2 18354 2142 18354 2142 0 net49
rlabel metal2 49174 32640 49174 32640 0 net5
rlabel metal1 20838 3094 20838 3094 0 net50
rlabel metal1 23966 2550 23966 2550 0 net51
rlabel metal1 20930 3060 20930 3060 0 net52
rlabel metal2 20930 2108 20930 2108 0 net53
rlabel metal1 27554 16218 27554 16218 0 net54
rlabel metal2 2438 2040 2438 2040 0 net55
rlabel metal2 3358 2006 3358 2006 0 net56
rlabel metal1 20148 17510 20148 17510 0 net57
rlabel via1 21022 21930 21022 21930 0 net58
rlabel via2 5474 2907 5474 2907 0 net59
rlabel metal1 39284 30702 39284 30702 0 net6
rlabel via2 6026 2363 6026 2363 0 net60
rlabel metal1 21206 18598 21206 18598 0 net61
rlabel metal2 12098 38012 12098 38012 0 net62
rlabel metal1 25392 53686 25392 53686 0 net63
rlabel metal1 30682 53958 30682 53958 0 net64
rlabel metal1 30268 54298 30268 54298 0 net65
rlabel metal1 33028 45526 33028 45526 0 net66
rlabel metal1 33120 45458 33120 45458 0 net67
rlabel metal1 33948 54026 33948 54026 0 net68
rlabel via2 35282 44693 35282 44693 0 net69
rlabel metal2 49174 34986 49174 34986 0 net7
rlabel metal1 35236 53414 35236 53414 0 net70
rlabel metal2 36570 44319 36570 44319 0 net71
rlabel metal1 37444 43690 37444 43690 0 net72
rlabel metal3 37467 44268 37467 44268 0 net73
rlabel metal1 25346 53482 25346 53482 0 net74
rlabel metal1 37260 44506 37260 44506 0 net75
rlabel metal1 40020 43282 40020 43282 0 net76
rlabel metal2 40434 42109 40434 42109 0 net77
rlabel metal1 41492 42194 41492 42194 0 net78
rlabel metal1 39652 54298 39652 54298 0 net79
rlabel metal1 49128 34918 49128 34918 0 net8
rlabel metal1 39974 44506 39974 44506 0 net80
rlabel metal1 38686 12206 38686 12206 0 net81
rlabel metal1 40986 54026 40986 54026 0 net82
rlabel metal1 41998 42670 41998 42670 0 net83
rlabel metal1 43470 42330 43470 42330 0 net84
rlabel metal1 25162 54026 25162 54026 0 net85
rlabel metal1 25898 53958 25898 53958 0 net86
rlabel metal1 28198 43690 28198 43690 0 net87
rlabel metal1 27416 53958 27416 53958 0 net88
rlabel metal1 28336 53958 28336 53958 0 net89
rlabel metal1 42182 32878 42182 32878 0 net9
rlabel metal1 29302 54026 29302 54026 0 net90
rlabel metal1 31234 45458 31234 45458 0 net91
rlabel metal3 29785 12852 29785 12852 0 net92
rlabel metal1 7544 25874 7544 25874 0 net93
rlabel metal2 7866 30838 7866 30838 0 net94
rlabel metal1 4600 36550 4600 36550 0 net95
rlabel metal1 4508 38726 4508 38726 0 net96
rlabel metal2 12650 20366 12650 20366 0 net97
rlabel metal1 21489 35734 21489 35734 0 net98
rlabel metal2 47426 4896 47426 4896 0 net99
rlabel metal2 44942 10360 44942 10360 0 prog_clk
rlabel metal2 45678 1554 45678 1554 0 prog_reset_bottom_in
rlabel metal2 46414 1792 46414 1792 0 prog_reset_bottom_out
rlabel metal3 49734 45764 49734 45764 0 prog_reset_right_out
rlabel metal1 47058 53618 47058 53618 0 prog_reset_top_out
rlabel metal2 47150 1860 47150 1860 0 reset_bottom_in
rlabel metal2 47886 1860 47886 1860 0 reset_bottom_out
rlabel metal2 48300 54604 48300 54604 0 reset_top_out
rlabel metal2 49082 47379 49082 47379 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 49082 47957 49082 47957 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 49082 48603 49082 48603 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel via2 49082 49181 49082 49181 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 49082 50065 49082 50065 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 48990 50711 48990 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 49082 51289 49082 51289 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 49082 51935 49082 51935 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 2062 4148 2062 4148 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 2062 6460 2062 6460 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 2016 8772 2016 8772 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 2062 11084 2062 11084 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 36662 17816 36662 17816 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel metal2 31786 21318 31786 21318 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 35466 19312 35466 19312 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 32246 23290 32246 23290 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal2 34270 23630 34270 23630 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal1 33948 26418 33948 26418 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal1 33856 25806 33856 25806 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal2 32522 26044 32522 26044 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal2 39514 25874 39514 25874 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal1 41170 32946 41170 32946 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 37720 25194 37720 25194 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal2 40802 26826 40802 26826 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal2 42274 32300 42274 32300 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal2 40710 27846 40710 27846 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal1 35650 29274 35650 29274 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 41722 27574 41722 27574 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 36478 28594 36478 28594 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal2 34270 20842 34270 20842 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 33902 26894 33902 26894 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 33442 21454 33442 21454 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal1 34582 33082 34582 33082 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal1 35742 31926 35742 31926 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 35282 32402 35282 32402 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal1 37069 34374 37069 34374 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal1 40894 33422 40894 33422 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal2 42090 32300 42090 32300 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal1 38134 20978 38134 20978 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal1 41538 30124 41538 30124 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 39974 23834 39974 23834 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal1 21942 41480 21942 41480 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal1 35696 28594 35696 28594 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal2 35190 23324 35190 23324 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal1 33948 35258 33948 35258 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal2 42734 30838 42734 30838 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal1 37996 31858 37996 31858 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal2 40526 29002 40526 29002 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal1 38962 42126 38962 42126 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal1 37030 41514 37030 41514 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 38134 43826 38134 43826 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal1 35236 38250 35236 38250 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal1 35512 41446 35512 41446 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal1 36432 42738 36432 42738 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal1 37306 42534 37306 42534 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal1 35328 40902 35328 40902 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal2 35558 43350 35558 43350 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal1 35282 41990 35282 41990 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal1 33718 41446 33718 41446 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel metal1 33297 43078 33297 43078 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 31464 41514 31464 41514 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal1 31878 41990 31878 41990 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal1 32154 43826 32154 43826 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal1 29854 42262 29854 42262 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal1 43003 37434 43003 37434 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal1 43056 35734 43056 35734 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 42642 36210 42642 36210 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal1 30774 34374 30774 34374 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel metal1 28750 43826 28750 43826 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal1 32223 37298 32223 37298 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel metal2 28842 29920 28842 29920 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 28290 35258 28290 35258 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal1 27784 34034 27784 34034 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal1 29394 26894 29394 26894 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal1 28060 28118 28060 28118 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal1 30084 25670 30084 25670 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal1 30222 26758 30222 26758 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 28244 22542 28244 22542 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal1 31234 24718 31234 24718 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 28290 24582 28290 24582 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 27501 24582 27501 24582 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal1 27002 27302 27002 27302 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal1 28888 25466 28888 25466 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal2 24242 27166 24242 27166 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal1 28382 28186 28382 28186 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal2 21206 15674 21206 15674 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 20815 21454 20815 21454 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal1 19136 19890 19136 19890 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel metal1 28520 14926 28520 14926 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal2 26174 15164 26174 15164 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal1 39928 35802 39928 35802 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 41722 37128 41722 37128 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel via1 38410 35581 38410 35581 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal2 32890 15402 32890 15402 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal1 29302 16014 29302 16014 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal2 33534 16320 33534 16320 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal2 30314 16541 30314 16541 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal1 35098 18190 35098 18190 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal1 32568 18326 32568 18326 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 37352 17850 37352 17850 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal1 35880 17578 35880 17578 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal1 38364 18190 38364 18190 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal1 37628 19278 37628 19278 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal2 37766 13906 37766 13906 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal1 36616 15538 36616 15538 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal2 35466 13328 35466 13328 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel metal2 33994 13668 33994 13668 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal1 35374 16626 35374 16626 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 43056 38454 43056 38454 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal2 41078 35258 41078 35258 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal2 41814 37230 41814 37230 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal1 39008 44302 39008 44302 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal1 39698 40562 39698 40562 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal2 27370 43044 27370 43044 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal2 21850 42245 21850 42245 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal2 25898 40426 25898 40426 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal1 24932 37638 24932 37638 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal1 22356 36346 22356 36346 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel metal1 32614 35632 32614 35632 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal1 20838 36040 20838 36040 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal2 25622 33286 25622 33286 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal2 36938 30566 36938 30566 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 28474 32266 28474 32266 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal2 30038 39644 30038 39644 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal1 35144 39474 35144 39474 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 32338 39542 32338 39542 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal1 24012 34034 24012 34034 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal1 33350 31178 33350 31178 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal1 23276 31858 23276 31858 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal1 21344 35802 21344 35802 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel via1 29026 31875 29026 31875 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal2 23322 35360 23322 35360 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal1 25024 40154 25024 40154 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 26634 39474 26634 39474 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal1 23552 39950 23552 39950 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal1 27646 37774 27646 37774 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 35282 33320 35282 33320 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal2 32338 36142 32338 36142 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 32430 39916 32430 39916 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal1 27416 41038 27416 41038 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal2 43194 37876 43194 37876 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal1 36478 36550 36478 36550 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal2 38042 36380 38042 36380 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal1 27646 38352 27646 38352 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 28474 16150 28474 16150 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal1 32154 25330 32154 25330 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33534 25262 33534 25262 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 25622 21726 25622 21726 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31096 20774 31096 20774 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 30682 21114 30682 21114 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 30176 17578 30176 17578 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 33810 7446 33810 7446 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal1 33488 28594 33488 28594 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37674 33082 37674 33082 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31924 26010 31924 26010 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27646 23902 27646 23902 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32936 24786 32936 24786 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 31050 25296 31050 25296 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 32476 17170 32476 17170 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 35512 9622 35512 9622 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal1 36478 28458 36478 28458 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40342 32742 40342 32742 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36938 25330 36938 25330 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37628 24786 37628 24786 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37214 24922 37214 24922 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 35236 19822 35236 19822 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 38226 8534 38226 8534 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal1 39744 28458 39744 28458 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 41354 32742 41354 32742 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 39008 25330 39008 25330 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40388 24242 40388 24242 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 40250 24174 40250 24174 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39514 16082 39514 16082 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 32246 9622 32246 9622 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal1 35052 31858 35052 31858 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38272 34510 38272 34510 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37030 28186 37030 28186 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 35466 30345 35466 30345 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35696 27438 35696 27438 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33580 20978 33580 20978 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 35006 6698 35006 6698 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal2 33994 26044 33994 26044 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34408 25194 34408 25194 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32844 20570 32844 20570 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32269 20502 32269 20502 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 32614 17850 32614 17850 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 27922 21318 27922 21318 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal2 35190 34476 35190 34476 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36432 32538 36432 32538 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34638 32198 34638 32198 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 27574 28612 27574 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 28428 21522 28428 21522 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 31832 16116 31832 16116 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal2 42182 35836 42182 35836 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 41446 31654 41446 31654 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 39974 29614 39974 29614 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36110 19822 36110 19822 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37122 6766 37122 6766 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal1 37628 26418 37628 26418 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39560 26350 39560 26350 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38088 23018 38088 23018 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38364 20774 38364 20774 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38272 20910 38272 20910 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 36386 16082 36386 16082 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 23828 17170 23828 17170 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal2 32246 37468 32246 37468 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32062 36618 32062 36618 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25024 27030 25024 27030 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34454 8534 34454 8534 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal1 35374 25194 35374 25194 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36018 25126 36018 25126 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34454 23766 34454 23766 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32706 23188 32706 23188 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 34178 23902 34178 23902 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 34316 22746 34316 22746 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 33028 22406 33028 22406 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 44022 26826 44022 26826 0 sb_0__1_.mux_right_track_0.out
rlabel metal1 39238 31926 39238 31926 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40434 30906 40434 30906 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 40664 29274 40664 29274 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 39928 27914 39928 27914 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 44206 28220 44206 28220 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 46138 28288 46138 28288 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 37628 39066 37628 39066 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37582 38930 37582 38930 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36984 35054 36984 35054 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 36386 34510 36386 34510 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36110 34918 36110 34918 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 41998 28220 41998 28220 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 36524 38930 36524 38930 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36616 36210 36616 36210 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32338 34476 32338 34476 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36386 36006 36386 36006 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 46046 28220 46046 28220 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 35466 44982 35466 44982 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 35558 36771 35558 36771 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32752 35462 32752 35462 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35834 36278 35834 36278 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 45310 28764 45310 28764 0 sb_0__1_.mux_right_track_16.out
rlabel metal1 33810 40562 33810 40562 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33902 39066 33902 39066 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 33350 38046 33350 38046 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 39422 31790 39422 31790 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 42941 25194 42941 25194 0 sb_0__1_.mux_right_track_18.out
rlabel metal1 32522 45254 32522 45254 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 34178 39406 34178 39406 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31970 36312 31970 36312 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34270 38454 34270 38454 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 46966 29614 46966 29614 0 sb_0__1_.mux_right_track_2.out
rlabel metal2 42366 39100 42366 39100 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 42274 35768 42274 35768 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 40894 34034 40894 34034 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 42366 36278 42366 36278 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 41354 34680 41354 34680 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 44298 32912 44298 32912 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43562 22678 43562 22678 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 30544 43962 30544 43962 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32154 34986 32154 34986 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29302 32538 29302 32538 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34408 27098 34408 27098 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 43838 22746 43838 22746 0 sb_0__1_.mux_right_track_22.out
rlabel metal1 29946 33422 29946 33422 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30084 29478 30084 29478 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30130 29648 30130 29648 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 36662 27166 36662 27166 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 44160 19822 44160 19822 0 sb_0__1_.mux_right_track_24.out
rlabel metal2 31188 26418 31188 26418 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 31142 26418 31142 26418 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35558 24752 35558 24752 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 44206 20298 44206 20298 0 sb_0__1_.mux_right_track_26.out
rlabel metal2 31970 27370 31970 27370 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26404 24650 26404 24650 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36846 22032 36846 22032 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 44482 18904 44482 18904 0 sb_0__1_.mux_right_track_28.out
rlabel metal1 30268 22746 30268 22746 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27508 22746 27508 22746 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 36938 21454 36938 21454 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43746 19142 43746 19142 0 sb_0__1_.mux_right_track_30.out
rlabel metal2 30222 25772 30222 25772 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28198 24174 28198 24174 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35788 20910 35788 20910 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43378 19482 43378 19482 0 sb_0__1_.mux_right_track_32.out
rlabel metal1 28934 25262 28934 25262 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28750 25296 28750 25296 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33166 21624 33166 21624 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 42826 19380 42826 19380 0 sb_0__1_.mux_right_track_34.out
rlabel metal1 28612 26350 28612 26350 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 28198 26588 28198 26588 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28198 22066 28198 22066 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35466 13872 35466 13872 0 sb_0__1_.mux_right_track_36.out
rlabel metal2 18630 20094 18630 20094 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20056 17748 20056 17748 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17066 13158 17066 13158 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20562 14688 20562 14688 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 38594 13464 38594 13464 0 sb_0__1_.mux_right_track_38.out
rlabel metal1 29578 14246 29578 14246 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34362 14280 34362 14280 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 47058 28764 47058 28764 0 sb_0__1_.mux_right_track_4.out
rlabel metal1 40388 37230 40388 37230 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39514 37162 39514 37162 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 39744 34714 39744 34714 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35650 33014 35650 33014 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 43286 30736 43286 30736 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 44482 12240 44482 12240 0 sb_0__1_.mux_right_track_40.out
rlabel metal2 29670 15368 29670 15368 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37766 13294 37766 13294 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 43746 11730 43746 11730 0 sb_0__1_.mux_right_track_44.out
rlabel metal1 33580 15402 33580 15402 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 39146 14790 39146 14790 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 45172 11730 45172 11730 0 sb_0__1_.mux_right_track_46.out
rlabel metal1 34822 17102 34822 17102 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40112 14382 40112 14382 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 44390 12444 44390 12444 0 sb_0__1_.mux_right_track_48.out
rlabel metal1 37858 16490 37858 16490 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 39514 15164 39514 15164 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 44206 13294 44206 13294 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 38318 18394 38318 18394 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34040 15946 34040 15946 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 39790 16524 39790 16524 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 44206 10540 44206 10540 0 sb_0__1_.mux_right_track_52.out
rlabel metal1 36570 14450 36570 14450 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40756 11730 40756 11730 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 42734 9486 42734 9486 0 sb_0__1_.mux_right_track_54.out
rlabel metal1 35420 12750 35420 12750 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40434 10642 40434 10642 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 43378 10506 43378 10506 0 sb_0__1_.mux_right_track_56.out
rlabel metal1 37766 15062 37766 15062 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 41400 12206 41400 12206 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 44850 29614 44850 29614 0 sb_0__1_.mux_right_track_6.out
rlabel metal1 40572 43078 40572 43078 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40618 38522 40618 38522 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38456 34170 38456 34170 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 42918 36822 42918 36822 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 40756 36346 40756 36346 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 42596 36550 42596 36550 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 47242 30090 47242 30090 0 sb_0__1_.mux_right_track_8.out
rlabel metal1 39008 40562 39008 40562 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39238 39066 39238 39066 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36708 35462 36708 35462 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 39008 39474 39008 39474 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38686 39066 38686 39066 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 43838 36244 43838 36244 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24196 47770 24196 47770 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 23368 41718 23368 41718 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33764 41514 33764 41514 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30774 34714 30774 34714 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24794 36346 24794 36346 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26680 41786 26680 41786 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 26128 43282 26128 43282 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 25346 47634 25346 47634 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21022 50218 21022 50218 0 sb_0__1_.mux_top_track_10.out
rlabel metal1 25438 37230 25438 37230 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 27002 36618 27002 36618 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26496 33490 26496 33490 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25300 33490 25300 33490 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 25530 37638 25530 37638 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 25116 33626 25116 33626 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 22172 43758 22172 43758 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21206 49130 21206 49130 0 sb_0__1_.mux_top_track_12.out
rlabel metal1 28980 32946 28980 32946 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36202 30838 36202 30838 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23322 30294 23322 30294 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28014 33082 28014 33082 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24840 33830 24840 33830 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22448 42194 22448 42194 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 26726 48756 26726 48756 0 sb_0__1_.mux_top_track_2.out
rlabel metal1 33396 39270 33396 39270 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37536 34918 37536 34918 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 26634 32606 26634 32606 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 30866 40358 30866 40358 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30866 37094 30866 37094 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 27370 45934 27370 45934 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19412 49198 19412 49198 0 sb_0__1_.mux_top_track_20.out
rlabel metal1 30590 32742 30590 32742 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37398 30600 37398 30600 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22218 29682 22218 29682 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 29762 32776 29762 32776 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23230 33830 23230 33830 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 20976 42194 20976 42194 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 16882 46614 16882 46614 0 sb_0__1_.mux_top_track_28.out
rlabel metal1 25668 35054 25668 35054 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28152 31994 28152 31994 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20976 36754 20976 36754 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18538 36754 18538 36754 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19458 40052 19458 40052 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 15962 48722 15962 48722 0 sb_0__1_.mux_top_track_36.out
rlabel metal1 28750 38386 28750 38386 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27738 38454 27738 38454 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22172 37094 22172 37094 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20148 45866 20148 45866 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24610 45050 24610 45050 0 sb_0__1_.mux_top_track_4.out
rlabel metal1 32614 36890 32614 36890 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36892 33626 36892 33626 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26450 34986 26450 34986 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32338 36856 32338 36856 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26036 35258 26036 35258 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 26220 44846 26220 44846 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19550 45832 19550 45832 0 sb_0__1_.mux_top_track_44.out
rlabel metal2 28934 39100 28934 39100 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23414 37094 23414 37094 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20884 45934 20884 45934 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20930 46648 20930 46648 0 sb_0__1_.mux_top_track_52.out
rlabel metal1 38870 35054 38870 35054 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36248 35258 36248 35258 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 28750 35190 28750 35190 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21114 43214 21114 43214 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22862 45050 22862 45050 0 sb_0__1_.mux_top_track_6.out
rlabel metal2 27554 38556 27554 38556 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37582 36346 37582 36346 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27232 34646 27232 34646 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23230 31382 23230 31382 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26726 38522 26726 38522 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 25116 34714 25116 34714 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 23828 44846 23828 44846 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 48622 2404 48622 2404 0 test_enable_bottom_in
rlabel metal2 49358 2098 49358 2098 0 test_enable_bottom_out
rlabel metal1 49450 53142 49450 53142 0 test_enable_top_out
rlabel metal3 820 45764 820 45764 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 820 48076 820 48076 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 820 50388 820 50388 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 820 52700 820 52700 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 57000
<< end >>
